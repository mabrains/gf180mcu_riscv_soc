magic
tech gf180mcuD
magscale 1 10
timestamp 1700952943
<< metal1 >>
rect 346882 35198 346894 35250
rect 346946 35247 346958 35250
rect 350018 35247 350030 35250
rect 346946 35201 350030 35247
rect 346946 35198 346958 35201
rect 350018 35198 350030 35201
rect 350082 35198 350094 35250
rect 344194 33630 344206 33682
rect 344258 33630 344270 33682
rect 344209 33231 344255 33630
rect 344306 33231 344318 33234
rect 344209 33185 344318 33231
rect 344306 33182 344318 33185
rect 344370 33182 344382 33234
rect 343410 23438 343422 23490
rect 343474 23487 343486 23490
rect 349682 23487 349694 23490
rect 343474 23441 349694 23487
rect 343474 23438 343486 23441
rect 349682 23438 349694 23441
rect 349746 23438 349758 23490
<< via1 >>
rect 346894 35198 346946 35250
rect 350030 35198 350082 35250
rect 344206 33630 344258 33682
rect 344318 33182 344370 33234
rect 343422 23438 343474 23490
rect 349694 23438 349746 23490
<< metal2 >>
rect 11032 595672 11256 597000
rect 33096 595672 33320 597000
rect 55160 595672 55384 597000
rect 11004 595560 11256 595672
rect 33068 595560 33320 595672
rect 55132 595560 55384 595672
rect 77224 595560 77448 597000
rect 99288 595672 99512 597000
rect 121352 595672 121576 597000
rect 143416 595672 143640 597000
rect 165480 595672 165704 597000
rect 187544 595672 187768 597000
rect 99260 595560 99512 595672
rect 121324 595560 121576 595672
rect 143388 595560 143640 595672
rect 165452 595560 165704 595672
rect 187516 595560 187768 595672
rect 209608 595672 209832 597000
rect 209608 595560 209860 595672
rect 231672 595560 231896 597000
rect 253736 595560 253960 597000
rect 275800 595672 276024 597000
rect 297864 595672 298088 597000
rect 275800 595560 276052 595672
rect 297864 595560 298116 595672
rect 319928 595560 320152 597000
rect 341992 595672 342216 597000
rect 364056 595672 364280 597000
rect 341992 595560 342244 595672
rect 364056 595560 364308 595672
rect 386120 595560 386344 597000
rect 408184 595672 408408 597000
rect 430248 595672 430472 597000
rect 408184 595560 408436 595672
rect 430248 595560 430500 595672
rect 452312 595560 452536 597000
rect 474376 595672 474600 597000
rect 496440 595672 496664 597000
rect 474376 595560 474628 595672
rect 496440 595560 496692 595672
rect 518504 595560 518728 597000
rect 540568 595672 540792 597000
rect 540568 595560 540820 595672
rect 562632 595560 562856 597000
rect 584696 595560 584920 597000
rect 11004 204148 11060 595560
rect 11004 204082 11060 204092
rect 33068 198548 33124 595560
rect 40908 590772 40964 590782
rect 40796 590660 40852 590670
rect 40684 590548 40740 590558
rect 40236 589652 40292 589662
rect 40236 209972 40292 589596
rect 40684 221396 40740 590492
rect 40796 225204 40852 590604
rect 40796 225138 40852 225148
rect 40684 221330 40740 221340
rect 40236 209906 40292 209916
rect 33068 198482 33124 198492
rect 40908 194740 40964 590716
rect 55132 590772 55188 595560
rect 55132 590706 55188 590716
rect 77308 589764 77364 595560
rect 77308 589698 77364 589708
rect 99260 589652 99316 595560
rect 99260 589586 99316 589596
rect 41132 589540 41188 589550
rect 41020 589428 41076 589438
rect 41020 217588 41076 589372
rect 41020 217522 41076 217532
rect 41132 206164 41188 589484
rect 121324 589540 121380 595560
rect 143388 590660 143444 595560
rect 143388 590594 143444 590604
rect 165452 590548 165508 595560
rect 165452 590482 165508 590492
rect 121324 589474 121380 589484
rect 187516 589428 187572 595560
rect 187516 589362 187572 589372
rect 209804 589428 209860 595560
rect 231756 590548 231812 595560
rect 231756 590482 231812 590492
rect 275996 589540 276052 595560
rect 298060 590660 298116 595560
rect 298060 590594 298116 590604
rect 342188 589652 342244 595560
rect 364252 590772 364308 595560
rect 364252 590706 364308 590716
rect 408380 589764 408436 595560
rect 430444 590884 430500 595560
rect 430444 590818 430500 590828
rect 408380 589698 408436 589708
rect 474572 589764 474628 595560
rect 496636 590996 496692 595560
rect 496636 590930 496692 590940
rect 474572 589698 474628 589708
rect 540764 589764 540820 595560
rect 540764 589698 540820 589708
rect 548828 590996 548884 591006
rect 342188 589586 342244 589596
rect 275996 589474 276052 589484
rect 209804 589362 209860 589372
rect 548716 589428 548772 589438
rect 43596 588868 43652 588878
rect 43596 213780 43652 588812
rect 548716 503300 548772 589372
rect 548828 583828 548884 590940
rect 548828 583762 548884 583772
rect 550172 590884 550228 590894
rect 550172 504868 550228 590828
rect 551852 590660 551908 590670
rect 551852 506548 551908 590604
rect 551852 506482 551908 506492
rect 553532 590548 553588 590558
rect 550172 504802 550228 504812
rect 548716 503234 548772 503244
rect 553532 503188 553588 590492
rect 562716 590548 562772 595560
rect 562716 590482 562772 590492
rect 575372 590772 575428 590782
rect 563612 589652 563668 589662
rect 553532 503122 553588 503132
rect 560252 589540 560308 589550
rect 560252 502740 560308 589484
rect 563612 503972 563668 589596
rect 570332 589092 570388 589102
rect 568540 588980 568596 588990
rect 566748 588868 566804 588878
rect 563612 503906 563668 503916
rect 564956 503972 565012 503982
rect 560252 502674 560308 502684
rect 561372 503300 561428 503310
rect 561372 499912 561428 503244
rect 563164 502740 563220 502750
rect 563164 499912 563220 502684
rect 564956 499912 565012 503916
rect 566748 499912 566804 588812
rect 568540 499912 568596 588924
rect 570332 499912 570388 589036
rect 572124 588644 572180 588654
rect 572124 499912 572180 588588
rect 573916 548996 573972 549006
rect 573916 499912 573972 548940
rect 575372 503972 575428 590716
rect 584668 590548 584724 590558
rect 582876 583828 582932 583838
rect 575372 503906 575428 503916
rect 577500 506548 577556 506558
rect 575708 503188 575764 503198
rect 575708 499912 575764 503132
rect 577500 499912 577556 506492
rect 581084 504868 581140 504878
rect 579292 503972 579348 503982
rect 579292 499912 579348 503916
rect 581084 499912 581140 504812
rect 582876 499912 582932 583772
rect 584668 499912 584724 590492
rect 586460 575428 586516 575438
rect 586460 499912 586516 575372
rect 588252 535780 588308 535790
rect 588252 499912 588308 535724
rect 551852 492324 551908 492334
rect 550172 449316 550228 449326
rect 221564 232708 221620 232718
rect 207228 232596 207284 232606
rect 200060 232484 200116 232494
rect 71036 232260 71092 232270
rect 71036 229880 71092 232204
rect 135548 232148 135604 232158
rect 106876 230804 106932 230814
rect 85372 230468 85428 230478
rect 85372 229880 85428 230412
rect 106876 229880 106932 230748
rect 114044 230692 114100 230702
rect 114044 229880 114100 230636
rect 135548 229880 135604 232092
rect 171388 230580 171444 230590
rect 149884 230244 149940 230254
rect 149884 229880 149940 230188
rect 157052 229908 157108 229918
rect 171388 229880 171444 230524
rect 185724 230356 185780 230366
rect 179228 230020 179284 230030
rect 179228 229908 179284 229964
rect 178584 229852 179284 229908
rect 185724 229880 185780 230300
rect 200060 229880 200116 232428
rect 207228 229880 207284 232540
rect 214396 232372 214452 232382
rect 214396 229880 214452 232316
rect 221564 229880 221620 232652
rect 242956 232708 243012 232718
rect 228732 232036 228788 232046
rect 228732 229880 228788 231980
rect 240156 232036 240212 232046
rect 235900 231924 235956 231934
rect 235900 229880 235956 231868
rect 157052 229842 157108 229852
rect 121212 229796 121268 229806
rect 121212 229730 121268 229740
rect 92540 229684 92596 229694
rect 92540 229618 92596 229628
rect 164220 229572 164276 229582
rect 164220 229506 164276 229516
rect 78652 229460 78708 229470
rect 78232 229404 78652 229460
rect 78652 229394 78708 229404
rect 128380 229460 128436 229470
rect 128380 229394 128436 229404
rect 63868 229348 63924 229358
rect 63868 229282 63924 229292
rect 192892 229348 192948 229358
rect 192892 229282 192948 229292
rect 240156 224308 240212 231980
rect 242732 231924 242788 231934
rect 240156 224242 240212 224252
rect 241948 229684 242004 229694
rect 241948 222740 242004 229628
rect 241948 222674 242004 222684
rect 242732 217588 242788 231868
rect 242956 217700 243012 232652
rect 549388 232484 549444 232494
rect 247772 232372 247828 232382
rect 243628 232260 243684 232270
rect 243628 224532 243684 232204
rect 246876 230804 246932 230814
rect 243628 224466 243684 224476
rect 244412 229796 244468 229806
rect 242956 217634 243012 217644
rect 242732 217522 242788 217532
rect 43596 213714 43652 213724
rect 41132 206098 41188 206108
rect 53788 204148 53844 204158
rect 53788 202356 53844 204092
rect 53788 202290 53844 202300
rect 40908 194674 40964 194684
rect 244412 172228 244468 229740
rect 246876 222628 246932 230748
rect 246876 222562 246932 222572
rect 247772 219492 247828 232316
rect 315868 232148 315924 232158
rect 247772 219426 247828 219436
rect 289884 230692 289940 230702
rect 244412 172162 244468 172172
rect 289884 169960 289940 230636
rect 315868 224420 315924 232092
rect 409836 230580 409892 230590
rect 391916 230468 391972 230478
rect 375340 227892 375396 227902
rect 315868 224354 315924 224364
rect 358764 224532 358820 224542
rect 358764 219912 358820 224476
rect 375340 219912 375396 227836
rect 391916 219912 391972 230412
rect 408492 222740 408548 222750
rect 408492 219912 408548 222684
rect 409836 222740 409892 230524
rect 505148 230356 505204 230366
rect 474796 230244 474852 230254
rect 456764 229908 456820 229918
rect 424956 227668 425012 227678
rect 424956 223412 425012 227612
rect 456764 223412 456820 229852
rect 424956 223356 425124 223412
rect 409836 222674 409892 222684
rect 425068 219912 425124 223356
rect 456764 223346 456820 223356
rect 458220 223412 458276 223422
rect 441644 222628 441700 222638
rect 441644 219912 441700 222572
rect 458220 219912 458276 223356
rect 474796 219912 474852 230188
rect 491372 229572 491428 229582
rect 491372 219912 491428 229516
rect 505148 223412 505204 230300
rect 524076 230020 524132 230030
rect 505148 223346 505204 223356
rect 507948 223412 508004 223422
rect 507948 219912 508004 223356
rect 524076 223300 524132 229964
rect 524076 223244 524580 223300
rect 524524 219912 524580 223244
rect 541100 222740 541156 222750
rect 541100 219912 541156 222684
rect 347228 219716 347284 219726
rect 343532 215908 343588 215918
rect 309820 172228 309876 172238
rect 309820 169960 309876 172172
rect 289884 67228 289940 70056
rect 289772 67172 289940 67228
rect 289772 65604 289828 67172
rect 242844 52948 242900 52958
rect 239372 51604 239428 51614
rect 239372 31108 239428 51548
rect 242732 49252 242788 49262
rect 240268 39508 240324 39518
rect 240156 34468 240212 34478
rect 240156 31332 240212 34412
rect 240268 32564 240324 39452
rect 241948 37828 242004 37838
rect 241388 37268 241444 37278
rect 241164 37156 241220 37166
rect 240268 32498 240324 32508
rect 241052 36148 241108 36158
rect 240156 31266 240212 31276
rect 239372 31042 239428 31052
rect 139132 30772 139188 30782
rect 139132 30706 139188 30716
rect 140924 30772 140980 30782
rect 140924 30706 140980 30716
rect 142716 30772 142772 30782
rect 142716 30706 142772 30716
rect 149884 30772 149940 30782
rect 149884 30706 149940 30716
rect 137340 30660 137396 30670
rect 137340 30548 137396 30604
rect 137228 30520 137396 30548
rect 151676 30660 151732 30670
rect 151676 30548 151732 30604
rect 153468 30660 153524 30670
rect 153468 30548 153524 30604
rect 158844 30660 158900 30670
rect 158844 30548 158900 30604
rect 160636 30660 160692 30670
rect 160636 30548 160692 30604
rect 162428 30660 162484 30670
rect 162428 30548 162484 30604
rect 185724 30660 185780 30670
rect 185724 30548 185780 30604
rect 191100 30660 191156 30670
rect 191100 30548 191156 30604
rect 196476 30660 196532 30670
rect 196476 30548 196532 30604
rect 151676 30520 151844 30548
rect 153468 30520 153636 30548
rect 158844 30520 159012 30548
rect 160636 30520 160804 30548
rect 162428 30520 162596 30548
rect 137228 30492 137368 30520
rect 151704 30492 151844 30520
rect 153496 30492 153636 30520
rect 158872 30492 159012 30520
rect 160664 30492 160804 30520
rect 162456 30492 162596 30520
rect 135548 30436 135604 30446
rect 105084 30324 105140 30334
rect 134428 30324 134484 30334
rect 133784 30268 134428 30324
rect 96124 30212 96180 30222
rect 81788 30100 81844 30110
rect 69272 30044 71064 30100
rect 74648 30072 78232 30100
rect 69692 26964 69748 30044
rect 58940 26628 58996 26638
rect 45612 26516 45668 26526
rect 13244 26068 13300 26078
rect 11340 12628 11396 12638
rect 11340 480 11396 12572
rect 13244 480 13300 26012
rect 27692 24500 27748 24510
rect 18956 19460 19012 19470
rect 15148 14308 15204 14318
rect 15148 480 15204 14252
rect 17276 6580 17332 6590
rect 17276 480 17332 6524
rect 11340 392 11592 480
rect 13244 392 13496 480
rect 15148 392 15400 480
rect 11368 -960 11592 392
rect 13272 -960 13496 392
rect 15176 -960 15400 392
rect 17080 392 17332 480
rect 18956 480 19012 19404
rect 22764 17892 22820 17902
rect 21980 7588 22036 7598
rect 21868 7532 21980 7588
rect 21868 3444 21924 7532
rect 21980 7522 22036 7532
rect 21756 3388 21924 3444
rect 21084 480 21252 532
rect 18956 392 19208 480
rect 17080 -960 17304 392
rect 18984 -960 19208 392
rect 20888 476 21252 480
rect 20888 392 21140 476
rect 21196 420 21252 476
rect 21756 420 21812 3388
rect 20888 -960 21112 392
rect 21196 364 21812 420
rect 22764 480 22820 17836
rect 24892 4340 24948 4350
rect 24892 480 24948 4284
rect 27692 4340 27748 24444
rect 27692 4274 27748 4284
rect 27916 24388 27972 24398
rect 26796 4228 26852 4238
rect 26796 480 26852 4172
rect 27916 4228 27972 24332
rect 41804 21252 41860 21262
rect 37996 19684 38052 19694
rect 32284 19348 32340 19358
rect 30380 16212 30436 16222
rect 27916 4162 27972 4172
rect 28700 7700 28756 7710
rect 28700 480 28756 7644
rect 22764 392 23016 480
rect 22792 -960 23016 392
rect 24696 392 24948 480
rect 26600 392 26852 480
rect 28504 392 28756 480
rect 30380 480 30436 16156
rect 32284 480 32340 19292
rect 34412 10948 34468 10958
rect 34412 480 34468 10892
rect 36316 9380 36372 9390
rect 36316 480 36372 9324
rect 30380 392 30632 480
rect 32284 392 32536 480
rect 24696 -960 24920 392
rect 26600 -960 26824 392
rect 28504 -960 28728 392
rect 30408 -960 30632 392
rect 32312 -960 32536 392
rect 34216 392 34468 480
rect 36120 392 36372 480
rect 37996 480 38052 19628
rect 41132 16100 41188 16110
rect 40124 4228 40180 4238
rect 40124 480 40180 4172
rect 41132 4228 41188 16044
rect 41132 4162 41188 4172
rect 37996 392 38248 480
rect 34216 -960 34440 392
rect 36120 -960 36344 392
rect 38024 -960 38248 392
rect 39928 392 40180 480
rect 41804 480 41860 21196
rect 43932 5908 43988 5918
rect 43932 480 43988 5852
rect 41804 392 42056 480
rect 39928 -960 40152 392
rect 41832 -960 42056 392
rect 43736 392 43988 480
rect 45612 480 45668 26460
rect 53228 24724 53284 24734
rect 47516 17668 47572 17678
rect 47516 480 47572 17612
rect 49420 14420 49476 14430
rect 49420 480 49476 14364
rect 51548 7812 51604 7822
rect 51548 480 51604 7756
rect 45612 392 45864 480
rect 47516 392 47768 480
rect 49420 392 49672 480
rect 43736 -960 43960 392
rect 45640 -960 45864 392
rect 47544 -960 47768 392
rect 49448 -960 49672 392
rect 51352 392 51604 480
rect 53228 480 53284 24668
rect 55132 21364 55188 21374
rect 55132 480 55188 21308
rect 57260 4228 57316 4238
rect 57260 480 57316 4172
rect 53228 392 53480 480
rect 55132 392 55384 480
rect 51352 -960 51576 392
rect 53256 -960 53480 392
rect 55160 -960 55384 392
rect 57064 392 57316 480
rect 58940 480 58996 26572
rect 66556 24612 66612 24622
rect 62748 15988 62804 15998
rect 59612 12740 59668 12750
rect 59612 4228 59668 12684
rect 59612 4162 59668 4172
rect 61068 4228 61124 4238
rect 61068 480 61124 4172
rect 58940 392 59192 480
rect 57064 -960 57288 392
rect 58968 -960 59192 392
rect 60872 392 61124 480
rect 62748 480 62804 15932
rect 62972 14532 63028 14542
rect 62972 4228 63028 14476
rect 62972 4162 63028 4172
rect 64652 12964 64708 12974
rect 64652 480 64708 12908
rect 66556 480 66612 24556
rect 68460 17780 68516 17790
rect 68460 480 68516 17724
rect 69692 12628 69748 26908
rect 72828 26964 72884 30072
rect 72828 26898 72884 26908
rect 74620 30044 78260 30072
rect 69692 12562 69748 12572
rect 72268 26292 72324 26302
rect 70476 6020 70532 6030
rect 70476 480 70532 5964
rect 72268 480 72324 26236
rect 74620 26068 74676 30044
rect 74620 26002 74676 26012
rect 77980 25956 78036 25966
rect 76300 6132 76356 6142
rect 74396 5012 74452 5022
rect 74396 480 74452 4956
rect 76300 480 76356 6076
rect 62748 392 63000 480
rect 64652 392 64904 480
rect 66556 392 66808 480
rect 68460 392 68712 480
rect 60872 -960 61096 392
rect 62776 -960 63000 392
rect 64680 -960 64904 392
rect 66584 -960 66808 392
rect 68488 -960 68712 392
rect 70392 -960 70616 480
rect 72268 392 72520 480
rect 72296 -960 72520 392
rect 74200 392 74452 480
rect 76104 392 76356 480
rect 77980 480 78036 25900
rect 78204 21700 78260 30044
rect 78204 21634 78260 21644
rect 79772 30044 80024 30100
rect 88956 30100 89012 30110
rect 79772 20188 79828 30044
rect 81788 27412 81844 30044
rect 81788 27346 81844 27356
rect 79212 20132 79828 20188
rect 79212 19460 79268 20132
rect 79212 10052 79268 19404
rect 79212 9986 79268 9996
rect 81452 19460 81508 19470
rect 81452 5012 81508 19404
rect 83580 7588 83636 30072
rect 83580 7522 83636 7532
rect 83692 19572 83748 19582
rect 81452 4946 81508 4956
rect 82012 6804 82068 6814
rect 80108 4228 80164 4238
rect 80108 480 80164 4172
rect 82012 480 82068 6748
rect 77980 392 78232 480
rect 74200 -960 74424 392
rect 76104 -960 76328 392
rect 78008 -960 78232 392
rect 79912 392 80164 480
rect 81816 392 82068 480
rect 83692 480 83748 19516
rect 85372 8260 85428 30072
rect 86492 13412 86548 13422
rect 85372 6804 85428 8204
rect 85372 6738 85428 6748
rect 85820 9268 85876 9278
rect 85820 480 85876 9212
rect 86492 6132 86548 13356
rect 87164 13412 87220 30072
rect 87164 13346 87220 13356
rect 86492 6066 86548 6076
rect 87500 7588 87556 7598
rect 83692 392 83944 480
rect 79912 -960 80136 392
rect 81816 -960 82040 392
rect 83720 -960 83944 392
rect 85624 392 85876 480
rect 87500 480 87556 7532
rect 88956 6020 89012 30044
rect 90748 28420 90804 30072
rect 90748 28354 90804 28364
rect 91532 28420 91588 28430
rect 91308 26180 91364 26190
rect 89852 24276 89908 24286
rect 88956 5954 89012 5964
rect 89404 12852 89460 12862
rect 89404 480 89460 12796
rect 89852 4228 89908 24220
rect 89852 4162 89908 4172
rect 91308 480 91364 26124
rect 91532 12964 91588 28364
rect 92540 28196 92596 30072
rect 92540 26628 92596 28140
rect 92540 26562 92596 26572
rect 94332 29876 94388 30072
rect 94332 24724 94388 29820
rect 96124 26516 96180 30156
rect 96124 26450 96180 26460
rect 97916 29876 97972 30072
rect 94332 24658 94388 24668
rect 95116 26068 95172 26078
rect 91532 12898 91588 12908
rect 93436 2548 93492 2558
rect 93436 480 93492 2492
rect 87500 392 87752 480
rect 89404 392 89656 480
rect 91308 392 91560 480
rect 85624 -960 85848 392
rect 87528 -960 87752 392
rect 89432 -960 89656 392
rect 91336 -960 91560 392
rect 93240 392 93492 480
rect 95116 480 95172 26012
rect 97916 19684 97972 29820
rect 97916 19618 97972 19628
rect 99708 23492 99764 30072
rect 99708 16212 99764 23436
rect 101500 24836 101556 30072
rect 99708 16146 99764 16156
rect 100828 18004 100884 18014
rect 97020 12628 97076 12638
rect 97020 480 97076 12572
rect 99036 2660 99092 2670
rect 99036 480 99092 2604
rect 100828 480 100884 17948
rect 101500 17892 101556 24780
rect 101500 17826 101556 17836
rect 103292 18452 103348 30072
rect 105084 27412 105140 30268
rect 105084 27346 105140 27356
rect 106652 30044 106904 30100
rect 108332 30044 108696 30100
rect 106652 28308 106708 30044
rect 102732 16212 102788 16222
rect 102732 480 102788 16156
rect 103292 7812 103348 18396
rect 103292 7746 103348 7756
rect 106540 16324 106596 16334
rect 104860 2772 104916 2782
rect 104860 480 104916 2716
rect 95116 392 95368 480
rect 97020 392 97272 480
rect 93240 -960 93464 392
rect 95144 -960 95368 392
rect 97048 -960 97272 392
rect 98952 -960 99176 480
rect 100828 392 101080 480
rect 102732 392 102984 480
rect 100856 -960 101080 392
rect 102760 -960 102984 392
rect 104664 392 104916 480
rect 106540 480 106596 16268
rect 106652 9380 106708 28252
rect 106652 9314 106708 9324
rect 108332 20132 108388 30044
rect 110460 28532 110516 30072
rect 110460 28466 110516 28476
rect 112252 28532 112308 30072
rect 112252 28466 112308 28476
rect 112588 28756 112644 28766
rect 112588 28196 112644 28700
rect 112588 28130 112644 28140
rect 114044 27748 114100 30072
rect 115836 27860 115892 30072
rect 117516 29428 117572 29438
rect 117516 28308 117572 29372
rect 117516 28242 117572 28252
rect 115836 27794 115892 27804
rect 114044 27682 114100 27692
rect 117628 27636 117684 30072
rect 117628 27570 117684 27580
rect 119420 22708 119476 30072
rect 121212 27524 121268 30072
rect 123004 28084 123060 30072
rect 124796 28196 124852 30072
rect 124796 28130 124852 28140
rect 123004 28018 123060 28028
rect 121212 27458 121268 27468
rect 119420 22642 119476 22652
rect 108332 7700 108388 20076
rect 125580 21588 125636 21598
rect 117964 19796 118020 19806
rect 114380 9492 114436 9502
rect 108332 7634 108388 7644
rect 108668 9380 108724 9390
rect 108668 480 108724 9324
rect 112476 6244 112532 6254
rect 110572 2884 110628 2894
rect 110572 480 110628 2828
rect 112476 480 112532 6188
rect 114380 480 114436 9436
rect 116284 2996 116340 3006
rect 116284 480 116340 2940
rect 106540 392 106792 480
rect 104664 -960 104888 392
rect 106568 -960 106792 392
rect 108472 392 108724 480
rect 110376 392 110628 480
rect 112280 392 112532 480
rect 114184 392 114436 480
rect 116088 392 116340 480
rect 117964 480 118020 19740
rect 119868 17892 119924 17902
rect 119868 480 119924 17836
rect 123676 13076 123732 13086
rect 121996 5908 122052 5918
rect 121996 480 122052 5852
rect 117964 392 118216 480
rect 119868 392 120120 480
rect 108472 -960 108696 392
rect 110376 -960 110600 392
rect 112280 -960 112504 392
rect 114184 -960 114408 392
rect 116088 -960 116312 392
rect 117992 -960 118216 392
rect 119896 -960 120120 392
rect 121800 392 122052 480
rect 123676 480 123732 13020
rect 125580 480 125636 21532
rect 126588 21140 126644 30072
rect 126588 21074 126644 21084
rect 128380 21028 128436 30072
rect 128380 20962 128436 20972
rect 129388 26964 129444 26974
rect 127596 6020 127652 6030
rect 127596 480 127652 5964
rect 129388 480 129444 26908
rect 130172 26516 130228 30072
rect 131964 28532 132020 30072
rect 131964 28466 132020 28476
rect 134428 26908 134484 30268
rect 135548 26964 135604 30380
rect 137228 30100 137284 30492
rect 151788 30100 151844 30492
rect 153580 30100 153636 30492
rect 158956 30100 159012 30492
rect 160748 30100 160804 30492
rect 162540 30100 162596 30492
rect 185612 30520 185780 30548
rect 190988 30520 191156 30548
rect 196364 30520 196532 30548
rect 198268 30660 198324 30670
rect 198268 30548 198324 30604
rect 200060 30660 200116 30670
rect 200060 30548 200116 30604
rect 198268 30520 198436 30548
rect 200060 30520 200228 30548
rect 185612 30492 185752 30520
rect 190988 30492 191128 30520
rect 196364 30492 196504 30520
rect 198296 30492 198436 30520
rect 200088 30492 200228 30520
rect 185612 30100 185668 30492
rect 190988 30100 191044 30492
rect 196364 30100 196420 30492
rect 198380 30100 198436 30492
rect 200172 30100 200228 30492
rect 137228 30072 137368 30100
rect 137228 30044 137396 30072
rect 134428 26852 134596 26908
rect 135548 26898 135604 26908
rect 130172 26450 130228 26460
rect 134540 20188 134596 26852
rect 134540 20132 135156 20188
rect 131292 19684 131348 19694
rect 131292 480 131348 19628
rect 133420 6132 133476 6142
rect 133420 480 133476 6076
rect 123676 392 123928 480
rect 125580 392 125832 480
rect 121800 -960 122024 392
rect 123704 -960 123928 392
rect 125608 -960 125832 392
rect 127512 -960 127736 480
rect 129388 392 129640 480
rect 131292 392 131544 480
rect 129416 -960 129640 392
rect 131320 -960 131544 392
rect 133224 392 133476 480
rect 135100 480 135156 20132
rect 137340 13076 137396 30044
rect 137340 13010 137396 13020
rect 140812 28420 140868 28430
rect 137004 12964 137060 12974
rect 137004 480 137060 12908
rect 139132 480 139300 532
rect 135100 392 135352 480
rect 137004 392 137256 480
rect 133224 -960 133448 392
rect 135128 -960 135352 392
rect 137032 -960 137256 392
rect 138936 476 139300 480
rect 138936 392 139188 476
rect 138936 -960 139160 392
rect 139244 84 139300 476
rect 140812 480 140868 28364
rect 144508 24948 144564 30072
rect 146300 26740 146356 30072
rect 147868 30044 148120 30100
rect 151704 30072 151844 30100
rect 153496 30072 153636 30100
rect 156268 30072 157080 30100
rect 158872 30072 159012 30100
rect 160664 30072 160804 30100
rect 162456 30072 162596 30100
rect 151676 30044 151844 30072
rect 153468 30044 153636 30072
rect 147868 29764 147924 30044
rect 147868 26964 147924 29708
rect 147868 26898 147924 26908
rect 146300 26674 146356 26684
rect 146188 26516 146244 26526
rect 146188 26068 146244 26460
rect 148428 26404 148484 26414
rect 146188 26002 146244 26012
rect 146524 26068 146580 26078
rect 144508 24882 144564 24892
rect 145292 24948 145348 24958
rect 145292 18004 145348 24892
rect 145292 17938 145348 17948
rect 142828 14644 142884 14654
rect 142828 480 142884 14588
rect 144844 480 145012 532
rect 140812 392 141064 480
rect 139244 18 139300 28
rect 140840 -960 141064 392
rect 142744 -960 142968 480
rect 144648 476 145012 480
rect 144648 392 144900 476
rect 144648 -960 144872 392
rect 144956 196 145012 476
rect 146524 480 146580 26012
rect 148428 480 148484 26348
rect 151676 25956 151732 30044
rect 153468 26292 153524 30044
rect 155260 28308 155316 30072
rect 155260 28242 155316 28252
rect 156268 30044 157108 30072
rect 156268 26964 156324 30044
rect 157052 29764 157108 30044
rect 157052 29698 157108 29708
rect 158844 30044 159012 30072
rect 160636 30044 160804 30072
rect 162428 30044 162596 30072
rect 163884 30044 164248 30100
rect 158844 27972 158900 30044
rect 158844 27906 158900 27916
rect 160636 27412 160692 30044
rect 160636 27346 160692 27356
rect 162428 27412 162484 30044
rect 162428 27346 162484 27356
rect 163660 28196 163716 28206
rect 156268 26898 156324 26908
rect 153468 26226 153524 26236
rect 151676 25890 151732 25900
rect 159852 25284 159908 25294
rect 157948 21140 158004 21150
rect 152236 21028 152292 21038
rect 150556 480 150724 532
rect 146524 392 146776 480
rect 148428 392 148680 480
rect 144956 130 145012 140
rect 146552 -960 146776 392
rect 148456 -960 148680 392
rect 150360 476 150724 480
rect 150360 392 150612 476
rect 150360 -960 150584 392
rect 150668 308 150724 476
rect 152236 480 152292 20972
rect 154140 18004 154196 18014
rect 154140 480 154196 17948
rect 156156 6244 156212 6254
rect 156156 480 156212 6188
rect 157948 480 158004 21084
rect 159852 480 159908 25228
rect 163660 24724 163716 28140
rect 161980 480 162148 532
rect 152236 392 152488 480
rect 154140 392 154392 480
rect 150668 242 150724 252
rect 152264 -960 152488 392
rect 154168 -960 154392 392
rect 156072 -960 156296 480
rect 157948 392 158200 480
rect 159852 392 160104 480
rect 157976 -960 158200 392
rect 159880 -960 160104 392
rect 161784 476 162148 480
rect 161784 392 162036 476
rect 162092 420 162148 476
rect 163660 480 163716 24668
rect 163884 25060 163940 30044
rect 163884 19348 163940 25004
rect 166012 25172 166068 30072
rect 167804 28196 167860 30072
rect 167804 28130 167860 28140
rect 166012 24500 166068 25116
rect 166012 24434 166068 24444
rect 169372 28084 169428 28094
rect 163884 19282 163940 19292
rect 169372 21812 169428 28028
rect 169596 28084 169652 30072
rect 171388 28308 171444 30072
rect 173180 28420 173236 30072
rect 173180 28354 173236 28364
rect 171388 28242 171444 28252
rect 169596 28018 169652 28028
rect 174972 27972 175028 30072
rect 174972 27906 175028 27916
rect 175084 27524 175140 27534
rect 165788 7700 165844 7710
rect 165788 480 165844 7644
rect 167692 6356 167748 6366
rect 167692 480 167748 6300
rect 162652 420 162708 430
rect 161784 -960 162008 392
rect 162092 364 162652 420
rect 163660 392 163912 480
rect 162652 354 162708 364
rect 163688 -960 163912 392
rect 165592 392 165844 480
rect 167496 392 167748 480
rect 169372 480 169428 21756
rect 171388 25396 171444 25406
rect 171388 480 171444 25340
rect 174636 7812 174692 7822
rect 174636 6580 174692 7756
rect 174636 6514 174692 6524
rect 173404 6468 173460 6478
rect 173404 480 173460 6412
rect 169372 392 169624 480
rect 165592 -960 165816 392
rect 167496 -960 167720 392
rect 169400 -960 169624 392
rect 171304 -960 171528 480
rect 173208 392 173460 480
rect 175084 480 175140 27468
rect 176316 27524 176372 27534
rect 176316 26628 176372 27468
rect 176316 26562 176372 26572
rect 176764 17668 176820 30072
rect 176764 17602 176820 17612
rect 176988 23380 177044 23390
rect 176988 17556 177044 23324
rect 178556 23380 178612 30072
rect 178556 23314 178612 23324
rect 180348 25396 180404 30072
rect 182168 30044 182308 30100
rect 180348 23044 180404 25340
rect 180348 22978 180404 22988
rect 176988 480 177044 17500
rect 180796 22708 180852 22718
rect 179116 3108 179172 3118
rect 179116 480 179172 3052
rect 175084 392 175336 480
rect 176988 392 177240 480
rect 173208 -960 173432 392
rect 175112 -960 175336 392
rect 177016 -960 177240 392
rect 178920 392 179172 480
rect 180796 480 180852 22652
rect 182252 20916 182308 30044
rect 183148 30044 183960 30100
rect 185612 30072 185752 30100
rect 185612 30044 185780 30072
rect 183148 25284 183204 30044
rect 183148 24612 183204 25228
rect 183148 24546 183204 24556
rect 182252 7700 182308 20860
rect 185724 18004 185780 30044
rect 186284 27972 186340 27982
rect 186284 27524 186340 27916
rect 186284 27458 186340 27468
rect 186508 27972 186564 27982
rect 186508 27636 186564 27916
rect 185724 17938 185780 17948
rect 182252 7634 182308 7644
rect 182700 17668 182756 17678
rect 182700 480 182756 17612
rect 184828 7700 184884 7710
rect 184828 5124 184884 7644
rect 184716 5068 184884 5124
rect 184716 480 184772 5068
rect 186508 480 186564 27580
rect 187516 26404 187572 30072
rect 187516 26338 187572 26348
rect 188412 29764 188468 29774
rect 188412 27524 188468 29708
rect 188412 480 188468 27468
rect 189308 23268 189364 30072
rect 189308 14644 189364 23212
rect 189308 14578 189364 14588
rect 190316 30044 191128 30100
rect 196364 30072 196504 30100
rect 198296 30072 198436 30100
rect 200088 30072 200228 30100
rect 190316 12964 190372 30044
rect 190316 12898 190372 12908
rect 192220 27972 192276 27982
rect 190540 7924 190596 7934
rect 190540 480 190596 7868
rect 180796 392 181048 480
rect 182700 392 182952 480
rect 178920 -960 179144 392
rect 180824 -960 181048 392
rect 182728 -960 182952 392
rect 184632 -960 184856 480
rect 186508 392 186760 480
rect 188412 392 188664 480
rect 186536 -960 186760 392
rect 188440 -960 188664 392
rect 190344 392 190596 480
rect 192220 480 192276 27916
rect 192332 24500 192388 24510
rect 192332 19684 192388 24444
rect 192892 24500 192948 30072
rect 194124 28532 194180 28542
rect 192892 24434 192948 24444
rect 193228 26292 193284 26302
rect 193228 21588 193284 26236
rect 193228 21522 193284 21532
rect 192332 19618 192388 19628
rect 194124 480 194180 28476
rect 194684 26292 194740 30072
rect 196364 30044 196532 30072
rect 194684 26226 194740 26236
rect 196476 17892 196532 30044
rect 198268 30044 198436 30072
rect 200060 30044 200228 30072
rect 196476 17826 196532 17836
rect 198156 27748 198212 27758
rect 198156 26516 198212 27692
rect 198156 8428 198212 26460
rect 198268 9492 198324 30044
rect 198268 9426 198324 9436
rect 199948 16884 200004 16894
rect 197932 8372 198212 8428
rect 196252 8036 196308 8046
rect 196252 480 196308 7980
rect 192220 392 192472 480
rect 194124 392 194376 480
rect 190344 -960 190568 392
rect 192248 -960 192472 392
rect 194152 -960 194376 392
rect 196056 392 196308 480
rect 197932 480 197988 8372
rect 199948 480 200004 16828
rect 200060 9380 200116 30044
rect 201852 28532 201908 30072
rect 203532 30044 203672 30100
rect 203532 29764 203588 30044
rect 201852 28466 201908 28476
rect 202412 28532 202468 28542
rect 200732 28308 200788 28318
rect 200732 18228 200788 28252
rect 200732 16884 200788 18172
rect 200732 16818 200788 16828
rect 202412 16212 202468 28476
rect 202412 16146 202468 16156
rect 203532 12628 203588 29708
rect 205436 29540 205492 30072
rect 207256 30044 207508 30100
rect 203532 12562 203588 12572
rect 203644 27636 203700 27646
rect 200060 9314 200116 9324
rect 201964 4228 202020 4238
rect 201964 480 202020 4172
rect 197932 392 198184 480
rect 196056 -960 196280 392
rect 197960 -960 198184 392
rect 199864 -960 200088 480
rect 201768 392 202020 480
rect 203644 480 203700 27580
rect 205436 26180 205492 29484
rect 205436 26114 205492 26124
rect 205548 28084 205604 28094
rect 205548 480 205604 28028
rect 207452 27412 207508 30044
rect 207452 9268 207508 27356
rect 209020 27860 209076 30072
rect 209020 24276 209076 27804
rect 209020 24210 209076 24220
rect 210812 28420 210868 30072
rect 207452 9202 207508 9212
rect 209356 21588 209412 21598
rect 207676 4340 207732 4350
rect 207676 480 207732 4284
rect 203644 392 203896 480
rect 205548 392 205800 480
rect 201768 -960 201992 392
rect 203672 -960 203896 392
rect 205576 -960 205800 392
rect 207480 392 207732 480
rect 209356 480 209412 21532
rect 210812 19460 210868 28364
rect 212492 30044 212632 30100
rect 214172 30044 214424 30100
rect 215852 30044 216216 30100
rect 217532 30044 218008 30100
rect 219800 30044 219940 30100
rect 212492 28308 212548 30044
rect 210812 19394 210868 19404
rect 211260 28196 211316 28206
rect 211260 18116 211316 28140
rect 211260 480 211316 18060
rect 212492 17780 212548 28252
rect 212492 17714 212548 17724
rect 214172 28196 214228 30044
rect 215852 28532 215908 30044
rect 215852 28466 215908 28476
rect 214172 15988 214228 28140
rect 214172 15922 214228 15932
rect 217532 27748 217588 30044
rect 219884 28532 219940 30044
rect 221564 29652 221620 30072
rect 221564 29586 221620 29596
rect 219884 28466 219940 28476
rect 217532 14420 217588 27692
rect 223356 26180 223412 30072
rect 225176 30044 225988 30100
rect 223356 24388 223412 26124
rect 223356 24322 223412 24332
rect 225932 24388 225988 30044
rect 217532 14354 217588 14364
rect 225932 14308 225988 24332
rect 225932 14242 225988 14252
rect 226940 9268 226996 30072
rect 228732 14308 228788 30072
rect 228732 14242 228788 14252
rect 230524 12628 230580 30072
rect 241052 27972 241108 36092
rect 241164 29876 241220 37100
rect 241388 30212 241444 37212
rect 241500 36260 241556 36270
rect 241500 31220 241556 36204
rect 241948 32900 242004 37772
rect 241948 32834 242004 32844
rect 241500 31154 241556 31164
rect 241388 30146 241444 30156
rect 241164 29810 241220 29820
rect 242732 28084 242788 49196
rect 242844 32452 242900 52892
rect 242844 32386 242900 32396
rect 242956 42868 243012 42878
rect 242956 30772 243012 42812
rect 242956 30706 243012 30716
rect 243068 37380 243124 37390
rect 243068 29988 243124 37324
rect 243068 29922 243124 29932
rect 242732 28018 242788 28028
rect 241052 27906 241108 27916
rect 289772 21700 289828 65548
rect 309820 26852 309876 70056
rect 309820 26786 309876 26796
rect 343420 53956 343476 53966
rect 289772 21634 289828 21644
rect 343420 23490 343476 53900
rect 343532 24388 343588 215852
rect 343644 210084 343700 210094
rect 343644 26180 343700 210028
rect 347228 189028 347284 219660
rect 347564 219604 347620 219614
rect 347340 216916 347396 216926
rect 347340 205828 347396 216860
rect 347340 205762 347396 205772
rect 347452 216804 347508 216814
rect 347452 199780 347508 216748
rect 347452 199714 347508 199724
rect 347564 194404 347620 219548
rect 347676 217028 347732 217038
rect 347676 210084 347732 216972
rect 347676 210018 347732 210028
rect 347564 194338 347620 194348
rect 347228 188962 347284 188972
rect 549388 184436 549444 232428
rect 549388 184370 549444 184380
rect 344316 156772 344372 156782
rect 344204 151396 344260 151406
rect 344092 146020 344148 146030
rect 343980 140644 344036 140654
rect 343868 135268 343924 135278
rect 343756 129892 343812 129902
rect 343756 36260 343812 129836
rect 343756 35588 343812 36204
rect 343756 35522 343812 35532
rect 343868 34244 343924 135212
rect 343868 34178 343924 34188
rect 343756 32900 343812 32910
rect 343980 32900 344036 140588
rect 343812 32844 344036 32900
rect 343756 32676 343812 32844
rect 343756 32610 343812 32620
rect 344092 31556 344148 145964
rect 344204 33682 344260 151340
rect 344316 33908 344372 156716
rect 347004 108388 347060 108398
rect 346780 97636 346836 97646
rect 346668 70756 346724 70766
rect 346108 53844 346164 53854
rect 346108 52948 346164 53788
rect 346108 52882 346164 52892
rect 346668 51940 346724 70700
rect 346668 51874 346724 51884
rect 346780 42868 346836 97580
rect 346780 42802 346836 42812
rect 347004 40964 347060 108332
rect 347452 92260 347508 92270
rect 347340 86884 347396 86894
rect 347228 81508 347284 81518
rect 347116 76132 347172 76142
rect 347116 52052 347172 76076
rect 347116 51986 347172 51996
rect 347228 50372 347284 81452
rect 347228 50306 347284 50316
rect 347340 48468 347396 86828
rect 347340 48402 347396 48412
rect 347452 45444 347508 92204
rect 347564 65380 347620 65390
rect 347564 51604 347620 65324
rect 347676 60004 347732 60014
rect 347676 53844 347732 59948
rect 347676 53778 347732 53788
rect 350364 53844 350420 53854
rect 349804 51940 349860 51950
rect 347564 51538 347620 51548
rect 349580 51604 349636 51614
rect 347452 45378 347508 45388
rect 346892 35250 346948 35262
rect 346892 35198 346894 35250
rect 346946 35198 346948 35250
rect 344316 33852 344484 33908
rect 344204 33630 344206 33682
rect 344258 33630 344260 33682
rect 344204 33618 344260 33630
rect 344428 33460 344484 33852
rect 344092 31490 344148 31500
rect 344204 33404 344484 33460
rect 344204 29540 344260 33404
rect 344316 33234 344372 33246
rect 344316 33182 344318 33234
rect 344370 33182 344372 33234
rect 344316 30212 344372 33182
rect 344316 29764 344372 30156
rect 344316 29698 344372 29708
rect 344204 28868 344260 29484
rect 344204 28802 344260 28812
rect 343644 26114 343700 26124
rect 346108 27860 346164 27870
rect 346108 26180 346164 27804
rect 346108 26114 346164 26124
rect 343532 24322 343588 24332
rect 343420 23438 343422 23490
rect 343474 23438 343476 23490
rect 343420 18228 343476 23438
rect 343420 18162 343476 18172
rect 346892 18116 346948 35198
rect 347004 23268 347060 40908
rect 347004 23202 347060 23212
rect 349580 21476 349636 51548
rect 349692 50372 349748 50382
rect 349692 35140 349748 50316
rect 349692 35074 349748 35084
rect 349580 21410 349636 21420
rect 349692 23490 349748 23502
rect 349692 23438 349694 23490
rect 349746 23438 349748 23490
rect 349692 21364 349748 23438
rect 349692 21298 349748 21308
rect 349804 23156 349860 51884
rect 350140 48804 350196 48814
rect 350028 43652 350084 43662
rect 350028 35250 350084 43596
rect 350028 35198 350030 35250
rect 350082 35198 350084 35250
rect 350028 35186 350084 35198
rect 350140 23380 350196 48748
rect 350140 23314 350196 23324
rect 350364 23268 350420 53788
rect 550060 53060 550116 53070
rect 549388 45556 549444 45566
rect 431788 40740 431844 40750
rect 431788 40674 431844 40684
rect 472108 40740 472164 40750
rect 443884 40628 443940 40638
rect 443884 40562 443940 40572
rect 444108 40628 444164 40638
rect 472108 40628 472164 40684
rect 472108 40600 472388 40628
rect 472136 40572 472388 40600
rect 436268 40516 436324 40526
rect 435148 40460 436268 40516
rect 415660 40068 415716 40078
rect 354508 40012 355208 40068
rect 354508 37716 354564 40012
rect 359212 37828 359268 40040
rect 359212 37762 359268 37772
rect 362908 40012 363272 40068
rect 367052 40012 367304 40068
rect 350364 23202 350420 23212
rect 350812 35140 350868 35150
rect 346892 18050 346948 18060
rect 349804 17668 349860 23100
rect 350812 23044 350868 35084
rect 350812 22978 350868 22988
rect 349804 17602 349860 17612
rect 230524 12562 230580 12572
rect 354508 10052 354564 37660
rect 362908 37044 362964 40012
rect 362908 13412 362964 36988
rect 367052 37492 367108 40012
rect 367052 30100 367108 37436
rect 367052 30034 367108 30044
rect 371308 28644 371364 40040
rect 375340 28756 375396 40040
rect 378812 40012 379400 40068
rect 383432 40012 383908 40068
rect 378812 37380 378868 40012
rect 378812 30100 378868 37324
rect 383852 37268 383908 40012
rect 383852 37044 383908 37212
rect 383852 36978 383908 36988
rect 387436 37156 387492 40040
rect 387436 31948 387492 37100
rect 378812 30034 378868 30044
rect 387212 31892 387492 31948
rect 375340 28690 375396 28700
rect 376236 28756 376292 28766
rect 371308 28578 371364 28588
rect 376236 26404 376292 28700
rect 376236 26338 376292 26348
rect 387212 25844 387268 31892
rect 387212 25778 387268 25788
rect 391468 25956 391524 40040
rect 391468 23492 391524 25900
rect 394828 40012 395528 40068
rect 394828 29652 394884 40012
rect 394828 24836 394884 29596
rect 394828 24770 394884 24780
rect 391468 23426 391524 23436
rect 399532 18452 399588 40040
rect 403564 33012 403620 40040
rect 403564 32946 403620 32956
rect 407596 29428 407652 40040
rect 407596 29362 407652 29372
rect 411628 20132 411684 40040
rect 415660 21588 415716 40012
rect 419692 39732 419748 40040
rect 419692 39666 419748 39676
rect 423388 40012 423752 40068
rect 423388 35364 423444 40012
rect 427756 39844 427812 40040
rect 427756 36148 427812 39788
rect 427756 36082 427812 36092
rect 423388 26516 423444 35308
rect 423388 26450 423444 26460
rect 435148 22708 435204 40460
rect 436268 40450 436324 40460
rect 439852 40180 439908 40190
rect 439852 26628 439908 40124
rect 444108 38668 444164 40572
rect 455980 40516 456036 40526
rect 455980 40450 456036 40460
rect 456204 40516 456260 40526
rect 443996 38612 444164 38668
rect 447916 39844 447972 40040
rect 443996 31948 444052 38612
rect 439852 26562 439908 26572
rect 443884 31892 444052 31948
rect 435148 22642 435204 22652
rect 443884 21812 443940 31892
rect 447916 24724 447972 39788
rect 447916 24658 447972 24668
rect 451948 39508 452004 40040
rect 443884 21746 443940 21756
rect 415660 21522 415716 21532
rect 451948 21140 452004 39452
rect 456204 31948 456260 40460
rect 464044 40404 464100 40414
rect 463708 40348 464044 40404
rect 459228 40040 460040 40068
rect 459228 40012 460068 40040
rect 459228 31948 459284 40012
rect 460012 39396 460068 40012
rect 460012 39330 460068 39340
rect 463708 37380 463764 40348
rect 464044 40338 464100 40348
rect 463708 37314 463764 37324
rect 468076 40292 468132 40302
rect 451948 21074 452004 21084
rect 455980 31892 456260 31948
rect 458668 31892 459284 31948
rect 455980 21028 456036 31892
rect 458668 26068 458724 31892
rect 468076 30324 468132 40236
rect 472332 38668 472388 40572
rect 536648 40124 536900 40180
rect 472108 38612 472388 38668
rect 476140 39284 476196 40040
rect 472108 30436 472164 38612
rect 476140 30548 476196 39228
rect 480172 39732 480228 40040
rect 480172 37716 480228 39676
rect 480172 37650 480228 37660
rect 483868 40012 484232 40068
rect 483868 39732 483924 40012
rect 483868 37716 483924 39676
rect 483868 37650 483924 37660
rect 488236 39732 488292 40040
rect 488236 37716 488292 39676
rect 488236 37650 488292 37660
rect 492268 39508 492324 40040
rect 476140 30482 476196 30492
rect 472108 30370 472164 30380
rect 468076 30258 468132 30268
rect 458668 26002 458724 26012
rect 492268 24948 492324 39452
rect 496300 39732 496356 40040
rect 496300 26740 496356 39676
rect 500332 38164 500388 40040
rect 504392 40012 504868 40068
rect 500332 37044 500388 38108
rect 500332 36978 500388 36988
rect 504812 38500 504868 40012
rect 504812 37044 504868 38444
rect 504812 36978 504868 36988
rect 508396 38388 508452 40040
rect 508396 32788 508452 38332
rect 512428 39396 512484 40040
rect 516460 39732 516516 40040
rect 520520 40012 520772 40068
rect 516460 39666 516516 39676
rect 512428 37044 512484 39340
rect 512428 36978 512484 36988
rect 520716 34580 520772 40012
rect 524524 38612 524580 40040
rect 524524 38546 524580 38556
rect 528556 37044 528612 40040
rect 532588 39732 532644 40040
rect 532588 38052 532644 39676
rect 532588 37986 532644 37996
rect 528556 36978 528612 36988
rect 536732 37940 536788 37950
rect 536844 37940 536900 40124
rect 536788 37884 536900 37940
rect 540092 40012 540680 40068
rect 544712 40012 545188 40068
rect 540092 38052 540148 40012
rect 520716 34514 520772 34524
rect 508396 32722 508452 32732
rect 496300 26674 496356 26684
rect 536732 25060 536788 37884
rect 540092 25172 540148 37996
rect 540092 25106 540148 25116
rect 545132 26852 545188 40012
rect 549388 36484 549444 45500
rect 549388 36418 549444 36428
rect 536732 24994 536788 25004
rect 492268 24882 492324 24892
rect 455980 20962 456036 20972
rect 411628 20066 411684 20076
rect 399532 18386 399588 18396
rect 362908 13346 362964 13356
rect 354508 9986 354564 9996
rect 545132 10052 545188 26796
rect 550060 23268 550116 53004
rect 550172 40628 550228 449260
rect 550172 40562 550228 40572
rect 550284 433188 550340 433198
rect 550284 40292 550340 433132
rect 550396 422436 550452 422446
rect 550396 41412 550452 422380
rect 550620 414372 550676 414382
rect 550396 41346 550452 41356
rect 550508 398244 550564 398254
rect 550284 40226 550340 40236
rect 550508 34580 550564 398188
rect 550620 41524 550676 414316
rect 550620 41458 550676 41468
rect 550732 403620 550788 403630
rect 550732 39396 550788 403564
rect 551404 60340 551460 60350
rect 550956 60228 551012 60238
rect 550732 39330 550788 39340
rect 550844 55748 550900 55758
rect 550508 34514 550564 34524
rect 550844 23380 550900 55692
rect 550956 38500 551012 60172
rect 551404 50428 551460 60284
rect 551404 50372 551684 50428
rect 550956 38434 551012 38444
rect 551628 28308 551684 50372
rect 551740 44996 551796 45006
rect 551740 34916 551796 44940
rect 551740 34850 551796 34860
rect 551852 31948 551908 492268
rect 556892 489636 556948 489646
rect 553644 473508 553700 473518
rect 551964 468132 552020 468142
rect 551964 40068 552020 468076
rect 553532 435876 553588 435886
rect 551964 40002 552020 40012
rect 552076 411684 552132 411694
rect 552076 38164 552132 411628
rect 552076 38098 552132 38108
rect 552188 393204 552244 393214
rect 552188 216916 552244 393148
rect 550844 23314 550900 23324
rect 551516 27076 551572 27086
rect 550060 23202 550116 23212
rect 551516 20804 551572 27020
rect 551628 23492 551684 28252
rect 551740 31892 551908 31948
rect 551740 28420 551796 31892
rect 551740 24836 551796 28364
rect 551740 24770 551796 24780
rect 551964 28532 552020 28542
rect 551628 23426 551684 23436
rect 551964 22148 552020 28476
rect 551964 22082 552020 22092
rect 551516 20738 551572 20748
rect 552188 16772 552244 216860
rect 552300 232596 552356 232606
rect 552300 205044 552356 232540
rect 553196 227780 553252 227790
rect 552972 224308 553028 224318
rect 552860 217588 552916 217598
rect 552300 204988 552804 205044
rect 552748 193956 552804 204988
rect 552748 193890 552804 193900
rect 552860 164388 552916 217532
rect 552972 174244 553028 224252
rect 553084 219492 553140 219502
rect 553084 203812 553140 219436
rect 553084 203746 553140 203756
rect 552972 174178 553028 174188
rect 552860 164322 552916 164332
rect 553196 154532 553252 227724
rect 553196 154466 553252 154476
rect 552524 60452 552580 60462
rect 552412 47684 552468 47694
rect 552300 46340 552356 46350
rect 552300 33572 552356 46284
rect 552412 35140 552468 47628
rect 552412 35074 552468 35084
rect 552300 33506 552356 33516
rect 552524 28532 552580 60396
rect 553532 40404 553588 435820
rect 553644 226884 553700 473452
rect 555212 470820 555268 470830
rect 553644 226818 553700 226828
rect 553756 446628 553812 446638
rect 553532 40338 553588 40348
rect 553756 39844 553812 446572
rect 554652 430500 554708 430510
rect 553868 425124 553924 425134
rect 553868 41188 553924 425068
rect 553868 41122 553924 41132
rect 553980 417060 554036 417070
rect 553756 39778 553812 39788
rect 553980 39508 554036 417004
rect 553980 39442 554036 39452
rect 554092 56532 554148 56542
rect 552524 28466 552580 28476
rect 552300 27748 552356 27758
rect 552300 19460 552356 27692
rect 552300 19394 552356 19404
rect 552636 26964 552692 26974
rect 552636 18116 552692 26908
rect 554092 20188 554148 56476
rect 554652 40740 554708 430444
rect 555212 216580 555268 470764
rect 555212 216514 555268 216524
rect 556108 218484 556164 218494
rect 556108 193284 556164 218428
rect 556220 216804 556276 216814
rect 556220 199892 556276 216748
rect 556220 199826 556276 199836
rect 556108 193218 556164 193228
rect 556668 63252 556724 63262
rect 556668 59864 556724 63196
rect 556892 60340 556948 489580
rect 558572 486948 558628 486958
rect 557676 484260 557732 484270
rect 557004 481572 557060 481582
rect 557004 219604 557060 481516
rect 557228 478884 557284 478894
rect 557004 218484 557060 219548
rect 557004 218418 557060 218428
rect 557116 408996 557172 409006
rect 556892 60274 556948 60284
rect 557116 60228 557172 408940
rect 557228 216804 557284 478828
rect 557452 476196 557508 476206
rect 557228 216738 557284 216748
rect 557340 406308 557396 406318
rect 557116 60162 557172 60172
rect 557340 60004 557396 406252
rect 557452 393204 557508 476140
rect 557452 393138 557508 393148
rect 557676 379764 557732 484204
rect 557676 379698 557732 379708
rect 558572 60452 558628 486892
rect 590492 430164 590548 430174
rect 559468 379764 559524 379774
rect 558684 378868 558740 378878
rect 558684 63252 558740 378812
rect 559468 219716 559524 379708
rect 559468 189812 559524 219660
rect 559468 189746 559524 189756
rect 562716 66388 562772 380072
rect 563388 376516 563444 380072
rect 564060 377524 564116 380072
rect 564060 377458 564116 377468
rect 564732 376852 564788 380072
rect 565404 377300 565460 380072
rect 566076 377412 566132 380072
rect 566076 377346 566132 377356
rect 565404 377234 565460 377244
rect 564732 376786 564788 376796
rect 566748 376628 566804 380072
rect 567420 377412 567476 380072
rect 567420 377346 567476 377356
rect 568092 377300 568148 380072
rect 568092 377234 568148 377244
rect 568764 376740 568820 380072
rect 568764 376674 568820 376684
rect 566748 376562 566804 376572
rect 563388 376450 563444 376460
rect 569436 376516 569492 380072
rect 570108 376628 570164 380072
rect 570808 380044 571060 380100
rect 570108 376562 570164 376572
rect 569436 376450 569492 376460
rect 571004 376516 571060 380044
rect 571452 376628 571508 380072
rect 572152 380044 572628 380100
rect 571452 376562 571508 376572
rect 571004 376450 571060 376460
rect 572572 376516 572628 380044
rect 572572 376450 572628 376460
rect 572796 376516 572852 380072
rect 573468 376628 573524 380072
rect 574168 380044 574532 380100
rect 573468 376562 573524 376572
rect 572796 376450 572852 376460
rect 574476 376516 574532 380044
rect 574812 376964 574868 380072
rect 574812 376898 574868 376908
rect 575484 376852 575540 380072
rect 575484 376786 575540 376796
rect 576156 376628 576212 380072
rect 576156 376562 576212 376572
rect 574476 376450 574532 376460
rect 576828 376516 576884 380072
rect 577500 376628 577556 380072
rect 577500 376562 577556 376572
rect 576828 376450 576884 376460
rect 578172 376404 578228 380072
rect 578844 377860 578900 380072
rect 578844 377794 578900 377804
rect 579516 376516 579572 380072
rect 579516 376450 579572 376460
rect 578172 376338 578228 376348
rect 580188 375620 580244 380072
rect 580860 376740 580916 380072
rect 580860 376674 580916 376684
rect 581532 376516 581588 380072
rect 581532 376450 581588 376460
rect 582204 376292 582260 380072
rect 582204 376226 582260 376236
rect 580188 375554 580244 375564
rect 562716 66322 562772 66332
rect 575372 375508 575428 375518
rect 558684 63186 558740 63196
rect 566524 63812 566580 63822
rect 558572 60386 558628 60396
rect 561596 63140 561652 63150
rect 557340 59938 557396 59948
rect 561596 59864 561652 63084
rect 566524 59864 566580 63756
rect 575372 63140 575428 375452
rect 576380 311108 576436 311118
rect 575596 246148 575652 246158
rect 575596 63812 575652 246092
rect 575596 63746 575652 63756
rect 575372 63074 575428 63084
rect 571452 63028 571508 63038
rect 571452 59864 571508 62972
rect 576380 59864 576436 311052
rect 581308 140420 581364 140430
rect 581308 59864 581364 140364
rect 582876 140308 582932 380072
rect 583548 377636 583604 380072
rect 583548 377570 583604 377580
rect 584220 376516 584276 380072
rect 584892 377188 584948 380072
rect 584892 377122 584948 377132
rect 584220 376450 584276 376460
rect 585564 376516 585620 380072
rect 586236 376628 586292 380072
rect 586236 376562 586292 376572
rect 585564 376450 585620 376460
rect 586908 376516 586964 380072
rect 586908 376450 586964 376460
rect 588812 379764 588868 379774
rect 582876 140242 582932 140252
rect 587132 350756 587188 350766
rect 586236 63252 586292 63262
rect 586236 59864 586292 63196
rect 587132 63252 587188 350700
rect 587132 63186 587188 63196
rect 588028 66388 588084 66398
rect 588028 60228 588084 66332
rect 588812 63028 588868 379708
rect 590156 377188 590212 377198
rect 590156 375508 590212 377132
rect 590156 375442 590212 375452
rect 588924 297892 588980 297902
rect 588924 140420 588980 297836
rect 590492 246148 590548 430108
rect 590604 416836 590660 416846
rect 590604 379764 590660 416780
rect 590604 379698 590660 379708
rect 590716 390404 590772 390414
rect 590716 378868 590772 390348
rect 590716 378802 590772 378812
rect 590492 246082 590548 246092
rect 591164 337540 591220 337550
rect 588924 140354 588980 140364
rect 588812 62962 588868 62972
rect 588028 60162 588084 60172
rect 591164 59864 591220 337484
rect 554652 40674 554708 40684
rect 553980 20132 554148 20188
rect 554316 37604 554372 37614
rect 554316 36260 554372 37548
rect 553980 18340 554036 20132
rect 553980 18274 554036 18284
rect 552636 18050 552692 18060
rect 552188 16706 552244 16716
rect 553532 14308 553588 14318
rect 545132 9986 545188 9996
rect 551852 12628 551908 12638
rect 226940 9202 226996 9212
rect 551852 4340 551908 12572
rect 553532 4452 553588 14252
rect 554316 10836 554372 36204
rect 554316 10770 554372 10780
rect 557340 10612 557396 10622
rect 557340 10546 557396 10556
rect 560252 10612 560308 10622
rect 567196 10612 567252 10622
rect 560308 10556 560952 10612
rect 560252 10546 560308 10556
rect 567196 10546 567252 10556
rect 574588 10612 574644 10622
rect 586012 10612 586068 10622
rect 574644 10556 575288 10612
rect 559132 10500 559188 10510
rect 559132 10434 559188 10444
rect 565404 10500 565460 10510
rect 565404 10434 565460 10444
rect 560028 10388 560084 10398
rect 560028 10322 560084 10332
rect 574364 10388 574420 10398
rect 574420 10332 574532 10388
rect 574364 10322 574420 10332
rect 563612 10276 563668 10286
rect 574476 10276 574532 10332
rect 574392 10248 574532 10276
rect 563612 10210 563668 10220
rect 574364 10220 574532 10248
rect 557788 10164 557844 10174
rect 562716 10164 562772 10174
rect 556444 9828 556500 10136
rect 557844 10108 558264 10164
rect 561484 10108 561848 10164
rect 557788 10098 557844 10108
rect 561484 9940 561540 10108
rect 562716 10098 562772 10108
rect 561484 9874 561540 9884
rect 556444 7812 556500 9772
rect 564508 9716 564564 10136
rect 566328 10108 567140 10164
rect 569912 10136 570724 10164
rect 567084 9940 567140 10108
rect 567084 9874 567140 9884
rect 564508 9650 564564 9660
rect 556444 7746 556500 7756
rect 562940 9268 562996 9278
rect 553532 4386 553588 4396
rect 559468 7252 559524 7262
rect 551852 4274 551908 4284
rect 559468 4228 559524 7196
rect 559468 4162 559524 4172
rect 562940 4228 562996 9212
rect 568092 8372 568148 10136
rect 568092 8306 568148 8316
rect 568988 9716 569044 10136
rect 568988 8260 569044 9660
rect 569884 10108 570724 10136
rect 568988 8194 569044 8204
rect 569212 8260 569268 8270
rect 564396 7812 564452 7822
rect 564396 5012 564452 7756
rect 564396 4946 564452 4956
rect 566972 7364 567028 7374
rect 562940 4162 562996 4172
rect 566972 3108 567028 7308
rect 566972 3042 567028 3052
rect 567980 7028 568036 7038
rect 209356 392 209608 480
rect 211260 392 211512 480
rect 207480 -960 207704 392
rect 209384 -960 209608 392
rect 211288 -960 211512 392
rect 213192 -960 213416 480
rect 215096 -960 215320 480
rect 217000 -960 217224 480
rect 218904 -960 219128 480
rect 220808 -960 221032 480
rect 222712 -960 222936 480
rect 224616 -960 224840 480
rect 226520 -960 226744 480
rect 228424 -960 228648 480
rect 230328 -960 230552 480
rect 232232 -960 232456 480
rect 234136 -960 234360 480
rect 236040 -960 236264 480
rect 237944 -960 238168 480
rect 239848 -960 240072 480
rect 241752 -960 241976 480
rect 243656 -960 243880 480
rect 245560 -960 245784 480
rect 247464 -960 247688 480
rect 249368 -960 249592 480
rect 251272 -960 251496 480
rect 253176 -960 253400 480
rect 255080 -960 255304 480
rect 256984 -960 257208 480
rect 258888 -960 259112 480
rect 260792 -960 261016 480
rect 262696 -960 262920 480
rect 264600 -960 264824 480
rect 266504 -960 266728 480
rect 268408 -960 268632 480
rect 270312 -960 270536 480
rect 272216 -960 272440 480
rect 274120 -960 274344 480
rect 276024 -960 276248 480
rect 277928 -960 278152 480
rect 279832 -960 280056 480
rect 281736 -960 281960 480
rect 283640 -960 283864 480
rect 285544 -960 285768 480
rect 287448 -960 287672 480
rect 289352 -960 289576 480
rect 291256 -960 291480 480
rect 293160 -960 293384 480
rect 295064 -960 295288 480
rect 296968 -960 297192 480
rect 298872 -960 299096 480
rect 300776 -960 301000 480
rect 302680 -960 302904 480
rect 304584 -960 304808 480
rect 306488 -960 306712 480
rect 308392 -960 308616 480
rect 310296 -960 310520 480
rect 312200 -960 312424 480
rect 314104 -960 314328 480
rect 316008 -960 316232 480
rect 317912 -960 318136 480
rect 319816 -960 320040 480
rect 321720 -960 321944 480
rect 323624 -960 323848 480
rect 325528 -960 325752 480
rect 327432 -960 327656 480
rect 329336 -960 329560 480
rect 331240 -960 331464 480
rect 333144 -960 333368 480
rect 335048 -960 335272 480
rect 336952 -960 337176 480
rect 338856 -960 339080 480
rect 340760 -960 340984 480
rect 342664 -960 342888 480
rect 344568 -960 344792 480
rect 346472 -960 346696 480
rect 348376 -960 348600 480
rect 350280 -960 350504 480
rect 352184 -960 352408 480
rect 354088 -960 354312 480
rect 355992 -960 356216 480
rect 357896 -960 358120 480
rect 359800 -960 360024 480
rect 361704 -960 361928 480
rect 363608 -960 363832 480
rect 365512 -960 365736 480
rect 367416 -960 367640 480
rect 369320 -960 369544 480
rect 371224 -960 371448 480
rect 373128 -960 373352 480
rect 375032 -960 375256 480
rect 376936 -960 377160 480
rect 378840 -960 379064 480
rect 380744 -960 380968 480
rect 382648 -960 382872 480
rect 384552 -960 384776 480
rect 386456 -960 386680 480
rect 388360 -960 388584 480
rect 390264 -960 390488 480
rect 392168 -960 392392 480
rect 394072 -960 394296 480
rect 395976 -960 396200 480
rect 397880 -960 398104 480
rect 399784 -960 400008 480
rect 401688 -960 401912 480
rect 403592 -960 403816 480
rect 405496 -960 405720 480
rect 407400 -960 407624 480
rect 409304 -960 409528 480
rect 411208 -960 411432 480
rect 413112 -960 413336 480
rect 415016 -960 415240 480
rect 416920 -960 417144 480
rect 418824 -960 419048 480
rect 420728 -960 420952 480
rect 422632 -960 422856 480
rect 424536 -960 424760 480
rect 426440 -960 426664 480
rect 428344 -960 428568 480
rect 430248 -960 430472 480
rect 432152 -960 432376 480
rect 434056 -960 434280 480
rect 435960 -960 436184 480
rect 437864 -960 438088 480
rect 439768 -960 439992 480
rect 441672 -960 441896 480
rect 443576 -960 443800 480
rect 445480 -960 445704 480
rect 447384 -960 447608 480
rect 449288 -960 449512 480
rect 451192 -960 451416 480
rect 453096 -960 453320 480
rect 455000 -960 455224 480
rect 456904 -960 457128 480
rect 458808 -960 459032 480
rect 460712 -960 460936 480
rect 462616 -960 462840 480
rect 464520 -960 464744 480
rect 466424 -960 466648 480
rect 468328 -960 468552 480
rect 470232 -960 470456 480
rect 472136 -960 472360 480
rect 474040 -960 474264 480
rect 475944 -960 476168 480
rect 477848 -960 478072 480
rect 479752 -960 479976 480
rect 481656 -960 481880 480
rect 483560 -960 483784 480
rect 485464 -960 485688 480
rect 487368 -960 487592 480
rect 489272 -960 489496 480
rect 491176 -960 491400 480
rect 493080 -960 493304 480
rect 494984 -960 495208 480
rect 496888 -960 497112 480
rect 498792 -960 499016 480
rect 500696 -960 500920 480
rect 502600 -960 502824 480
rect 504504 -960 504728 480
rect 506408 -960 506632 480
rect 508312 -960 508536 480
rect 510216 -960 510440 480
rect 512120 -960 512344 480
rect 514024 -960 514248 480
rect 515928 -960 516152 480
rect 517832 -960 518056 480
rect 519736 -960 519960 480
rect 521640 -960 521864 480
rect 523544 -960 523768 480
rect 525448 -960 525672 480
rect 527352 -960 527576 480
rect 529256 -960 529480 480
rect 531160 -960 531384 480
rect 533064 -960 533288 480
rect 534968 -960 535192 480
rect 536872 -960 537096 480
rect 538776 -960 539000 480
rect 540680 -960 540904 480
rect 542584 -960 542808 480
rect 544488 -960 544712 480
rect 546392 -960 546616 480
rect 548296 -960 548520 480
rect 550200 -960 550424 480
rect 552104 -960 552328 480
rect 554008 -960 554232 480
rect 555912 -960 556136 480
rect 557816 -960 558040 480
rect 559720 -960 559944 480
rect 561624 -960 561848 480
rect 563528 -960 563752 480
rect 565432 -960 565656 480
rect 567336 -960 567560 480
rect 567980 420 568036 6972
rect 569212 6468 569268 8204
rect 569884 7588 569940 10108
rect 570668 9940 570724 10108
rect 570668 9874 570724 9884
rect 569884 7522 569940 7532
rect 570780 9268 570836 10136
rect 569212 6402 569268 6412
rect 570780 2548 570836 9212
rect 571676 9380 571732 10136
rect 571676 2660 571732 9324
rect 572572 9604 572628 10136
rect 572572 2772 572628 9548
rect 573468 9492 573524 10136
rect 573468 2884 573524 9436
rect 574364 2996 574420 10220
rect 574588 6916 574644 10556
rect 586012 10546 586068 10556
rect 591388 10612 591444 10622
rect 591388 10546 591444 10556
rect 575596 10500 575652 10510
rect 575652 10444 576184 10500
rect 575596 10434 575652 10444
rect 577052 8260 577108 10136
rect 577052 8194 577108 8204
rect 577948 8148 578004 10136
rect 577948 8082 578004 8092
rect 578844 8148 578900 10136
rect 579768 10108 579908 10164
rect 578844 8082 578900 8092
rect 579852 8148 579908 10108
rect 579852 8082 579908 8092
rect 580636 7924 580692 10136
rect 581532 8036 581588 10136
rect 582428 8260 582484 10136
rect 583324 8372 583380 10136
rect 583324 8306 583380 8316
rect 582428 8194 582484 8204
rect 581532 7970 581588 7980
rect 580636 7858 580692 7868
rect 578620 7700 578676 7710
rect 578620 7252 578676 7644
rect 578956 7364 579012 7374
rect 578620 7186 578676 7196
rect 578732 7308 578956 7364
rect 574588 6850 574644 6860
rect 574364 2930 574420 2940
rect 578732 6804 578788 7308
rect 578956 7298 579012 7308
rect 584220 7140 584276 10136
rect 585116 7700 585172 10136
rect 586908 9156 586964 10136
rect 586908 9090 586964 9100
rect 585116 7634 585172 7644
rect 587804 7252 587860 10136
rect 588700 7812 588756 10136
rect 588924 10108 589624 10164
rect 588924 10052 588980 10108
rect 588924 9986 588980 9996
rect 588700 7746 588756 7756
rect 590492 7364 590548 10136
rect 590492 7298 590548 7308
rect 587804 7186 587860 7196
rect 584220 7074 584276 7084
rect 573468 2818 573524 2828
rect 572572 2706 572628 2716
rect 571676 2594 571732 2604
rect 570780 2482 570836 2492
rect 578732 480 578788 6748
rect 582540 4452 582596 4462
rect 580636 4228 580692 4238
rect 580636 480 580692 4172
rect 582540 480 582596 4396
rect 584444 4340 584500 4350
rect 584444 480 584500 4284
rect 567980 354 568036 364
rect 569240 -960 569464 480
rect 571144 -960 571368 480
rect 573048 -960 573272 480
rect 574952 -960 575176 480
rect 576856 -960 577080 480
rect 578732 392 578984 480
rect 580636 392 580888 480
rect 582540 392 582792 480
rect 584444 392 584696 480
rect 578760 -960 578984 392
rect 580664 -960 580888 392
rect 582568 -960 582792 392
rect 584472 -960 584696 392
<< via2 >>
rect 11004 204092 11060 204148
rect 40908 590716 40964 590772
rect 40796 590604 40852 590660
rect 40684 590492 40740 590548
rect 40236 589596 40292 589652
rect 40796 225148 40852 225204
rect 40684 221340 40740 221396
rect 40236 209916 40292 209972
rect 33068 198492 33124 198548
rect 55132 590716 55188 590772
rect 77308 589708 77364 589764
rect 99260 589596 99316 589652
rect 41132 589484 41188 589540
rect 41020 589372 41076 589428
rect 41020 217532 41076 217588
rect 143388 590604 143444 590660
rect 165452 590492 165508 590548
rect 121324 589484 121380 589540
rect 187516 589372 187572 589428
rect 231756 590492 231812 590548
rect 298060 590604 298116 590660
rect 364252 590716 364308 590772
rect 430444 590828 430500 590884
rect 408380 589708 408436 589764
rect 496636 590940 496692 590996
rect 474572 589708 474628 589764
rect 540764 589708 540820 589764
rect 548828 590940 548884 590996
rect 342188 589596 342244 589652
rect 275996 589484 276052 589540
rect 209804 589372 209860 589428
rect 548716 589372 548772 589428
rect 43596 588812 43652 588868
rect 548828 583772 548884 583828
rect 550172 590828 550228 590884
rect 551852 590604 551908 590660
rect 551852 506492 551908 506548
rect 553532 590492 553588 590548
rect 550172 504812 550228 504868
rect 548716 503244 548772 503300
rect 562716 590492 562772 590548
rect 575372 590716 575428 590772
rect 563612 589596 563668 589652
rect 553532 503132 553588 503188
rect 560252 589484 560308 589540
rect 570332 589036 570388 589092
rect 568540 588924 568596 588980
rect 566748 588812 566804 588868
rect 563612 503916 563668 503972
rect 564956 503916 565012 503972
rect 560252 502684 560308 502740
rect 561372 503244 561428 503300
rect 563164 502684 563220 502740
rect 572124 588588 572180 588644
rect 573916 548940 573972 548996
rect 584668 590492 584724 590548
rect 582876 583772 582932 583828
rect 575372 503916 575428 503972
rect 577500 506492 577556 506548
rect 575708 503132 575764 503188
rect 581084 504812 581140 504868
rect 579292 503916 579348 503972
rect 586460 575372 586516 575428
rect 588252 535724 588308 535780
rect 551852 492268 551908 492324
rect 550172 449260 550228 449316
rect 221564 232652 221620 232708
rect 207228 232540 207284 232596
rect 200060 232428 200116 232484
rect 71036 232204 71092 232260
rect 135548 232092 135604 232148
rect 106876 230748 106932 230804
rect 85372 230412 85428 230468
rect 114044 230636 114100 230692
rect 171388 230524 171444 230580
rect 149884 230188 149940 230244
rect 157052 229852 157108 229908
rect 185724 230300 185780 230356
rect 179228 229964 179284 230020
rect 214396 232316 214452 232372
rect 242956 232652 243012 232708
rect 228732 231980 228788 232036
rect 240156 231980 240212 232036
rect 235900 231868 235956 231924
rect 121212 229740 121268 229796
rect 92540 229628 92596 229684
rect 164220 229516 164276 229572
rect 78652 229404 78708 229460
rect 128380 229404 128436 229460
rect 63868 229292 63924 229348
rect 192892 229292 192948 229348
rect 242732 231868 242788 231924
rect 240156 224252 240212 224308
rect 241948 229628 242004 229684
rect 241948 222684 242004 222740
rect 549388 232428 549444 232484
rect 247772 232316 247828 232372
rect 243628 232204 243684 232260
rect 246876 230748 246932 230804
rect 243628 224476 243684 224532
rect 244412 229740 244468 229796
rect 242956 217644 243012 217700
rect 242732 217532 242788 217588
rect 43596 213724 43652 213780
rect 41132 206108 41188 206164
rect 53788 204092 53844 204148
rect 53788 202300 53844 202356
rect 40908 194684 40964 194740
rect 246876 222572 246932 222628
rect 315868 232092 315924 232148
rect 247772 219436 247828 219492
rect 289884 230636 289940 230692
rect 244412 172172 244468 172228
rect 409836 230524 409892 230580
rect 391916 230412 391972 230468
rect 375340 227836 375396 227892
rect 315868 224364 315924 224420
rect 358764 224476 358820 224532
rect 408492 222684 408548 222740
rect 505148 230300 505204 230356
rect 474796 230188 474852 230244
rect 456764 229852 456820 229908
rect 424956 227612 425012 227668
rect 409836 222684 409892 222740
rect 456764 223356 456820 223412
rect 458220 223356 458276 223412
rect 441644 222572 441700 222628
rect 491372 229516 491428 229572
rect 524076 229964 524132 230020
rect 505148 223356 505204 223412
rect 507948 223356 508004 223412
rect 541100 222684 541156 222740
rect 347228 219660 347284 219716
rect 343532 215852 343588 215908
rect 309820 172172 309876 172228
rect 289772 65548 289828 65604
rect 242844 52892 242900 52948
rect 239372 51548 239428 51604
rect 242732 49196 242788 49252
rect 240268 39452 240324 39508
rect 240156 34412 240212 34468
rect 241948 37772 242004 37828
rect 241388 37212 241444 37268
rect 241164 37100 241220 37156
rect 240268 32508 240324 32564
rect 241052 36092 241108 36148
rect 240156 31276 240212 31332
rect 239372 31052 239428 31108
rect 139132 30716 139188 30772
rect 140924 30716 140980 30772
rect 142716 30716 142772 30772
rect 149884 30716 149940 30772
rect 137340 30604 137396 30660
rect 151676 30604 151732 30660
rect 153468 30604 153524 30660
rect 158844 30604 158900 30660
rect 160636 30604 160692 30660
rect 162428 30604 162484 30660
rect 185724 30604 185780 30660
rect 191100 30604 191156 30660
rect 196476 30604 196532 30660
rect 135548 30380 135604 30436
rect 105084 30268 105140 30324
rect 134428 30268 134484 30324
rect 96124 30156 96180 30212
rect 69692 26908 69748 26964
rect 58940 26572 58996 26628
rect 45612 26460 45668 26516
rect 13244 26012 13300 26068
rect 11340 12572 11396 12628
rect 27692 24444 27748 24500
rect 18956 19404 19012 19460
rect 15148 14252 15204 14308
rect 17276 6524 17332 6580
rect 22764 17836 22820 17892
rect 21980 7532 22036 7588
rect 24892 4284 24948 4340
rect 27692 4284 27748 4340
rect 27916 24332 27972 24388
rect 26796 4172 26852 4228
rect 41804 21196 41860 21252
rect 37996 19628 38052 19684
rect 32284 19292 32340 19348
rect 30380 16156 30436 16212
rect 27916 4172 27972 4228
rect 28700 7644 28756 7700
rect 34412 10892 34468 10948
rect 36316 9324 36372 9380
rect 41132 16044 41188 16100
rect 40124 4172 40180 4228
rect 41132 4172 41188 4228
rect 43932 5852 43988 5908
rect 53228 24668 53284 24724
rect 47516 17612 47572 17668
rect 49420 14364 49476 14420
rect 51548 7756 51604 7812
rect 55132 21308 55188 21364
rect 57260 4172 57316 4228
rect 66556 24556 66612 24612
rect 62748 15932 62804 15988
rect 59612 12684 59668 12740
rect 59612 4172 59668 4228
rect 61068 4172 61124 4228
rect 62972 14476 63028 14532
rect 62972 4172 63028 4228
rect 64652 12908 64708 12964
rect 68460 17724 68516 17780
rect 72828 26908 72884 26964
rect 69692 12572 69748 12628
rect 72268 26236 72324 26292
rect 70476 5964 70532 6020
rect 74620 26012 74676 26068
rect 77980 25900 78036 25956
rect 76300 6076 76356 6132
rect 74396 4956 74452 5012
rect 78204 21644 78260 21700
rect 81788 30044 81844 30100
rect 81788 27356 81844 27412
rect 79212 19404 79268 19460
rect 79212 9996 79268 10052
rect 81452 19404 81508 19460
rect 83580 7532 83636 7588
rect 83692 19516 83748 19572
rect 81452 4956 81508 5012
rect 82012 6748 82068 6804
rect 80108 4172 80164 4228
rect 86492 13356 86548 13412
rect 85372 8204 85428 8260
rect 85372 6748 85428 6804
rect 85820 9212 85876 9268
rect 87164 13356 87220 13412
rect 88956 30044 89012 30100
rect 86492 6076 86548 6132
rect 87500 7532 87556 7588
rect 90748 28364 90804 28420
rect 91532 28364 91588 28420
rect 91308 26124 91364 26180
rect 89852 24220 89908 24276
rect 88956 5964 89012 6020
rect 89404 12796 89460 12852
rect 89852 4172 89908 4228
rect 92540 28140 92596 28196
rect 92540 26572 92596 26628
rect 94332 29820 94388 29876
rect 96124 26460 96180 26516
rect 97916 29820 97972 29876
rect 94332 24668 94388 24724
rect 95116 26012 95172 26068
rect 91532 12908 91588 12964
rect 93436 2492 93492 2548
rect 97916 19628 97972 19684
rect 99708 23436 99764 23492
rect 101500 24780 101556 24836
rect 99708 16156 99764 16212
rect 100828 17948 100884 18004
rect 97020 12572 97076 12628
rect 99036 2604 99092 2660
rect 101500 17836 101556 17892
rect 105084 27356 105140 27412
rect 106652 28252 106708 28308
rect 103292 18396 103348 18452
rect 102732 16156 102788 16212
rect 103292 7756 103348 7812
rect 106540 16268 106596 16324
rect 104860 2716 104916 2772
rect 106652 9324 106708 9380
rect 110460 28476 110516 28532
rect 112252 28476 112308 28532
rect 112588 28700 112644 28756
rect 112588 28140 112644 28196
rect 117516 29372 117572 29428
rect 117516 28252 117572 28308
rect 115836 27804 115892 27860
rect 114044 27692 114100 27748
rect 117628 27580 117684 27636
rect 124796 28140 124852 28196
rect 123004 28028 123060 28084
rect 121212 27468 121268 27524
rect 119420 22652 119476 22708
rect 108332 20076 108388 20132
rect 125580 21532 125636 21588
rect 117964 19740 118020 19796
rect 114380 9436 114436 9492
rect 108332 7644 108388 7700
rect 108668 9324 108724 9380
rect 112476 6188 112532 6244
rect 110572 2828 110628 2884
rect 116284 2940 116340 2996
rect 119868 17836 119924 17892
rect 123676 13020 123732 13076
rect 121996 5852 122052 5908
rect 126588 21084 126644 21140
rect 128380 20972 128436 21028
rect 129388 26908 129444 26964
rect 127596 5964 127652 6020
rect 131964 28476 132020 28532
rect 198268 30604 198324 30660
rect 200060 30604 200116 30660
rect 135548 26908 135604 26964
rect 130172 26460 130228 26516
rect 131292 19628 131348 19684
rect 133420 6076 133476 6132
rect 137340 13020 137396 13076
rect 140812 28364 140868 28420
rect 137004 12908 137060 12964
rect 147868 29708 147924 29764
rect 147868 26908 147924 26964
rect 146300 26684 146356 26740
rect 146188 26460 146244 26516
rect 148428 26348 148484 26404
rect 146188 26012 146244 26068
rect 146524 26012 146580 26068
rect 144508 24892 144564 24948
rect 145292 24892 145348 24948
rect 145292 17948 145348 18004
rect 142828 14588 142884 14644
rect 139244 28 139300 84
rect 155260 28252 155316 28308
rect 157052 29708 157108 29764
rect 158844 27916 158900 27972
rect 160636 27356 160692 27412
rect 162428 27356 162484 27412
rect 163660 28140 163716 28196
rect 156268 26908 156324 26964
rect 153468 26236 153524 26292
rect 151676 25900 151732 25956
rect 159852 25228 159908 25284
rect 157948 21084 158004 21140
rect 152236 20972 152292 21028
rect 144956 140 145012 196
rect 154140 17948 154196 18004
rect 156156 6188 156212 6244
rect 163660 24668 163716 24724
rect 150668 252 150724 308
rect 163884 25004 163940 25060
rect 167804 28140 167860 28196
rect 166012 25116 166068 25172
rect 166012 24444 166068 24500
rect 169372 28028 169428 28084
rect 163884 19292 163940 19348
rect 173180 28364 173236 28420
rect 171388 28252 171444 28308
rect 169596 28028 169652 28084
rect 174972 27916 175028 27972
rect 175084 27468 175140 27524
rect 169372 21756 169428 21812
rect 165788 7644 165844 7700
rect 167692 6300 167748 6356
rect 162652 364 162708 420
rect 171388 25340 171444 25396
rect 174636 7756 174692 7812
rect 174636 6524 174692 6580
rect 173404 6412 173460 6468
rect 176316 27468 176372 27524
rect 176316 26572 176372 26628
rect 176764 17612 176820 17668
rect 176988 23324 177044 23380
rect 178556 23324 178612 23380
rect 180348 25340 180404 25396
rect 180348 22988 180404 23044
rect 176988 17500 177044 17556
rect 180796 22652 180852 22708
rect 179116 3052 179172 3108
rect 183148 25228 183204 25284
rect 183148 24556 183204 24612
rect 182252 20860 182308 20916
rect 186284 27916 186340 27972
rect 186284 27468 186340 27524
rect 186508 27916 186564 27972
rect 186508 27580 186564 27636
rect 185724 17948 185780 18004
rect 182252 7644 182308 7700
rect 182700 17612 182756 17668
rect 184828 7644 184884 7700
rect 187516 26348 187572 26404
rect 188412 29708 188468 29764
rect 188412 27468 188468 27524
rect 189308 23212 189364 23268
rect 189308 14588 189364 14644
rect 190316 12908 190372 12964
rect 192220 27916 192276 27972
rect 190540 7868 190596 7924
rect 192332 24444 192388 24500
rect 194124 28476 194180 28532
rect 192892 24444 192948 24500
rect 193228 26236 193284 26292
rect 193228 21532 193284 21588
rect 192332 19628 192388 19684
rect 194684 26236 194740 26292
rect 196476 17836 196532 17892
rect 198156 27692 198212 27748
rect 198156 26460 198212 26516
rect 198268 9436 198324 9492
rect 199948 16828 200004 16884
rect 196252 7980 196308 8036
rect 203532 29708 203588 29764
rect 201852 28476 201908 28532
rect 202412 28476 202468 28532
rect 200732 28252 200788 28308
rect 200732 18172 200788 18228
rect 200732 16828 200788 16884
rect 202412 16156 202468 16212
rect 205436 29484 205492 29540
rect 203532 12572 203588 12628
rect 203644 27580 203700 27636
rect 200060 9324 200116 9380
rect 201964 4172 202020 4228
rect 205436 26124 205492 26180
rect 205548 28028 205604 28084
rect 207452 27356 207508 27412
rect 209020 27804 209076 27860
rect 209020 24220 209076 24276
rect 210812 28364 210868 28420
rect 207452 9212 207508 9268
rect 209356 21532 209412 21588
rect 207676 4284 207732 4340
rect 212492 28252 212548 28308
rect 210812 19404 210868 19460
rect 211260 28140 211316 28196
rect 211260 18060 211316 18116
rect 212492 17724 212548 17780
rect 215852 28476 215908 28532
rect 214172 28140 214228 28196
rect 214172 15932 214228 15988
rect 221564 29596 221620 29652
rect 219884 28476 219940 28532
rect 217532 27692 217588 27748
rect 223356 26124 223412 26180
rect 223356 24332 223412 24388
rect 225932 24332 225988 24388
rect 217532 14364 217588 14420
rect 225932 14252 225988 14308
rect 228732 14252 228788 14308
rect 241500 36204 241556 36260
rect 241948 32844 242004 32900
rect 241500 31164 241556 31220
rect 241388 30156 241444 30212
rect 241164 29820 241220 29876
rect 242844 32396 242900 32452
rect 242956 42812 243012 42868
rect 242956 30716 243012 30772
rect 243068 37324 243124 37380
rect 243068 29932 243124 29988
rect 242732 28028 242788 28084
rect 241052 27916 241108 27972
rect 309820 26796 309876 26852
rect 343420 53900 343476 53956
rect 289772 21644 289828 21700
rect 343644 210028 343700 210084
rect 347564 219548 347620 219604
rect 347340 216860 347396 216916
rect 347340 205772 347396 205828
rect 347452 216748 347508 216804
rect 347452 199724 347508 199780
rect 347676 216972 347732 217028
rect 347676 210028 347732 210084
rect 347564 194348 347620 194404
rect 347228 188972 347284 189028
rect 549388 184380 549444 184436
rect 344316 156716 344372 156772
rect 344204 151340 344260 151396
rect 344092 145964 344148 146020
rect 343980 140588 344036 140644
rect 343868 135212 343924 135268
rect 343756 129836 343812 129892
rect 343756 36204 343812 36260
rect 343756 35532 343812 35588
rect 343868 34188 343924 34244
rect 343756 32844 343812 32900
rect 343756 32620 343812 32676
rect 347004 108332 347060 108388
rect 346780 97580 346836 97636
rect 346668 70700 346724 70756
rect 346108 53788 346164 53844
rect 346108 52892 346164 52948
rect 346668 51884 346724 51940
rect 346780 42812 346836 42868
rect 347452 92204 347508 92260
rect 347340 86828 347396 86884
rect 347228 81452 347284 81508
rect 347116 76076 347172 76132
rect 347116 51996 347172 52052
rect 347228 50316 347284 50372
rect 347340 48412 347396 48468
rect 347564 65324 347620 65380
rect 347676 59948 347732 60004
rect 347676 53788 347732 53844
rect 350364 53788 350420 53844
rect 349804 51884 349860 51940
rect 347564 51548 347620 51604
rect 349580 51548 349636 51604
rect 347452 45388 347508 45444
rect 347004 40908 347060 40964
rect 344092 31500 344148 31556
rect 344316 30156 344372 30212
rect 344316 29708 344372 29764
rect 344204 29484 344260 29540
rect 344204 28812 344260 28868
rect 343644 26124 343700 26180
rect 346108 27804 346164 27860
rect 346108 26124 346164 26180
rect 343532 24332 343588 24388
rect 343420 18172 343476 18228
rect 347004 23212 347060 23268
rect 349692 50316 349748 50372
rect 349692 35084 349748 35140
rect 349580 21420 349636 21476
rect 349692 21308 349748 21364
rect 350140 48748 350196 48804
rect 350028 43596 350084 43652
rect 350140 23324 350196 23380
rect 550060 53004 550116 53060
rect 549388 45500 549444 45556
rect 431788 40684 431844 40740
rect 472108 40684 472164 40740
rect 443884 40572 443940 40628
rect 444108 40572 444164 40628
rect 436268 40460 436324 40516
rect 359212 37772 359268 37828
rect 354508 37660 354564 37716
rect 350364 23212 350420 23268
rect 350812 35084 350868 35140
rect 349804 23100 349860 23156
rect 346892 18060 346948 18116
rect 350812 22988 350868 23044
rect 349804 17612 349860 17668
rect 230524 12572 230580 12628
rect 362908 36988 362964 37044
rect 367052 37436 367108 37492
rect 367052 30044 367108 30100
rect 378812 37324 378868 37380
rect 383852 37212 383908 37268
rect 383852 36988 383908 37044
rect 387436 37100 387492 37156
rect 378812 30044 378868 30100
rect 375340 28700 375396 28756
rect 376236 28700 376292 28756
rect 371308 28588 371364 28644
rect 376236 26348 376292 26404
rect 387212 25788 387268 25844
rect 391468 25900 391524 25956
rect 394828 29596 394884 29652
rect 394828 24780 394884 24836
rect 391468 23436 391524 23492
rect 403564 32956 403620 33012
rect 407596 29372 407652 29428
rect 415660 40012 415716 40068
rect 419692 39676 419748 39732
rect 427756 39788 427812 39844
rect 427756 36092 427812 36148
rect 423388 35308 423444 35364
rect 423388 26460 423444 26516
rect 439852 40124 439908 40180
rect 455980 40460 456036 40516
rect 456204 40460 456260 40516
rect 447916 39788 447972 39844
rect 439852 26572 439908 26628
rect 435148 22652 435204 22708
rect 447916 24668 447972 24724
rect 451948 39452 452004 39508
rect 443884 21756 443940 21812
rect 415660 21532 415716 21588
rect 464044 40348 464100 40404
rect 460012 39340 460068 39396
rect 463708 37324 463764 37380
rect 468076 40236 468132 40292
rect 451948 21084 452004 21140
rect 476140 39228 476196 39284
rect 480172 39676 480228 39732
rect 480172 37660 480228 37716
rect 483868 39676 483924 39732
rect 483868 37660 483924 37716
rect 488236 39676 488292 39732
rect 488236 37660 488292 37716
rect 492268 39452 492324 39508
rect 476140 30492 476196 30548
rect 472108 30380 472164 30436
rect 468076 30268 468132 30324
rect 458668 26012 458724 26068
rect 496300 39676 496356 39732
rect 500332 38108 500388 38164
rect 500332 36988 500388 37044
rect 504812 38444 504868 38500
rect 504812 36988 504868 37044
rect 508396 38332 508452 38388
rect 516460 39676 516516 39732
rect 512428 39340 512484 39396
rect 512428 36988 512484 37044
rect 524524 38556 524580 38612
rect 532588 39676 532644 39732
rect 532588 37996 532644 38052
rect 528556 36988 528612 37044
rect 536732 37884 536788 37940
rect 540092 37996 540148 38052
rect 520716 34524 520772 34580
rect 508396 32732 508452 32788
rect 496300 26684 496356 26740
rect 540092 25116 540148 25172
rect 549388 36428 549444 36484
rect 545132 26796 545188 26852
rect 536732 25004 536788 25060
rect 492268 24892 492324 24948
rect 455980 20972 456036 21028
rect 411628 20076 411684 20132
rect 399532 18396 399588 18452
rect 362908 13356 362964 13412
rect 354508 9996 354564 10052
rect 550172 40572 550228 40628
rect 550284 433132 550340 433188
rect 550396 422380 550452 422436
rect 550620 414316 550676 414372
rect 550396 41356 550452 41412
rect 550508 398188 550564 398244
rect 550284 40236 550340 40292
rect 550620 41468 550676 41524
rect 550732 403564 550788 403620
rect 551404 60284 551460 60340
rect 550956 60172 551012 60228
rect 550732 39340 550788 39396
rect 550844 55692 550900 55748
rect 550508 34524 550564 34580
rect 550956 38444 551012 38500
rect 551740 44940 551796 44996
rect 551740 34860 551796 34916
rect 556892 489580 556948 489636
rect 553644 473452 553700 473508
rect 551964 468076 552020 468132
rect 553532 435820 553588 435876
rect 551964 40012 552020 40068
rect 552076 411628 552132 411684
rect 552076 38108 552132 38164
rect 552188 393148 552244 393204
rect 552188 216860 552244 216916
rect 551628 28252 551684 28308
rect 550844 23324 550900 23380
rect 551516 27020 551572 27076
rect 550060 23212 550116 23268
rect 551740 28364 551796 28420
rect 551740 24780 551796 24836
rect 551964 28476 552020 28532
rect 551628 23436 551684 23492
rect 551964 22092 552020 22148
rect 551516 20748 551572 20804
rect 552300 232540 552356 232596
rect 553196 227724 553252 227780
rect 552972 224252 553028 224308
rect 552860 217532 552916 217588
rect 552748 193900 552804 193956
rect 553084 219436 553140 219492
rect 553084 203756 553140 203812
rect 552972 174188 553028 174244
rect 552860 164332 552916 164388
rect 553196 154476 553252 154532
rect 552524 60396 552580 60452
rect 552412 47628 552468 47684
rect 552300 46284 552356 46340
rect 552412 35084 552468 35140
rect 552300 33516 552356 33572
rect 555212 470764 555268 470820
rect 553644 226828 553700 226884
rect 553756 446572 553812 446628
rect 553532 40348 553588 40404
rect 554652 430444 554708 430500
rect 553868 425068 553924 425124
rect 553868 41132 553924 41188
rect 553980 417004 554036 417060
rect 553756 39788 553812 39844
rect 553980 39452 554036 39508
rect 554092 56476 554148 56532
rect 552524 28476 552580 28532
rect 552300 27692 552356 27748
rect 552300 19404 552356 19460
rect 552636 26908 552692 26964
rect 555212 216524 555268 216580
rect 556108 218428 556164 218484
rect 556220 216748 556276 216804
rect 556220 199836 556276 199892
rect 556108 193228 556164 193284
rect 556668 63196 556724 63252
rect 558572 486892 558628 486948
rect 557676 484204 557732 484260
rect 557004 481516 557060 481572
rect 557228 478828 557284 478884
rect 557004 219548 557060 219604
rect 557004 218428 557060 218484
rect 557116 408940 557172 408996
rect 556892 60284 556948 60340
rect 557452 476140 557508 476196
rect 557228 216748 557284 216804
rect 557340 406252 557396 406308
rect 557116 60172 557172 60228
rect 557452 393148 557508 393204
rect 557676 379708 557732 379764
rect 590492 430108 590548 430164
rect 559468 379708 559524 379764
rect 558684 378812 558740 378868
rect 559468 219660 559524 219716
rect 559468 189756 559524 189812
rect 564060 377468 564116 377524
rect 566076 377356 566132 377412
rect 565404 377244 565460 377300
rect 564732 376796 564788 376852
rect 567420 377356 567476 377412
rect 568092 377244 568148 377300
rect 568764 376684 568820 376740
rect 566748 376572 566804 376628
rect 563388 376460 563444 376516
rect 570108 376572 570164 376628
rect 569436 376460 569492 376516
rect 571452 376572 571508 376628
rect 571004 376460 571060 376516
rect 572572 376460 572628 376516
rect 573468 376572 573524 376628
rect 572796 376460 572852 376516
rect 574812 376908 574868 376964
rect 575484 376796 575540 376852
rect 576156 376572 576212 376628
rect 574476 376460 574532 376516
rect 577500 376572 577556 376628
rect 576828 376460 576884 376516
rect 578844 377804 578900 377860
rect 579516 376460 579572 376516
rect 578172 376348 578228 376404
rect 580860 376684 580916 376740
rect 581532 376460 581588 376516
rect 582204 376236 582260 376292
rect 580188 375564 580244 375620
rect 562716 66332 562772 66388
rect 575372 375452 575428 375508
rect 558684 63196 558740 63252
rect 566524 63756 566580 63812
rect 558572 60396 558628 60452
rect 561596 63084 561652 63140
rect 557340 59948 557396 60004
rect 576380 311052 576436 311108
rect 575596 246092 575652 246148
rect 575596 63756 575652 63812
rect 575372 63084 575428 63140
rect 571452 62972 571508 63028
rect 581308 140364 581364 140420
rect 583548 377580 583604 377636
rect 584892 377132 584948 377188
rect 584220 376460 584276 376516
rect 586236 376572 586292 376628
rect 585564 376460 585620 376516
rect 586908 376460 586964 376516
rect 588812 379708 588868 379764
rect 582876 140252 582932 140308
rect 587132 350700 587188 350756
rect 586236 63196 586292 63252
rect 587132 63196 587188 63252
rect 588028 66332 588084 66388
rect 590156 377132 590212 377188
rect 590156 375452 590212 375508
rect 588924 297836 588980 297892
rect 590604 416780 590660 416836
rect 590604 379708 590660 379764
rect 590716 390348 590772 390404
rect 590716 378812 590772 378868
rect 590492 246092 590548 246148
rect 591164 337484 591220 337540
rect 588924 140364 588980 140420
rect 588812 62972 588868 63028
rect 588028 60172 588084 60228
rect 554652 40684 554708 40740
rect 554316 37548 554372 37604
rect 554316 36204 554372 36260
rect 553980 18284 554036 18340
rect 552636 18060 552692 18116
rect 552188 16716 552244 16772
rect 553532 14252 553588 14308
rect 545132 9996 545188 10052
rect 551852 12572 551908 12628
rect 226940 9212 226996 9268
rect 554316 10780 554372 10836
rect 557340 10556 557396 10612
rect 560252 10556 560308 10612
rect 567196 10556 567252 10612
rect 574588 10556 574644 10612
rect 586012 10556 586068 10612
rect 559132 10444 559188 10500
rect 565404 10444 565460 10500
rect 560028 10332 560084 10388
rect 574364 10332 574420 10388
rect 563612 10220 563668 10276
rect 557788 10108 557844 10164
rect 562716 10108 562772 10164
rect 561484 9884 561540 9940
rect 556444 9772 556500 9828
rect 567084 9884 567140 9940
rect 564508 9660 564564 9716
rect 556444 7756 556500 7812
rect 562940 9212 562996 9268
rect 553532 4396 553588 4452
rect 559468 7196 559524 7252
rect 551852 4284 551908 4340
rect 559468 4172 559524 4228
rect 568092 8316 568148 8372
rect 568988 9660 569044 9716
rect 568988 8204 569044 8260
rect 569212 8204 569268 8260
rect 564396 7756 564452 7812
rect 564396 4956 564452 5012
rect 566972 7308 567028 7364
rect 562940 4172 562996 4228
rect 566972 3052 567028 3108
rect 567980 6972 568036 7028
rect 570668 9884 570724 9940
rect 569884 7532 569940 7588
rect 570780 9212 570836 9268
rect 569212 6412 569268 6468
rect 571676 9324 571732 9380
rect 572572 9548 572628 9604
rect 573468 9436 573524 9492
rect 591388 10556 591444 10612
rect 575596 10444 575652 10500
rect 577052 8204 577108 8260
rect 577948 8092 578004 8148
rect 578844 8092 578900 8148
rect 579852 8092 579908 8148
rect 583324 8316 583380 8372
rect 582428 8204 582484 8260
rect 581532 7980 581588 8036
rect 580636 7868 580692 7924
rect 578620 7644 578676 7700
rect 578620 7196 578676 7252
rect 578956 7308 579012 7364
rect 574588 6860 574644 6916
rect 574364 2940 574420 2996
rect 586908 9100 586964 9156
rect 585116 7644 585172 7700
rect 588924 9996 588980 10052
rect 588700 7756 588756 7812
rect 590492 7308 590548 7364
rect 587804 7196 587860 7252
rect 584220 7084 584276 7140
rect 578732 6748 578788 6804
rect 573468 2828 573524 2884
rect 572572 2716 572628 2772
rect 571676 2604 571732 2660
rect 570780 2492 570836 2548
rect 582540 4396 582596 4452
rect 580636 4172 580692 4228
rect 584444 4284 584500 4340
rect 567980 364 568036 420
<< metal3 >>
rect 496626 590940 496636 590996
rect 496692 590940 548828 590996
rect 548884 590940 548894 590996
rect 430434 590828 430444 590884
rect 430500 590828 550172 590884
rect 550228 590828 550238 590884
rect 40898 590716 40908 590772
rect 40964 590716 55132 590772
rect 55188 590716 55198 590772
rect 364242 590716 364252 590772
rect 364308 590716 575372 590772
rect 575428 590716 575438 590772
rect 40786 590604 40796 590660
rect 40852 590604 143388 590660
rect 143444 590604 143454 590660
rect 298050 590604 298060 590660
rect 298116 590604 551852 590660
rect 551908 590604 551918 590660
rect 40674 590492 40684 590548
rect 40740 590492 165452 590548
rect 165508 590492 165518 590548
rect 231746 590492 231756 590548
rect 231812 590492 553532 590548
rect 553588 590492 553598 590548
rect 562706 590492 562716 590548
rect 562772 590492 584668 590548
rect 584724 590492 584734 590548
rect 77270 589708 77308 589764
rect 77364 589708 77374 589764
rect 408342 589708 408380 589764
rect 408436 589708 408446 589764
rect 474534 589708 474572 589764
rect 474628 589708 474638 589764
rect 540726 589708 540764 589764
rect 540820 589708 540830 589764
rect 40226 589596 40236 589652
rect 40292 589596 99260 589652
rect 99316 589596 99326 589652
rect 342178 589596 342188 589652
rect 342244 589596 563612 589652
rect 563668 589596 563678 589652
rect 41122 589484 41132 589540
rect 41188 589484 121324 589540
rect 121380 589484 121390 589540
rect 275986 589484 275996 589540
rect 276052 589484 560252 589540
rect 560308 589484 560318 589540
rect 41010 589372 41020 589428
rect 41076 589372 187516 589428
rect 187572 589372 187582 589428
rect 209794 589372 209804 589428
rect 209860 589372 548716 589428
rect 548772 589372 548782 589428
rect 474562 589260 474572 589316
rect 474628 589260 478828 589316
rect 540754 589260 540764 589316
rect 540820 589260 549388 589316
rect 478772 588980 478828 589260
rect 549332 589092 549388 589260
rect 549332 589036 570332 589092
rect 570388 589036 570398 589092
rect 478772 588924 568540 588980
rect 568596 588924 568606 588980
rect 43586 588812 43596 588868
rect 43652 588812 77308 588868
rect 77364 588812 77374 588868
rect 408370 588812 408380 588868
rect 408436 588812 566748 588868
rect 566804 588812 566814 588868
rect 595560 588644 597000 588840
rect 572114 588588 572124 588644
rect 572180 588616 597000 588644
rect 572180 588588 595672 588616
rect -960 587188 480 587384
rect -960 587160 37772 587188
rect 392 587132 37772 587160
rect 37828 587132 37838 587188
rect 548818 583772 548828 583828
rect 548884 583772 582876 583828
rect 582932 583772 582942 583828
rect 595560 575428 597000 575624
rect 586450 575372 586460 575428
rect 586516 575400 597000 575428
rect 586516 575372 595672 575400
rect -960 573076 480 573272
rect -960 573048 27692 573076
rect 392 573020 27692 573048
rect 27748 573020 27758 573076
rect 595560 562184 597000 562408
rect -960 558964 480 559160
rect -960 558936 36092 558964
rect 392 558908 36092 558936
rect 36148 558908 36158 558964
rect 595560 548996 597000 549192
rect 573906 548940 573916 548996
rect 573972 548968 597000 548996
rect 573972 548940 595672 548968
rect -960 544852 480 545048
rect -960 544824 5852 544852
rect 392 544796 5852 544824
rect 5908 544796 5918 544852
rect 595560 535780 597000 535976
rect 588242 535724 588252 535780
rect 588308 535752 597000 535780
rect 588308 535724 595672 535752
rect -960 530740 480 530936
rect -960 530712 22652 530740
rect 392 530684 22652 530712
rect 22708 530684 22718 530740
rect 595560 522536 597000 522760
rect -960 516628 480 516824
rect -960 516600 34412 516628
rect 392 516572 34412 516600
rect 34468 516572 34478 516628
rect 595560 509320 597000 509544
rect 551842 506492 551852 506548
rect 551908 506492 577500 506548
rect 577556 506492 577566 506548
rect 550162 504812 550172 504868
rect 550228 504812 581084 504868
rect 581140 504812 581150 504868
rect 563602 503916 563612 503972
rect 563668 503916 564956 503972
rect 565012 503916 565022 503972
rect 575362 503916 575372 503972
rect 575428 503916 579292 503972
rect 579348 503916 579358 503972
rect 548706 503244 548716 503300
rect 548772 503244 561372 503300
rect 561428 503244 561438 503300
rect 553522 503132 553532 503188
rect 553588 503132 575708 503188
rect 575764 503132 575774 503188
rect -960 502516 480 502712
rect 560242 502684 560252 502740
rect 560308 502684 563164 502740
rect 563220 502684 563230 502740
rect -960 502488 12572 502516
rect 392 502460 12572 502488
rect 12628 502460 12638 502516
rect 595560 496104 597000 496328
rect 551842 492268 551852 492324
rect 551908 492268 560056 492324
rect 556882 489580 556892 489636
rect 556948 489580 560056 489636
rect -960 488404 480 488600
rect -960 488376 4172 488404
rect 392 488348 4172 488376
rect 4228 488348 4238 488404
rect 558562 486892 558572 486948
rect 558628 486892 560056 486948
rect 557666 484204 557676 484260
rect 557732 484204 560056 484260
rect 595560 482888 597000 483112
rect 556994 481516 557004 481572
rect 557060 481516 560056 481572
rect 557218 478828 557228 478884
rect 557284 478828 560056 478884
rect 557442 476140 557452 476196
rect 557508 476140 560056 476196
rect -960 474292 480 474488
rect -960 474264 5964 474292
rect 392 474236 5964 474264
rect 6020 474236 6030 474292
rect 553634 473452 553644 473508
rect 553700 473452 560056 473508
rect 555202 470764 555212 470820
rect 555268 470764 560056 470820
rect 595560 469672 597000 469896
rect 551954 468076 551964 468132
rect 552020 468076 560056 468132
rect 560242 465388 560252 465444
rect 560308 465388 560318 465444
rect 549266 462700 549276 462756
rect 549332 462700 560056 462756
rect -960 460180 480 460376
rect -960 460152 14252 460180
rect 392 460124 14252 460152
rect 14308 460124 14318 460180
rect 553522 460012 553532 460068
rect 553588 460012 560056 460068
rect 560018 457324 560028 457380
rect 560084 457324 560094 457380
rect 595560 456456 597000 456680
rect 554530 454636 554540 454692
rect 554596 454636 560056 454692
rect 554642 451948 554652 452004
rect 554708 451948 560056 452004
rect 550162 449260 550172 449316
rect 550228 449260 560056 449316
rect 553746 446572 553756 446628
rect 553812 446572 560056 446628
rect -960 446068 480 446264
rect -960 446040 19292 446068
rect 392 446012 19292 446040
rect 19348 446012 19358 446068
rect 559794 443884 559804 443940
rect 559860 443884 560056 443940
rect 595560 443240 597000 443464
rect 554418 441196 554428 441252
rect 554484 441196 560056 441252
rect 559682 438508 559692 438564
rect 559748 438508 560056 438564
rect 553522 435820 553532 435876
rect 553588 435820 560056 435876
rect 550274 433132 550284 433188
rect 550340 433132 560056 433188
rect -960 431956 480 432152
rect -960 431928 31052 431956
rect 392 431900 31052 431928
rect 31108 431900 31118 431956
rect 554642 430444 554652 430500
rect 554708 430444 560056 430500
rect 595560 430164 597000 430248
rect 590482 430108 590492 430164
rect 590548 430108 597000 430164
rect 595560 430024 597000 430108
rect 555202 427756 555212 427812
rect 555268 427756 560056 427812
rect 553858 425068 553868 425124
rect 553924 425068 560056 425124
rect 550386 422380 550396 422436
rect 550452 422380 560056 422436
rect 555314 419692 555324 419748
rect 555380 419692 560056 419748
rect -960 417844 480 418040
rect -960 417816 15932 417844
rect 392 417788 15932 417816
rect 15988 417788 15998 417844
rect 553970 417004 553980 417060
rect 554036 417004 560056 417060
rect 595560 416836 597000 417032
rect 590594 416780 590604 416836
rect 590660 416808 597000 416836
rect 590660 416780 595672 416808
rect 550610 414316 550620 414372
rect 550676 414316 560056 414372
rect 552066 411628 552076 411684
rect 552132 411628 560056 411684
rect 557106 408940 557116 408996
rect 557172 408940 560056 408996
rect 557330 406252 557340 406308
rect 557396 406252 560056 406308
rect -960 403732 480 403928
rect -960 403704 4284 403732
rect 392 403676 4284 403704
rect 4340 403676 4350 403732
rect 550722 403564 550732 403620
rect 550788 403564 560056 403620
rect 595560 403592 597000 403816
rect 556882 400876 556892 400932
rect 556948 400876 560056 400932
rect 550498 398188 550508 398244
rect 550564 398188 560056 398244
rect 559346 395500 559356 395556
rect 559412 395500 560056 395556
rect 552178 393148 552188 393204
rect 552244 393148 557452 393204
rect 557508 393148 557518 393204
rect 550162 392812 550172 392868
rect 550228 392812 560056 392868
rect 595560 390404 597000 390600
rect 590706 390348 590716 390404
rect 590772 390376 597000 390404
rect 590772 390348 595672 390376
rect 550274 390124 550284 390180
rect 550340 390124 560056 390180
rect -960 389620 480 389816
rect -960 389592 9212 389620
rect 392 389564 9212 389592
rect 9268 389564 9278 389620
rect 556994 387436 557004 387492
rect 557060 387436 560056 387492
rect 557106 384748 557116 384804
rect 557172 384748 560056 384804
rect 557666 379708 557676 379764
rect 557732 379708 559468 379764
rect 559524 379708 559534 379764
rect 588802 379708 588812 379764
rect 588868 379708 590604 379764
rect 590660 379708 590670 379764
rect 558674 378812 558684 378868
rect 558740 378812 590716 378868
rect 590772 378812 590782 378868
rect 578834 377804 578844 377860
rect 578900 377804 584668 377860
rect 584724 377804 584734 377860
rect 583538 377580 583548 377636
rect 583604 377580 586460 377636
rect 586516 377580 586526 377636
rect 550946 377468 550956 377524
rect 551012 377468 564060 377524
rect 564116 377468 564126 377524
rect 552626 377356 552636 377412
rect 552692 377356 566076 377412
rect 566132 377356 566142 377412
rect 567410 377356 567420 377412
rect 567476 377356 573244 377412
rect 573300 377356 573310 377412
rect 549042 377244 549052 377300
rect 549108 377244 565404 377300
rect 565460 377244 565470 377300
rect 568082 377244 568092 377300
rect 568148 377244 574812 377300
rect 574868 377244 574878 377300
rect 595560 377188 597000 377384
rect 557666 377132 557676 377188
rect 557732 377132 584892 377188
rect 584948 377132 584958 377188
rect 590146 377132 590156 377188
rect 590212 377160 597000 377188
rect 590212 377132 595672 377160
rect 574802 376908 574812 376964
rect 574868 376908 579964 376964
rect 580020 376908 580030 376964
rect 564722 376796 564732 376852
rect 564788 376796 571340 376852
rect 571396 376796 571406 376852
rect 575474 376796 575484 376852
rect 575540 376796 581308 376852
rect 581364 376796 581374 376852
rect 568754 376684 568764 376740
rect 568820 376684 571228 376740
rect 571284 376684 571294 376740
rect 577042 376684 577052 376740
rect 577108 376684 580860 376740
rect 580916 376684 580926 376740
rect 566738 376572 566748 376628
rect 566804 376572 569884 376628
rect 569940 376572 569950 376628
rect 570098 376572 570108 376628
rect 570164 376572 571116 376628
rect 571172 376572 571182 376628
rect 571442 376572 571452 376628
rect 571508 376572 572684 376628
rect 572740 376572 572750 376628
rect 573458 376572 573468 376628
rect 573524 376572 574364 376628
rect 574420 376572 574430 376628
rect 574578 376572 574588 376628
rect 574644 376572 576156 376628
rect 576212 376572 576222 376628
rect 577490 376572 577500 376628
rect 577556 376572 579852 376628
rect 579908 376572 579918 376628
rect 584882 376572 584892 376628
rect 584948 376572 586236 376628
rect 586292 376572 586302 376628
rect 563378 376460 563388 376516
rect 563444 376460 564396 376516
rect 564452 376460 564462 376516
rect 569426 376460 569436 376516
rect 569492 376460 569996 376516
rect 570052 376460 570062 376516
rect 570966 376460 571004 376516
rect 571060 376460 571070 376516
rect 572534 376460 572572 376516
rect 572628 376460 572638 376516
rect 572758 376460 572796 376516
rect 572852 376460 572862 376516
rect 574438 376460 574476 376516
rect 574532 376460 574542 376516
rect 576258 376460 576268 376516
rect 576324 376460 576828 376516
rect 576884 376460 576894 376516
rect 577938 376460 577948 376516
rect 578004 376460 579516 376516
rect 579572 376460 579582 376516
rect 581494 376460 581532 376516
rect 581588 376460 581598 376516
rect 582082 376460 582092 376516
rect 582148 376460 584220 376516
rect 584276 376460 584286 376516
rect 584770 376460 584780 376516
rect 584836 376460 585564 376516
rect 585620 376460 585630 376516
rect 586338 376460 586348 376516
rect 586404 376460 586908 376516
rect 586964 376460 586974 376516
rect 575362 376348 575372 376404
rect 575428 376348 578172 376404
rect 578228 376348 578238 376404
rect 573682 376236 573692 376292
rect 573748 376236 582204 376292
rect 582260 376236 582270 376292
rect -960 375508 480 375704
rect 566962 375564 566972 375620
rect 567028 375564 580188 375620
rect 580244 375564 580254 375620
rect -960 375480 17612 375508
rect 392 375452 17612 375480
rect 17668 375452 17678 375508
rect 575362 375452 575372 375508
rect 575428 375452 590156 375508
rect 590212 375452 590222 375508
rect 595560 363944 597000 364168
rect -960 361396 480 361592
rect -960 361368 37884 361396
rect 392 361340 37884 361368
rect 37940 361340 37950 361396
rect 595560 350756 597000 350952
rect 587122 350700 587132 350756
rect 587188 350728 597000 350756
rect 587188 350700 595672 350728
rect -960 347284 480 347480
rect -960 347256 29372 347284
rect 392 347228 29372 347256
rect 29428 347228 29438 347284
rect 595560 337540 597000 337736
rect 591154 337484 591164 337540
rect 591220 337512 597000 337540
rect 591220 337484 595672 337512
rect -960 333172 480 333368
rect -960 333144 19404 333172
rect 392 333116 19404 333144
rect 19460 333116 19470 333172
rect 595560 324296 597000 324520
rect -960 319060 480 319256
rect -960 319032 36204 319060
rect 392 319004 36204 319032
rect 36260 319004 36270 319060
rect 595560 311108 597000 311304
rect 576370 311052 576380 311108
rect 576436 311080 597000 311108
rect 576436 311052 595672 311080
rect -960 304948 480 305144
rect -960 304920 32732 304948
rect 392 304892 32732 304920
rect 32788 304892 32798 304948
rect 595560 297892 597000 298088
rect 588914 297836 588924 297892
rect 588980 297864 597000 297892
rect 588980 297836 595672 297864
rect -960 290836 480 291032
rect -960 290808 22764 290836
rect 392 290780 22764 290808
rect 22820 290780 22830 290836
rect 595560 284648 597000 284872
rect -960 276724 480 276920
rect -960 276696 34524 276724
rect 392 276668 34524 276696
rect 34580 276668 34590 276724
rect 595560 271460 597000 271656
rect 591266 271404 591276 271460
rect 591332 271432 597000 271460
rect 591332 271404 595672 271432
rect -960 262612 480 262808
rect -960 262584 6076 262612
rect 392 262556 6076 262584
rect 6132 262556 6142 262612
rect 595560 258216 597000 258440
rect -960 248500 480 248696
rect -960 248472 27804 248500
rect 392 248444 27804 248472
rect 27860 248444 27870 248500
rect 575586 246092 575596 246148
rect 575652 246092 590492 246148
rect 590548 246092 590558 246148
rect 595560 245028 597000 245224
rect 591154 244972 591164 245028
rect 591220 245000 597000 245028
rect 591220 244972 595672 245000
rect -960 234388 480 234584
rect -960 234360 44492 234388
rect 392 234332 44492 234360
rect 44548 234332 44558 234388
rect 221554 232652 221564 232708
rect 221620 232652 242956 232708
rect 243012 232652 243022 232708
rect 207218 232540 207228 232596
rect 207284 232540 552300 232596
rect 552356 232540 552366 232596
rect 200050 232428 200060 232484
rect 200116 232428 549388 232484
rect 549444 232428 549454 232484
rect 214386 232316 214396 232372
rect 214452 232316 247772 232372
rect 247828 232316 247838 232372
rect 71026 232204 71036 232260
rect 71092 232204 243628 232260
rect 243684 232204 243694 232260
rect 135538 232092 135548 232148
rect 135604 232092 315868 232148
rect 315924 232092 315934 232148
rect 228722 231980 228732 232036
rect 228788 231980 240156 232036
rect 240212 231980 240222 232036
rect 595560 231924 597000 232008
rect 235890 231868 235900 231924
rect 235956 231868 242732 231924
rect 242788 231868 242798 231924
rect 592946 231868 592956 231924
rect 593012 231868 597000 231924
rect 595560 231784 597000 231868
rect 106866 230748 106876 230804
rect 106932 230748 246876 230804
rect 246932 230748 246942 230804
rect 114034 230636 114044 230692
rect 114100 230636 289884 230692
rect 289940 230636 289950 230692
rect 171378 230524 171388 230580
rect 171444 230524 409836 230580
rect 409892 230524 409902 230580
rect 85362 230412 85372 230468
rect 85428 230412 391916 230468
rect 391972 230412 391982 230468
rect 185714 230300 185724 230356
rect 185780 230300 505148 230356
rect 505204 230300 505214 230356
rect 149874 230188 149884 230244
rect 149940 230188 474796 230244
rect 474852 230188 474862 230244
rect 179218 229964 179228 230020
rect 179284 229964 524076 230020
rect 524132 229964 524142 230020
rect 157042 229852 157052 229908
rect 157108 229852 456764 229908
rect 456820 229852 456830 229908
rect 121202 229740 121212 229796
rect 121268 229740 244412 229796
rect 244468 229740 244478 229796
rect 92530 229628 92540 229684
rect 92596 229628 241948 229684
rect 242004 229628 242014 229684
rect 164210 229516 164220 229572
rect 164276 229516 491372 229572
rect 491428 229516 491438 229572
rect 78642 229404 78652 229460
rect 78708 229404 80892 229460
rect 80948 229404 80958 229460
rect 128370 229404 128380 229460
rect 128436 229404 552748 229460
rect 552804 229404 552814 229460
rect 63830 229292 63868 229348
rect 63924 229292 63934 229348
rect 192882 229292 192892 229348
rect 192948 229292 193228 229348
rect 193284 229292 193294 229348
rect 80882 227836 80892 227892
rect 80948 227836 375340 227892
rect 375396 227836 375406 227892
rect 193218 227724 193228 227780
rect 193284 227724 553196 227780
rect 553252 227724 553262 227780
rect 63858 227612 63868 227668
rect 63924 227612 424956 227668
rect 425012 227612 425022 227668
rect 551842 226828 551852 226884
rect 551908 226828 553644 226884
rect 553700 226828 553710 226884
rect 40786 225148 40796 225204
rect 40852 225148 60088 225204
rect 243618 224476 243628 224532
rect 243684 224476 358764 224532
rect 358820 224476 358830 224532
rect 315858 224364 315868 224420
rect 315924 224364 552860 224420
rect 552916 224364 552926 224420
rect 240146 224252 240156 224308
rect 240212 224252 552972 224308
rect 553028 224252 553038 224308
rect 456754 223356 456764 223412
rect 456820 223356 458220 223412
rect 458276 223356 458286 223412
rect 505138 223356 505148 223412
rect 505204 223356 507948 223412
rect 508004 223356 508014 223412
rect 241938 222684 241948 222740
rect 242004 222684 408492 222740
rect 408548 222684 408558 222740
rect 409826 222684 409836 222740
rect 409892 222684 541100 222740
rect 541156 222684 541166 222740
rect 246866 222572 246876 222628
rect 246932 222572 441644 222628
rect 441700 222572 441710 222628
rect 40674 221340 40684 221396
rect 40740 221340 60088 221396
rect 239960 220668 243068 220724
rect 243124 220668 243134 220724
rect -960 220276 480 220472
rect -960 220248 4396 220276
rect 392 220220 4396 220248
rect 4452 220220 4462 220276
rect 347218 219660 347228 219716
rect 347284 219660 559468 219716
rect 559524 219660 559534 219716
rect 347554 219548 347564 219604
rect 347620 219548 557004 219604
rect 557060 219548 557070 219604
rect 247762 219436 247772 219492
rect 247828 219436 553084 219492
rect 553140 219436 553150 219492
rect 239960 218652 246092 218708
rect 246148 218652 246158 218708
rect 595560 218568 597000 218792
rect 556098 218428 556108 218484
rect 556164 218428 557004 218484
rect 557060 218428 557070 218484
rect 243058 217756 243068 217812
rect 243124 217756 274652 217812
rect 274708 217756 274718 217812
rect 242946 217644 242956 217700
rect 243012 217644 549388 217700
rect 549444 217644 549454 217700
rect 41010 217532 41020 217588
rect 41076 217532 60088 217588
rect 242722 217532 242732 217588
rect 242788 217532 552860 217588
rect 552916 217532 552926 217588
rect 347666 216972 347676 217028
rect 347732 216972 551852 217028
rect 551908 216972 551918 217028
rect 347330 216860 347340 216916
rect 347396 216860 552188 216916
rect 552244 216860 552254 216916
rect 347442 216748 347452 216804
rect 347508 216748 556220 216804
rect 556276 216748 557228 216804
rect 557284 216748 557294 216804
rect 239960 216636 266252 216692
rect 266308 216636 266318 216692
rect 408212 216636 431788 216692
rect 408212 216580 408268 216636
rect 350588 216524 408268 216580
rect 431732 216580 431788 216636
rect 478772 216636 502348 216692
rect 478772 216580 478828 216636
rect 431732 216524 478828 216580
rect 502292 216580 502348 216636
rect 502292 216524 552524 216580
rect 552580 216524 555212 216580
rect 555268 216524 555278 216580
rect 350588 215908 350644 216524
rect 343522 215852 343532 215908
rect 343588 215880 350644 215908
rect 343588 215852 350616 215880
rect 239960 214620 252812 214676
rect 252868 214620 252878 214676
rect 549378 214284 549388 214340
rect 549444 214284 549454 214340
rect 43586 213724 43596 213780
rect 43652 213724 60088 213780
rect 549388 213640 549444 214284
rect 239960 212604 242956 212660
rect 243012 212604 243022 212660
rect 239960 210588 251132 210644
rect 251188 210588 251198 210644
rect 350028 210084 350084 210504
rect 343634 210028 343644 210084
rect 343700 210028 347676 210084
rect 347732 210028 350084 210084
rect 40226 209916 40236 209972
rect 40292 209916 60088 209972
rect 239960 208572 242732 208628
rect 242788 208572 242798 208628
rect 239960 206556 243068 206612
rect 243124 206556 243134 206612
rect -960 206164 480 206360
rect -960 206136 29484 206164
rect 392 206108 29484 206136
rect 29540 206108 29550 206164
rect 41122 206108 41132 206164
rect 41188 206108 60088 206164
rect 244402 205772 244412 205828
rect 244468 205772 347340 205828
rect 347396 205772 350084 205828
rect 350028 205128 350084 205772
rect 595560 205380 597000 205576
rect 591042 205324 591052 205380
rect 591108 205352 597000 205380
rect 591108 205324 595672 205352
rect 239960 204540 242844 204596
rect 242900 204540 242910 204596
rect 10994 204092 11004 204148
rect 11060 204092 53788 204148
rect 53844 204092 53854 204148
rect 549864 203756 553084 203812
rect 553140 203756 553150 203812
rect 239960 202524 243180 202580
rect 243236 202524 243246 202580
rect 53778 202300 53788 202356
rect 53844 202300 60088 202356
rect 239960 200508 264572 200564
rect 264628 200508 264638 200564
rect 552066 199836 552076 199892
rect 552132 199836 556220 199892
rect 556276 199836 556286 199892
rect 347442 199724 347452 199780
rect 347508 199724 350056 199780
rect 33058 198492 33068 198548
rect 33124 198492 60088 198548
rect 239960 198492 271292 198548
rect 271348 198492 271358 198548
rect 239960 196476 261212 196532
rect 261268 196476 261278 196532
rect 40898 194684 40908 194740
rect 40964 194684 60088 194740
rect 239960 194460 269612 194516
rect 269668 194460 269678 194516
rect 347554 194348 347564 194404
rect 347620 194348 350056 194404
rect 549864 193900 552748 193956
rect 552804 193900 552814 193956
rect 552290 193228 552300 193284
rect 552356 193228 556108 193284
rect 556164 193228 556174 193284
rect 239960 192444 262892 192500
rect 262948 192444 262958 192500
rect -960 192052 480 192248
rect 595560 192136 597000 192360
rect -960 192024 41132 192052
rect 392 191996 41132 192024
rect 41188 191996 41198 192052
rect 37762 190876 37772 190932
rect 37828 190876 60088 190932
rect 239960 190428 257852 190484
rect 257908 190428 257918 190484
rect 551618 189756 551628 189812
rect 551684 189756 559468 189812
rect 559524 189756 559534 189812
rect 243170 188972 243180 189028
rect 243236 188972 276332 189028
rect 276388 188972 276398 189028
rect 347218 188972 347228 189028
rect 347284 188972 350056 189028
rect 239960 188412 247772 188468
rect 247828 188412 247838 188468
rect 27682 187068 27692 187124
rect 27748 187068 60088 187124
rect 239960 186396 267932 186452
rect 267988 186396 267998 186452
rect 243058 185612 243068 185668
rect 243124 185612 276444 185668
rect 276500 185612 276510 185668
rect 239960 184380 249452 184436
rect 249508 184380 249518 184436
rect 549378 184380 549388 184436
rect 549444 184380 549454 184436
rect 549388 184072 549444 184380
rect 347666 183596 347676 183652
rect 347732 183596 350056 183652
rect 36082 183260 36092 183316
rect 36148 183260 60088 183316
rect 239960 182364 264684 182420
rect 264740 182364 264750 182420
rect 239960 180348 251244 180404
rect 251300 180348 251310 180404
rect 5842 179452 5852 179508
rect 5908 179452 60088 179508
rect 595560 178920 597000 179144
rect 239960 178332 252924 178388
rect 252980 178332 252990 178388
rect 347554 178220 347564 178276
rect 347620 178220 350056 178276
rect -960 177940 480 178136
rect -960 177912 9324 177940
rect 392 177884 9324 177912
rect 9380 177884 9390 177940
rect 239960 176316 274764 176372
rect 274820 176316 274830 176372
rect 22642 175644 22652 175700
rect 22708 175644 60088 175700
rect 242946 175532 242956 175588
rect 243012 175532 276556 175588
rect 276612 175532 276622 175588
rect 239960 174300 246204 174356
rect 246260 174300 246270 174356
rect 549864 174188 552972 174244
rect 553028 174188 553038 174244
rect 347442 172844 347452 172900
rect 347508 172844 350056 172900
rect 239960 172284 241948 172340
rect 242004 172284 242014 172340
rect 244402 172172 244412 172228
rect 244468 172172 309820 172228
rect 309876 172172 309886 172228
rect 34402 171836 34412 171892
rect 34468 171836 60088 171892
rect 241938 170492 241948 170548
rect 242004 170492 266364 170548
rect 266420 170492 266430 170548
rect 239960 170268 271404 170324
rect 271460 170268 271470 170324
rect 239960 168252 261324 168308
rect 261380 168252 261390 168308
rect 12562 168028 12572 168084
rect 12628 168028 60088 168084
rect 346882 167468 346892 167524
rect 346948 167468 350056 167524
rect 239960 166236 247884 166292
rect 247940 166236 247950 166292
rect 595560 165704 597000 165928
rect 274642 165228 274652 165284
rect 274708 165228 280056 165284
rect 549864 164332 552860 164388
rect 552916 164332 552926 164388
rect 4162 164220 4172 164276
rect 4228 164220 60088 164276
rect 239960 164220 263004 164276
rect 263060 164220 263070 164276
rect 246082 164108 246092 164164
rect 246148 164108 280056 164164
rect -960 163828 480 164024
rect -960 163800 12572 163828
rect 392 163772 12572 163800
rect 12628 163772 12638 163828
rect 266242 162988 266252 163044
rect 266308 162988 280056 163044
rect 239960 162204 244524 162260
rect 244580 162204 244590 162260
rect 347330 162092 347340 162148
rect 347396 162092 350056 162148
rect 252802 161868 252812 161924
rect 252868 161868 280056 161924
rect 276546 160748 276556 160804
rect 276612 160748 280056 160804
rect 5954 160412 5964 160468
rect 6020 160412 60088 160468
rect 239960 160188 269724 160244
rect 269780 160188 269790 160244
rect 251122 159628 251132 159684
rect 251188 159628 280056 159684
rect 242722 158508 242732 158564
rect 242788 158508 280056 158564
rect 239960 158172 257964 158228
rect 258020 158172 258030 158228
rect 276434 157388 276444 157444
rect 276500 157388 280056 157444
rect 344306 156716 344316 156772
rect 344372 156716 350056 156772
rect 14242 156604 14252 156660
rect 14308 156604 60088 156660
rect 242834 156268 242844 156324
rect 242900 156268 280056 156324
rect 239960 156156 274652 156212
rect 274708 156156 274718 156212
rect 264562 155372 264572 155428
rect 264628 155372 275548 155428
rect 275604 155372 275614 155428
rect 276322 155148 276332 155204
rect 276388 155148 280056 155204
rect 549864 154476 553196 154532
rect 553252 154476 553262 154532
rect 239960 154140 241948 154196
rect 242004 154140 242014 154196
rect 275538 154028 275548 154084
rect 275604 154028 280056 154084
rect 271282 152908 271292 152964
rect 271348 152908 280056 152964
rect 19282 152796 19292 152852
rect 19348 152796 60088 152852
rect 595560 152488 597000 152712
rect 239960 152124 264572 152180
rect 264628 152124 264638 152180
rect 261202 151788 261212 151844
rect 261268 151788 280056 151844
rect 344194 151340 344204 151396
rect 344260 151340 350056 151396
rect 269602 150668 269612 150724
rect 269668 150668 280056 150724
rect 31042 150332 31052 150388
rect 31108 150332 55468 150388
rect 55524 150332 55534 150388
rect 241938 150332 241948 150388
rect 242004 150332 268044 150388
rect 268100 150332 268110 150388
rect 239960 150108 243068 150164
rect 243124 150108 243134 150164
rect -960 149716 480 149912
rect -960 149688 10892 149716
rect 392 149660 10892 149688
rect 10948 149660 10958 149716
rect 262882 149548 262892 149604
rect 262948 149548 280056 149604
rect 55458 148988 55468 149044
rect 55524 148988 60088 149044
rect 257842 148428 257852 148484
rect 257908 148428 280056 148484
rect 239960 148092 242732 148148
rect 242788 148092 242798 148148
rect 247762 147308 247772 147364
rect 247828 147308 280056 147364
rect 267922 146188 267932 146244
rect 267988 146188 280056 146244
rect 239960 146076 242844 146132
rect 242900 146076 242910 146132
rect 344082 145964 344092 146020
rect 344148 145964 350056 146020
rect 243058 145292 243068 145348
rect 243124 145292 249676 145348
rect 249732 145292 249742 145348
rect 15922 145180 15932 145236
rect 15988 145180 60088 145236
rect 249442 145068 249452 145124
rect 249508 145068 280056 145124
rect 549864 144620 552860 144676
rect 552916 144620 552926 144676
rect 239960 144060 243068 144116
rect 243124 144060 243134 144116
rect 264674 143948 264684 144004
rect 264740 143948 280056 144004
rect 251234 142828 251244 142884
rect 251300 142828 280056 142884
rect 239960 142044 242956 142100
rect 243012 142044 243022 142100
rect 252914 141708 252924 141764
rect 252980 141708 280056 141764
rect 4274 141372 4284 141428
rect 4340 141372 60088 141428
rect 274754 140588 274764 140644
rect 274820 140588 280056 140644
rect 343970 140588 343980 140644
rect 344036 140588 350056 140644
rect 581298 140364 581308 140420
rect 581364 140364 588924 140420
rect 588980 140364 588990 140420
rect 563602 140252 563612 140308
rect 563668 140252 582876 140308
rect 582932 140252 582942 140308
rect 239960 140028 243180 140084
rect 243236 140028 243246 140084
rect 246194 139468 246204 139524
rect 246260 139468 280056 139524
rect 595560 139272 597000 139496
rect 261314 138572 261324 138628
rect 261380 138572 275548 138628
rect 275604 138572 275614 138628
rect 266354 138348 266364 138404
rect 266420 138348 280056 138404
rect 239960 138012 243404 138068
rect 243460 138012 243470 138068
rect 9202 137564 9212 137620
rect 9268 137564 60088 137620
rect 271394 137228 271404 137284
rect 271460 137228 280056 137284
rect 275538 136108 275548 136164
rect 275604 136108 280056 136164
rect 239960 135996 248108 136052
rect 248164 135996 248174 136052
rect -960 135604 480 135800
rect -960 135576 4172 135604
rect 392 135548 4172 135576
rect 4228 135548 4238 135604
rect 343858 135212 343868 135268
rect 343924 135212 350056 135268
rect 247874 134988 247884 135044
rect 247940 134988 280056 135044
rect 549864 134764 552748 134820
rect 552804 134764 552814 134820
rect 239960 133980 252812 134036
rect 252868 133980 252878 134036
rect 262994 133868 263004 133924
rect 263060 133868 280056 133924
rect 17602 133756 17612 133812
rect 17668 133756 60088 133812
rect 244514 132748 244524 132804
rect 244580 132748 280056 132804
rect 239960 131964 258188 132020
rect 258244 131964 258254 132020
rect 37874 131852 37884 131908
rect 37940 131852 57036 131908
rect 57092 131852 57102 131908
rect 257954 131852 257964 131908
rect 258020 131852 275548 131908
rect 275604 131852 275614 131908
rect 269714 131628 269724 131684
rect 269780 131628 280056 131684
rect 275538 130508 275548 130564
rect 275604 130508 280056 130564
rect 57026 129948 57036 130004
rect 57092 129948 60088 130004
rect 239960 129948 244524 130004
rect 244580 129948 244590 130004
rect 343746 129836 343756 129892
rect 343812 129836 350056 129892
rect 274642 129388 274652 129444
rect 274708 129388 280056 129444
rect 268034 128268 268044 128324
rect 268100 128268 280056 128324
rect 239960 127932 268268 127988
rect 268324 127932 268334 127988
rect 264562 127148 264572 127204
rect 264628 127148 280056 127204
rect 29362 126140 29372 126196
rect 29428 126140 60088 126196
rect 249666 126028 249676 126084
rect 249732 126028 280056 126084
rect 595560 126056 597000 126280
rect 239960 125916 243292 125972
rect 243348 125916 243358 125972
rect 242722 124908 242732 124964
rect 242788 124908 280056 124964
rect 549378 124908 549388 124964
rect 549444 124908 549454 124964
rect 347218 124460 347228 124516
rect 347284 124460 350056 124516
rect 239960 123900 246092 123956
rect 246148 123900 246158 123956
rect 242834 123788 242844 123844
rect 242900 123788 280056 123844
rect 243058 122668 243068 122724
rect 243124 122668 280056 122724
rect 19394 122332 19404 122388
rect 19460 122332 60088 122388
rect 239960 121884 242732 121940
rect 242788 121884 242798 121940
rect 248098 121772 248108 121828
rect 248164 121772 275548 121828
rect 275604 121772 275614 121828
rect -960 121492 480 121688
rect 242946 121548 242956 121604
rect 243012 121548 280056 121604
rect -960 121464 14252 121492
rect 392 121436 14252 121464
rect 14308 121436 14318 121492
rect 243170 120428 243180 120484
rect 243236 120428 280056 120484
rect 36194 120092 36204 120148
rect 36260 120092 57036 120148
rect 57092 120092 57102 120148
rect 239960 119868 242956 119924
rect 243012 119868 243022 119924
rect 243394 119308 243404 119364
rect 243460 119308 280056 119364
rect 347106 119084 347116 119140
rect 347172 119084 350056 119140
rect 57026 118524 57036 118580
rect 57092 118524 60088 118580
rect 275538 118188 275548 118244
rect 275604 118188 280056 118244
rect 239960 117852 243068 117908
rect 243124 117852 243134 117908
rect 252802 117068 252812 117124
rect 252868 117068 280056 117124
rect 258178 115948 258188 116004
rect 258244 115948 280056 116004
rect 239960 115836 243516 115892
rect 243572 115836 243582 115892
rect 549864 115052 553308 115108
rect 553364 115052 553374 115108
rect 244514 114828 244524 114884
rect 244580 114828 280056 114884
rect 32722 114716 32732 114772
rect 32788 114716 60088 114772
rect 239960 113820 242172 113876
rect 242228 113820 242238 113876
rect 268258 113708 268268 113764
rect 268324 113708 280056 113764
rect 346994 113708 347004 113764
rect 347060 113708 350056 113764
rect 22754 113372 22764 113428
rect 22820 113372 57036 113428
rect 57092 113372 57102 113428
rect 246082 113372 246092 113428
rect 246148 113372 275548 113428
rect 275604 113372 275614 113428
rect 595560 112840 597000 113064
rect 243282 112588 243292 112644
rect 243348 112588 280056 112644
rect 239960 111804 242060 111860
rect 242116 111804 242126 111860
rect 275538 111468 275548 111524
rect 275604 111468 280056 111524
rect 57026 110908 57036 110964
rect 57092 110908 60088 110964
rect 242722 110348 242732 110404
rect 242788 110348 280056 110404
rect 239960 109788 242284 109844
rect 242340 109788 242350 109844
rect 242946 109228 242956 109284
rect 243012 109228 280056 109284
rect 346994 108332 347004 108388
rect 347060 108332 350056 108388
rect 243058 108108 243068 108164
rect 243124 108108 280056 108164
rect 239960 107772 241948 107828
rect 242004 107772 242014 107828
rect -960 107380 480 107576
rect -960 107352 4284 107380
rect 392 107324 4284 107352
rect 4340 107324 4350 107380
rect 34514 107100 34524 107156
rect 34580 107100 60088 107156
rect 243506 106988 243516 107044
rect 243572 106988 280056 107044
rect 242162 105868 242172 105924
rect 242228 105868 280056 105924
rect 239960 105756 243068 105812
rect 243124 105756 243134 105812
rect 549864 105196 553420 105252
rect 553476 105196 553486 105252
rect 242050 104748 242060 104804
rect 242116 104748 280056 104804
rect 239960 103740 243628 103796
rect 243684 103740 243694 103796
rect 242274 103628 242284 103684
rect 242340 103628 280056 103684
rect 6066 103292 6076 103348
rect 6132 103292 60088 103348
rect 346770 102956 346780 103012
rect 346836 102956 350056 103012
rect 241938 102508 241948 102564
rect 242004 102508 280056 102564
rect 239960 101724 273868 101780
rect 273924 101724 273934 101780
rect 27794 101612 27804 101668
rect 27860 101612 57036 101668
rect 57092 101612 57102 101668
rect 243618 101612 243628 101668
rect 243684 101612 275548 101668
rect 275604 101612 275614 101668
rect 243058 101388 243068 101444
rect 243124 101388 280056 101444
rect 275538 100268 275548 100324
rect 275604 100268 280056 100324
rect 239960 99708 241948 99764
rect 242004 99708 242014 99764
rect 595560 99624 597000 99848
rect 57026 99484 57036 99540
rect 57092 99484 60088 99540
rect 273858 99148 273868 99204
rect 273924 99148 280056 99204
rect 241938 98028 241948 98084
rect 242004 98028 280056 98084
rect 239932 97524 239988 97720
rect 346770 97580 346780 97636
rect 346836 97580 350056 97636
rect 239932 97468 243628 97524
rect 243572 96964 243628 97468
rect 243572 96908 280056 96964
rect 44482 96572 44492 96628
rect 44548 96572 57036 96628
rect 57092 96572 57102 96628
rect 243572 95788 280056 95844
rect 243572 95732 243628 95788
rect 57026 95676 57036 95732
rect 57092 95676 60088 95732
rect 239960 95676 243628 95732
rect 549864 95340 552972 95396
rect 553028 95340 553038 95396
rect 243572 94668 280056 94724
rect 243572 94052 243628 94668
rect 239932 93996 243628 94052
rect 239932 93688 239988 93996
rect 241938 93548 241948 93604
rect 242004 93548 280056 93604
rect -960 93268 480 93464
rect -960 93240 5852 93268
rect 392 93212 5852 93240
rect 5908 93212 5918 93268
rect 243170 92428 243180 92484
rect 243236 92428 280056 92484
rect 347442 92204 347452 92260
rect 347508 92204 350056 92260
rect 4386 91868 4396 91924
rect 4452 91868 60088 91924
rect 239960 91644 241948 91700
rect 242004 91644 242014 91700
rect 243058 91308 243068 91364
rect 243124 91308 280056 91364
rect 242050 90188 242060 90244
rect 242116 90188 280056 90244
rect 41122 89852 41132 89908
rect 41188 89852 57036 89908
rect 57092 89852 57102 89908
rect 239960 89628 243180 89684
rect 243236 89628 243246 89684
rect 241938 89068 241948 89124
rect 242004 89068 280056 89124
rect 29474 88060 29484 88116
rect 29540 88060 60088 88116
rect 242162 87948 242172 88004
rect 242228 87948 280056 88004
rect 239960 87612 243068 87668
rect 243124 87612 243134 87668
rect 242274 86828 242284 86884
rect 242340 86828 280056 86884
rect 347330 86828 347340 86884
rect 347396 86828 350056 86884
rect 595560 86408 597000 86632
rect 242722 85708 242732 85764
rect 242788 85708 280056 85764
rect 239960 85596 242060 85652
rect 242116 85596 242126 85652
rect 549864 85484 553084 85540
rect 553140 85484 553150 85540
rect 12562 84812 12572 84868
rect 12628 84812 56252 84868
rect 56308 84812 56318 84868
rect 244514 84588 244524 84644
rect 244580 84588 280056 84644
rect 57026 84252 57036 84308
rect 57092 84252 60088 84308
rect 239960 83580 241948 83636
rect 242004 83580 242014 83636
rect 274754 83468 274764 83524
rect 274820 83468 280056 83524
rect 243170 82348 243180 82404
rect 243236 82348 280056 82404
rect 239960 81564 242172 81620
rect 242228 81564 242238 81620
rect 347218 81452 347228 81508
rect 347284 81452 350056 81508
rect 243282 81228 243292 81284
rect 243348 81228 280056 81284
rect 9314 80444 9324 80500
rect 9380 80444 60088 80500
rect 243058 80108 243068 80164
rect 243124 80108 280056 80164
rect 239960 79548 242284 79604
rect 242340 79548 242350 79604
rect -960 79156 480 79352
rect -960 79128 4396 79156
rect 392 79100 4396 79128
rect 4452 79100 4462 79156
rect 242834 78988 242844 79044
rect 242900 78988 280056 79044
rect 242946 77868 242956 77924
rect 243012 77868 280056 77924
rect 239960 77532 242732 77588
rect 242788 77532 242798 77588
rect 275538 76748 275548 76804
rect 275604 76748 280056 76804
rect 56242 76636 56252 76692
rect 56308 76636 60088 76692
rect 347106 76076 347116 76132
rect 347172 76076 350056 76132
rect 274642 75628 274652 75684
rect 274708 75628 280056 75684
rect 549490 75628 549500 75684
rect 549556 75628 549566 75684
rect 239960 75516 244524 75572
rect 244580 75516 244590 75572
rect 242722 74508 242732 74564
rect 242788 74508 280056 74564
rect 239960 73500 274764 73556
rect 274820 73500 274830 73556
rect 595560 73192 597000 73416
rect 244514 73052 244524 73108
rect 244580 73052 275548 73108
rect 275604 73052 275614 73108
rect 10882 72828 10892 72884
rect 10948 72828 60088 72884
rect 239960 71484 243180 71540
rect 243236 71484 243246 71540
rect 346658 70700 346668 70756
rect 346724 70700 350056 70756
rect 239960 69468 243292 69524
rect 243348 69468 243358 69524
rect 4162 69020 4172 69076
rect 4228 69020 60088 69076
rect 14242 68012 14252 68068
rect 14308 68012 55468 68068
rect 55524 68012 55534 68068
rect 239960 67452 243068 67508
rect 243124 67452 243134 67508
rect 562706 66332 562716 66388
rect 562772 66332 588028 66388
rect 588084 66332 588094 66388
rect 549864 65772 553196 65828
rect 553252 65772 553262 65828
rect 289762 65548 289772 65604
rect 289828 65548 349916 65604
rect 349972 65548 349982 65604
rect 239960 65436 242844 65492
rect 242900 65436 242910 65492
rect 347554 65324 347564 65380
rect 347620 65324 350056 65380
rect -960 65044 480 65240
rect 55458 65212 55468 65268
rect 55524 65212 60088 65268
rect -960 65016 4172 65044
rect 392 64988 4172 65016
rect 4228 64988 4238 65044
rect 566514 63756 566524 63812
rect 566580 63756 575596 63812
rect 575652 63756 575662 63812
rect 239960 63420 242956 63476
rect 243012 63420 243022 63476
rect 556658 63196 556668 63252
rect 556724 63196 558684 63252
rect 558740 63196 558750 63252
rect 586226 63196 586236 63252
rect 586292 63196 587132 63252
rect 587188 63196 587198 63252
rect 561586 63084 561596 63140
rect 561652 63084 575372 63140
rect 575428 63084 575438 63140
rect 571442 62972 571452 63028
rect 571508 62972 588812 63028
rect 588868 62972 588878 63028
rect 4274 61404 4284 61460
rect 4340 61404 60088 61460
rect 239960 61404 244524 61460
rect 244580 61404 244590 61460
rect 552514 60396 552524 60452
rect 552580 60396 558572 60452
rect 558628 60396 558638 60452
rect 591042 60396 591052 60452
rect 591108 60396 593404 60452
rect 593460 60396 593470 60452
rect 551394 60284 551404 60340
rect 551460 60284 556892 60340
rect 556948 60284 556958 60340
rect 591154 60284 591164 60340
rect 591220 60284 593516 60340
rect 593572 60284 593582 60340
rect 550946 60172 550956 60228
rect 551012 60172 557116 60228
rect 557172 60172 557182 60228
rect 588018 60172 588028 60228
rect 588084 60172 591388 60228
rect 591444 60172 591454 60228
rect 347666 59948 347676 60004
rect 347732 59948 350056 60004
rect 550050 59948 550060 60004
rect 550116 59948 557340 60004
rect 557396 59948 557406 60004
rect 595560 59976 597000 60200
rect 5842 59612 5852 59668
rect 5908 59612 57036 59668
rect 57092 59612 57102 59668
rect 239960 59388 274652 59444
rect 274708 59388 274718 59444
rect 57026 57596 57036 57652
rect 57092 57596 60088 57652
rect 239960 57372 242732 57428
rect 242788 57372 242798 57428
rect 554092 56532 554148 57064
rect 554082 56476 554092 56532
rect 554148 56476 554158 56532
rect 549864 55916 552748 55972
rect 552804 55916 552814 55972
rect 550834 55692 550844 55748
rect 550900 55692 554120 55748
rect 239960 55356 343980 55412
rect 344036 55356 344046 55412
rect 350028 53956 350084 54600
rect 549378 54348 549388 54404
rect 549444 54348 554120 54404
rect 343410 53900 343420 53956
rect 343476 53900 350084 53956
rect 4386 53788 4396 53844
rect 4452 53788 60088 53844
rect 346098 53788 346108 53844
rect 346164 53788 347676 53844
rect 347732 53788 350364 53844
rect 350420 53788 350430 53844
rect 239960 53340 350588 53396
rect 350644 53340 350654 53396
rect 593282 53228 593292 53284
rect 593348 53228 593358 53284
rect 550050 53004 550060 53060
rect 550116 53004 554120 53060
rect 242834 52892 242844 52948
rect 242900 52892 346108 52948
rect 346164 52892 346174 52948
rect 347106 51996 347116 52052
rect 347172 51996 350476 52052
rect 350532 51996 350542 52052
rect 346658 51884 346668 51940
rect 346724 51884 349804 51940
rect 349860 51884 349870 51940
rect 549378 51660 549388 51716
rect 549444 51660 554120 51716
rect 239362 51548 239372 51604
rect 239428 51548 347564 51604
rect 347620 51548 349580 51604
rect 349636 51548 349646 51604
rect 239960 51324 350140 51380
rect 350196 51324 350206 51380
rect -960 50932 480 51128
rect -960 50904 5068 50932
rect 392 50876 5068 50904
rect 5124 50876 5134 50932
rect 347218 50316 347228 50372
rect 347284 50316 349692 50372
rect 349748 50316 349758 50372
rect 4162 49980 4172 50036
rect 4228 49980 60088 50036
rect 554092 49812 554148 50344
rect 549378 49756 549388 49812
rect 549444 49756 554148 49812
rect 239960 49308 242956 49364
rect 243012 49308 243022 49364
rect 242722 49196 242732 49252
rect 242788 49224 350168 49252
rect 242788 49196 350196 49224
rect 350140 48804 350196 49196
rect 554092 48804 554148 49000
rect 350130 48748 350140 48804
rect 350196 48748 350206 48804
rect 549276 48748 554148 48804
rect 549276 48692 549332 48748
rect 549266 48636 549276 48692
rect 549332 48636 549342 48692
rect 347330 48412 347340 48468
rect 347396 48412 350364 48468
rect 350420 48412 350430 48468
rect 5058 47852 5068 47908
rect 5124 47852 57036 47908
rect 57092 47852 57102 47908
rect 552402 47628 552412 47684
rect 552468 47628 554120 47684
rect 239960 47292 343532 47348
rect 343588 47292 343598 47348
rect 595560 46760 597000 46984
rect 552290 46284 552300 46340
rect 552356 46284 554120 46340
rect 57026 46172 57036 46228
rect 57092 46172 60088 46228
rect 549388 45556 549444 46088
rect 549378 45500 549388 45556
rect 549444 45500 549454 45556
rect 347442 45388 347452 45444
rect 347508 45388 349916 45444
rect 349972 45388 349982 45444
rect 239960 45276 349580 45332
rect 349636 45276 349646 45332
rect 551730 44940 551740 44996
rect 551796 44940 554120 44996
rect 350028 43652 350084 43848
rect 350018 43596 350028 43652
rect 350084 43596 350094 43652
rect 239960 43260 241948 43316
rect 242004 43260 242014 43316
rect 242946 42812 242956 42868
rect 243012 42812 346780 42868
rect 346836 42812 349468 42868
rect 349412 42420 349468 42812
rect 554092 42644 554148 43624
rect 549276 42588 554148 42644
rect 549276 42420 549332 42588
rect 4162 42364 4172 42420
rect 4228 42364 60088 42420
rect 349412 42364 549332 42420
rect 548930 42252 548940 42308
rect 548996 42252 549276 42308
rect 549332 42252 549342 42308
rect 551058 42252 551068 42308
rect 551124 42252 554120 42308
rect 496290 41468 496300 41524
rect 496356 41468 550620 41524
rect 550676 41468 550686 41524
rect 483868 41356 550396 41412
rect 550452 41356 550462 41412
rect 483868 41300 483924 41356
rect 239932 40516 239988 41272
rect 483858 41244 483868 41300
rect 483924 41244 483934 41300
rect 488226 41244 488236 41300
rect 488292 41244 553980 41300
rect 554036 41244 554046 41300
rect 480162 41132 480172 41188
rect 480228 41132 553868 41188
rect 553924 41132 553934 41188
rect 488348 41020 490588 41076
rect 488348 40964 488404 41020
rect 346994 40908 347004 40964
rect 347060 40908 488404 40964
rect 490532 40964 490588 41020
rect 490532 40908 554120 40964
rect 593506 40908 593516 40964
rect 593572 40908 593582 40964
rect 431778 40684 431788 40740
rect 431844 40684 431882 40740
rect 472098 40684 472108 40740
rect 472164 40684 554652 40740
rect 554708 40684 554718 40740
rect 443874 40572 443884 40628
rect 443940 40572 444108 40628
rect 444164 40572 550172 40628
rect 550228 40572 550238 40628
rect 239932 40460 243628 40516
rect 436230 40460 436268 40516
rect 436324 40460 436334 40516
rect 455970 40460 455980 40516
rect 456036 40460 456204 40516
rect 456260 40460 554428 40516
rect 554484 40460 554494 40516
rect 243572 40404 243628 40460
rect 243572 40348 461132 40404
rect 461188 40348 461198 40404
rect 464034 40348 464044 40404
rect 464100 40348 553532 40404
rect 553588 40348 553598 40404
rect 468066 40236 468076 40292
rect 468132 40236 550284 40292
rect 550340 40236 550350 40292
rect 552692 40236 554652 40292
rect 554708 40236 554718 40292
rect 552692 40180 552748 40236
rect 439842 40124 439852 40180
rect 439908 40124 552748 40180
rect 415650 40012 415660 40068
rect 415716 40012 551964 40068
rect 552020 40012 552030 40068
rect 431732 39900 553532 39956
rect 553588 39900 553598 39956
rect 431732 39844 431788 39900
rect 427746 39788 427756 39844
rect 427812 39788 431788 39844
rect 447906 39788 447916 39844
rect 447972 39788 553756 39844
rect 553812 39788 553822 39844
rect 419654 39676 419692 39732
rect 419748 39676 419758 39732
rect 480134 39676 480172 39732
rect 480228 39676 480238 39732
rect 483830 39676 483868 39732
rect 483924 39676 483934 39732
rect 488198 39676 488236 39732
rect 488292 39676 488302 39732
rect 496262 39676 496300 39732
rect 496356 39676 496366 39732
rect 516422 39676 516460 39732
rect 516516 39676 516526 39732
rect 532578 39676 532588 39732
rect 532644 39676 532700 39732
rect 532756 39676 532766 39732
rect 349412 39564 554120 39620
rect 349412 39508 349468 39564
rect 240258 39452 240268 39508
rect 240324 39452 347004 39508
rect 347060 39452 349468 39508
rect 451910 39452 451948 39508
rect 452004 39452 452014 39508
rect 492258 39452 492268 39508
rect 492324 39452 553980 39508
rect 554036 39452 554046 39508
rect 459974 39340 460012 39396
rect 460068 39340 460078 39396
rect 512418 39340 512428 39396
rect 512484 39340 550732 39396
rect 550788 39340 550798 39396
rect 239960 39228 437612 39284
rect 437668 39228 437678 39284
rect 476130 39228 476140 39284
rect 476196 39228 554652 39284
rect 554708 39228 554718 39284
rect 519708 38668 520100 38724
rect 519708 38612 519764 38668
rect 4274 38556 4284 38612
rect 4340 38556 60088 38612
rect 505652 38556 519764 38612
rect 520044 38612 520100 38668
rect 520044 38556 520828 38612
rect 524486 38556 524524 38612
rect 524580 38556 524972 38612
rect 525028 38556 525038 38612
rect 505652 38500 505708 38556
rect 504802 38444 504812 38500
rect 504868 38444 505708 38500
rect 520772 38500 520828 38556
rect 520772 38444 550956 38500
rect 551012 38444 551022 38500
rect 508386 38332 508396 38388
rect 508452 38332 548828 38388
rect 548884 38332 548894 38388
rect 346994 38220 347004 38276
rect 347060 38220 554120 38276
rect 500322 38108 500332 38164
rect 500388 38108 552076 38164
rect 552132 38108 552142 38164
rect 532550 37996 532588 38052
rect 532644 37996 532654 38052
rect 540082 37996 540092 38052
rect 540148 37996 550844 38052
rect 550900 37996 550910 38052
rect 536722 37884 536732 37940
rect 536788 37884 546028 37940
rect 546084 37884 546094 37940
rect 241938 37772 241948 37828
rect 242004 37772 359212 37828
rect 359268 37772 554596 37828
rect 354470 37660 354508 37716
rect 354564 37660 354574 37716
rect 478818 37660 478828 37716
rect 478884 37660 480172 37716
rect 480228 37660 480238 37716
rect 483830 37660 483868 37716
rect 483924 37660 483934 37716
rect 487218 37660 487228 37716
rect 487284 37660 488236 37716
rect 488292 37660 488302 37716
rect 554540 37604 554596 37772
rect 549332 37548 554316 37604
rect 554372 37548 554382 37604
rect 554530 37548 554540 37604
rect 554596 37548 554606 37604
rect 549332 37492 549388 37548
rect 367042 37436 367052 37492
rect 367108 37436 549388 37492
rect 243058 37324 243068 37380
rect 243124 37324 378812 37380
rect 378868 37324 378878 37380
rect 463670 37324 463708 37380
rect 463764 37324 463774 37380
rect 241378 37212 241388 37268
rect 241444 37212 383852 37268
rect 383908 37212 383918 37268
rect 241154 37100 241164 37156
rect 241220 37100 387436 37156
rect 387492 37100 387502 37156
rect -960 36932 480 37016
rect 362870 36988 362908 37044
rect 362964 36988 362974 37044
rect 383814 36988 383852 37044
rect 383908 36988 383918 37044
rect 500294 36988 500332 37044
rect 500388 36988 500398 37044
rect 504774 36988 504812 37044
rect 504868 36988 504878 37044
rect 512390 36988 512428 37044
rect 512484 36988 512494 37044
rect 528518 36988 528556 37044
rect 528612 36988 528622 37044
rect -960 36876 4172 36932
rect 4228 36876 4238 36932
rect 347218 36876 347228 36932
rect 347284 36876 554120 36932
rect -960 36792 480 36876
rect 241938 36764 241948 36820
rect 242004 36764 549500 36820
rect 549556 36764 549566 36820
rect 242946 36652 242956 36708
rect 243012 36652 549612 36708
rect 549668 36652 549678 36708
rect 343522 36540 343532 36596
rect 343588 36540 552972 36596
rect 553028 36540 553038 36596
rect 343970 36428 343980 36484
rect 344036 36428 549388 36484
rect 549444 36428 549454 36484
rect 349570 36316 349580 36372
rect 349636 36316 553084 36372
rect 553140 36316 553150 36372
rect 241490 36204 241500 36260
rect 241556 36204 343756 36260
rect 343812 36204 343822 36260
rect 554278 36204 554316 36260
rect 554372 36204 554382 36260
rect 241042 36092 241052 36148
rect 241108 36092 427756 36148
rect 427812 36092 427822 36148
rect 343746 35532 343756 35588
rect 343812 35532 554120 35588
rect 423350 35308 423388 35364
rect 423444 35308 423454 35364
rect 350130 35196 350140 35252
rect 350196 35196 553196 35252
rect 553252 35196 553262 35252
rect 349682 35084 349692 35140
rect 349748 35084 350812 35140
rect 350868 35084 552412 35140
rect 552468 35084 552478 35140
rect 350578 34972 350588 35028
rect 350644 34972 552748 35028
rect 552804 34972 552814 35028
rect 349906 34860 349916 34916
rect 349972 34860 551740 34916
rect 551796 34860 551806 34916
rect 4162 34748 4172 34804
rect 4228 34748 60088 34804
rect 437602 34748 437612 34804
rect 437668 34748 553420 34804
rect 553476 34748 553486 34804
rect 461122 34636 461132 34692
rect 461188 34636 553308 34692
rect 553364 34636 553374 34692
rect 519138 34524 519148 34580
rect 519204 34524 520716 34580
rect 520772 34524 550508 34580
rect 550564 34524 550574 34580
rect 240146 34412 240156 34468
rect 240212 34412 337708 34468
rect 528546 34412 528556 34468
rect 528612 34412 550172 34468
rect 550228 34412 550238 34468
rect 337652 34244 337708 34412
rect 337652 34188 343868 34244
rect 343924 34188 554120 34244
rect 350354 33516 350364 33572
rect 350420 33516 552300 33572
rect 552356 33516 552366 33572
rect 595560 33544 597000 33768
rect 105074 32956 105084 33012
rect 105140 32956 403564 33012
rect 403620 32956 403630 33012
rect 81778 32844 81788 32900
rect 81844 32844 241948 32900
rect 242004 32844 242014 32900
rect 343746 32844 343756 32900
rect 343812 32844 554120 32900
rect 151666 32732 151676 32788
rect 151732 32732 508396 32788
rect 508452 32732 508462 32788
rect 223570 32620 223580 32676
rect 223636 32620 343756 32676
rect 343812 32620 343822 32676
rect 191090 32508 191100 32564
rect 191156 32508 240268 32564
rect 240324 32508 240334 32564
rect 194114 32396 194124 32452
rect 194180 32396 242844 32452
rect 242900 32396 242910 32452
rect 209906 31500 209916 31556
rect 209972 31500 344092 31556
rect 344148 31500 554120 31556
rect 200050 31388 200060 31444
rect 200116 31388 223580 31444
rect 223636 31388 223646 31444
rect 198258 31276 198268 31332
rect 198324 31276 240156 31332
rect 240212 31276 240222 31332
rect 196466 31164 196476 31220
rect 196532 31164 241500 31220
rect 241556 31164 241566 31220
rect 191492 31052 239372 31108
rect 239428 31052 239438 31108
rect 191492 30884 191548 31052
rect 188402 30828 188412 30884
rect 188468 30828 191548 30884
rect 139094 30716 139132 30772
rect 139188 30716 139198 30772
rect 140886 30716 140924 30772
rect 140980 30716 140990 30772
rect 142678 30716 142716 30772
rect 142772 30716 142782 30772
rect 144452 30716 149548 30772
rect 149846 30716 149884 30772
rect 149940 30716 149950 30772
rect 185724 30716 242956 30772
rect 243012 30716 243022 30772
rect 144452 30660 144508 30716
rect 137330 30604 137340 30660
rect 137396 30604 144508 30660
rect 149492 30548 149548 30716
rect 185724 30660 185780 30716
rect 151638 30604 151676 30660
rect 151732 30604 151742 30660
rect 153430 30604 153468 30660
rect 153524 30604 153534 30660
rect 158806 30604 158844 30660
rect 158900 30604 158910 30660
rect 160598 30604 160636 30660
rect 160692 30604 160702 30660
rect 162390 30604 162428 30660
rect 162484 30604 162494 30660
rect 185714 30604 185724 30660
rect 185780 30604 185790 30660
rect 191062 30604 191100 30660
rect 191156 30604 191166 30660
rect 196438 30604 196476 30660
rect 196532 30604 196542 30660
rect 198230 30604 198268 30660
rect 198324 30604 198334 30660
rect 200022 30604 200060 30660
rect 200116 30604 200126 30660
rect 149492 30492 476140 30548
rect 476196 30492 476206 30548
rect 135538 30380 135548 30436
rect 135604 30380 472108 30436
rect 472164 30380 472174 30436
rect 105046 30268 105084 30324
rect 105140 30268 105150 30324
rect 134418 30268 134428 30324
rect 134484 30268 468076 30324
rect 468132 30268 468142 30324
rect 96114 30156 96124 30212
rect 96180 30156 241388 30212
rect 241444 30156 241454 30212
rect 344306 30156 344316 30212
rect 344372 30156 554120 30212
rect 81750 30044 81788 30100
rect 81844 30044 81854 30100
rect 88946 30044 88956 30100
rect 89012 30044 367052 30100
rect 367108 30044 367118 30100
rect 378802 30044 378812 30100
rect 378868 30044 554540 30100
rect 554596 30044 554606 30100
rect 94332 29932 243068 29988
rect 243124 29932 243134 29988
rect 94332 29876 94388 29932
rect 94322 29820 94332 29876
rect 94388 29820 94398 29876
rect 97906 29820 97916 29876
rect 97972 29820 241164 29876
rect 241220 29820 241230 29876
rect 147830 29708 147868 29764
rect 147924 29708 147934 29764
rect 157014 29708 157052 29764
rect 157108 29708 157118 29764
rect 188374 29708 188412 29764
rect 188468 29708 188478 29764
rect 203522 29708 203532 29764
rect 203588 29708 344316 29764
rect 344372 29708 344382 29764
rect 221526 29596 221564 29652
rect 221620 29596 221630 29652
rect 394790 29596 394828 29652
rect 394884 29596 394894 29652
rect 205426 29484 205436 29540
rect 205492 29484 344204 29540
rect 344260 29484 344270 29540
rect 117506 29372 117516 29428
rect 117572 29372 407596 29428
rect 407652 29372 407662 29428
rect 344194 28812 344204 28868
rect 344260 28812 554120 28868
rect 112578 28700 112588 28756
rect 112644 28700 375340 28756
rect 375396 28700 376236 28756
rect 376292 28700 376302 28756
rect 109228 28588 371308 28644
rect 371364 28588 371374 28644
rect 593282 28588 593292 28644
rect 593348 28588 593358 28644
rect 109228 28420 109284 28588
rect 110422 28476 110460 28532
rect 110516 28476 110526 28532
rect 112214 28476 112252 28532
rect 112308 28476 112318 28532
rect 131954 28476 131964 28532
rect 132020 28476 132748 28532
rect 137778 28476 137788 28532
rect 137844 28476 139132 28532
rect 139188 28476 139198 28532
rect 139570 28476 139580 28532
rect 139636 28476 140924 28532
rect 140980 28476 140990 28532
rect 141138 28476 141148 28532
rect 141204 28476 142716 28532
rect 142772 28476 142782 28532
rect 191492 28476 194124 28532
rect 194180 28476 194190 28532
rect 201842 28476 201852 28532
rect 201908 28476 202412 28532
rect 202468 28476 209916 28532
rect 209972 28476 209982 28532
rect 215814 28476 215852 28532
rect 215908 28476 215918 28532
rect 219846 28476 219884 28532
rect 219940 28476 219950 28532
rect 220098 28476 220108 28532
rect 220164 28476 221564 28532
rect 221620 28476 221630 28532
rect 346098 28476 346108 28532
rect 346164 28476 347676 28532
rect 347732 28476 551964 28532
rect 552020 28476 552524 28532
rect 552580 28476 552590 28532
rect 90738 28364 90748 28420
rect 90804 28364 91532 28420
rect 91588 28364 109284 28420
rect 132692 28420 132748 28476
rect 191492 28420 191548 28476
rect 132692 28364 140812 28420
rect 140868 28364 140878 28420
rect 173170 28364 173180 28420
rect 173236 28364 191548 28420
rect 210802 28364 210812 28420
rect 210868 28364 347452 28420
rect 347508 28364 551740 28420
rect 551796 28364 551806 28420
rect 106642 28252 106652 28308
rect 106708 28252 117516 28308
rect 117572 28252 117582 28308
rect 155222 28252 155260 28308
rect 155316 28252 155326 28308
rect 171378 28252 171388 28308
rect 171444 28252 200732 28308
rect 200788 28252 200798 28308
rect 212482 28252 212492 28308
rect 212548 28252 347564 28308
rect 347620 28252 551628 28308
rect 551684 28252 551694 28308
rect 92530 28140 92540 28196
rect 92596 28140 112588 28196
rect 112644 28140 112654 28196
rect 124786 28140 124796 28196
rect 124852 28140 163660 28196
rect 163716 28140 163726 28196
rect 167794 28140 167804 28196
rect 167860 28140 211260 28196
rect 211316 28140 211326 28196
rect 214162 28140 214172 28196
rect 214228 28140 346108 28196
rect 346164 28140 346174 28196
rect 122994 28028 123004 28084
rect 123060 28028 169372 28084
rect 169428 28028 169438 28084
rect 169586 28028 169596 28084
rect 169652 28028 205548 28084
rect 205604 28028 242732 28084
rect 242788 28028 242798 28084
rect 158806 27916 158844 27972
rect 158900 27916 158910 27972
rect 174962 27916 174972 27972
rect 175028 27916 186284 27972
rect 186340 27916 186350 27972
rect 186470 27916 186508 27972
rect 186564 27916 186574 27972
rect 191492 27916 192220 27972
rect 192276 27916 241052 27972
rect 241108 27916 241118 27972
rect 191492 27860 191548 27916
rect 115826 27804 115836 27860
rect 115892 27804 191548 27860
rect 209010 27804 209020 27860
rect 209076 27804 346108 27860
rect 346164 27804 346892 27860
rect 346948 27804 346958 27860
rect 114034 27692 114044 27748
rect 114100 27692 198156 27748
rect 198212 27692 198222 27748
rect 217522 27692 217532 27748
rect 217588 27692 552300 27748
rect 552356 27692 552366 27748
rect 117618 27580 117628 27636
rect 117684 27580 186508 27636
rect 186564 27580 186574 27636
rect 203298 27580 203308 27636
rect 203364 27580 203644 27636
rect 203700 27580 238476 27636
rect 238532 27580 238542 27636
rect 121202 27468 121212 27524
rect 121268 27468 175084 27524
rect 175140 27468 176316 27524
rect 176372 27468 176382 27524
rect 186274 27468 186284 27524
rect 186340 27468 188412 27524
rect 188468 27468 188478 27524
rect 349412 27468 554120 27524
rect 349412 27412 349468 27468
rect 80658 27356 80668 27412
rect 80724 27356 81788 27412
rect 81844 27356 81854 27412
rect 104178 27356 104188 27412
rect 104244 27356 105084 27412
rect 105140 27356 105150 27412
rect 159618 27356 159628 27412
rect 159684 27356 160636 27412
rect 160692 27356 160702 27412
rect 161410 27356 161420 27412
rect 161476 27356 162428 27412
rect 162484 27356 162494 27412
rect 207442 27356 207452 27412
rect 207508 27356 347340 27412
rect 347396 27356 349468 27412
rect 551478 27020 551516 27076
rect 551572 27020 551582 27076
rect 69682 26908 69692 26964
rect 69748 26908 72212 26964
rect 72818 26908 72828 26964
rect 72884 26908 73836 26964
rect 73892 26908 73902 26964
rect 129378 26908 129388 26964
rect 129444 26908 135548 26964
rect 135604 26908 135614 26964
rect 147830 26908 147868 26964
rect 147924 26908 147934 26964
rect 156230 26908 156268 26964
rect 156324 26908 156334 26964
rect 551282 26908 551292 26964
rect 551348 26908 552076 26964
rect 552132 26908 552636 26964
rect 552692 26908 552702 26964
rect 72156 26852 72212 26908
rect 72156 26796 309820 26852
rect 309876 26796 545132 26852
rect 545188 26796 545198 26852
rect 144508 26684 146300 26740
rect 146356 26684 496300 26740
rect 496356 26684 496366 26740
rect 144508 26628 144564 26684
rect 58930 26572 58940 26628
rect 58996 26572 92540 26628
rect 92596 26572 92606 26628
rect 144498 26572 144508 26628
rect 144564 26572 144574 26628
rect 176306 26572 176316 26628
rect 176372 26572 439852 26628
rect 439908 26572 439918 26628
rect 45602 26460 45612 26516
rect 45668 26460 96124 26516
rect 96180 26460 96190 26516
rect 130162 26460 130172 26516
rect 130228 26460 146188 26516
rect 146244 26460 146254 26516
rect 198146 26460 198156 26516
rect 198212 26460 423388 26516
rect 423444 26460 423454 26516
rect 148418 26348 148428 26404
rect 148484 26348 187516 26404
rect 187572 26348 346780 26404
rect 346836 26348 346846 26404
rect 376226 26348 376236 26404
rect 376292 26348 554540 26404
rect 554596 26348 554606 26404
rect 72258 26236 72268 26292
rect 72324 26236 153468 26292
rect 153524 26236 153534 26292
rect 193218 26236 193228 26292
rect 193284 26236 194684 26292
rect 194740 26236 347116 26292
rect 347172 26236 347182 26292
rect 91298 26124 91308 26180
rect 91364 26124 205436 26180
rect 205492 26124 205502 26180
rect 223346 26124 223356 26180
rect 223412 26124 343644 26180
rect 343700 26124 343710 26180
rect 346098 26124 346108 26180
rect 346164 26124 554120 26180
rect 13234 26012 13244 26068
rect 13300 26012 74620 26068
rect 74676 26012 74686 26068
rect 95106 26012 95116 26068
rect 95172 26012 144508 26068
rect 144564 26012 144574 26068
rect 146178 26012 146188 26068
rect 146244 26012 146524 26068
rect 146580 26012 458668 26068
rect 458724 26012 458734 26068
rect 77970 25900 77980 25956
rect 78036 25900 151676 25956
rect 151732 25900 151742 25956
rect 391458 25900 391468 25956
rect 391524 25900 554708 25956
rect 387202 25788 387212 25844
rect 387268 25788 554428 25844
rect 554484 25788 554494 25844
rect 554652 25508 554708 25900
rect 554530 25452 554540 25508
rect 554596 25452 554708 25508
rect 171378 25340 171388 25396
rect 171444 25340 180348 25396
rect 180404 25340 180414 25396
rect 159842 25228 159852 25284
rect 159908 25228 183148 25284
rect 183204 25228 183214 25284
rect 166002 25116 166012 25172
rect 166068 25116 540092 25172
rect 540148 25116 540158 25172
rect 163874 25004 163884 25060
rect 163940 25004 536732 25060
rect 536788 25004 536798 25060
rect 144498 24892 144508 24948
rect 144564 24892 145292 24948
rect 145348 24892 492268 24948
rect 492324 24892 492334 24948
rect 101490 24780 101500 24836
rect 101556 24780 394828 24836
rect 394884 24780 394894 24836
rect 551730 24780 551740 24836
rect 551796 24780 554120 24836
rect 53218 24668 53228 24724
rect 53284 24668 94332 24724
rect 94388 24668 94398 24724
rect 163650 24668 163660 24724
rect 163716 24668 447916 24724
rect 447972 24668 447982 24724
rect 66546 24556 66556 24612
rect 66612 24556 155260 24612
rect 155316 24556 155326 24612
rect 183138 24556 183148 24612
rect 183204 24556 349916 24612
rect 349972 24556 349982 24612
rect 27682 24444 27692 24500
rect 27748 24444 166012 24500
rect 166068 24444 166078 24500
rect 192322 24444 192332 24500
rect 192388 24444 192892 24500
rect 192948 24444 347004 24500
rect 347060 24444 347070 24500
rect 27906 24332 27916 24388
rect 27972 24332 223356 24388
rect 223412 24332 223422 24388
rect 225922 24332 225932 24388
rect 225988 24332 343532 24388
rect 343588 24332 343598 24388
rect 89842 24220 89852 24276
rect 89908 24220 209020 24276
rect 209076 24220 209086 24276
rect 99698 23436 99708 23492
rect 99764 23436 391468 23492
rect 391524 23436 391534 23492
rect 551618 23436 551628 23492
rect 551684 23436 554120 23492
rect 176978 23324 176988 23380
rect 177044 23324 178556 23380
rect 178612 23324 178622 23380
rect 350130 23324 350140 23380
rect 350196 23324 550844 23380
rect 550900 23324 550910 23380
rect 189298 23212 189308 23268
rect 189364 23212 347004 23268
rect 347060 23212 347070 23268
rect 350354 23212 350364 23268
rect 350420 23212 550060 23268
rect 550116 23212 550126 23268
rect 349794 23100 349804 23156
rect 349860 23100 548604 23156
rect 548660 23100 548670 23156
rect 180338 22988 180348 23044
rect 180404 22988 350812 23044
rect 350868 22988 350878 23044
rect 392 22904 4284 22932
rect -960 22876 4284 22904
rect 4340 22876 4350 22932
rect -960 22680 480 22876
rect 119410 22652 119420 22708
rect 119476 22652 180796 22708
rect 180852 22652 435148 22708
rect 435204 22652 435214 22708
rect 551954 22092 551964 22148
rect 552020 22092 554120 22148
rect 169362 21756 169372 21812
rect 169428 21756 443884 21812
rect 443940 21756 443950 21812
rect 78194 21644 78204 21700
rect 78260 21644 289772 21700
rect 289828 21644 289838 21700
rect 350466 21644 350476 21700
rect 350532 21644 548940 21700
rect 548996 21644 549006 21700
rect 125570 21532 125580 21588
rect 125636 21532 193228 21588
rect 193284 21532 193294 21588
rect 209318 21532 209356 21588
rect 209412 21532 415660 21588
rect 415716 21532 415726 21588
rect 349570 21420 349580 21476
rect 349636 21420 548716 21476
rect 548772 21420 548782 21476
rect 55122 21308 55132 21364
rect 55188 21308 158844 21364
rect 158900 21308 158910 21364
rect 349682 21308 349692 21364
rect 349748 21308 548492 21364
rect 548548 21308 548558 21364
rect 41794 21196 41804 21252
rect 41860 21196 218428 21252
rect 218484 21196 218494 21252
rect 126578 21084 126588 21140
rect 126644 21084 157948 21140
rect 158004 21084 451948 21140
rect 452004 21084 452014 21140
rect 128370 20972 128380 21028
rect 128436 20972 152236 21028
rect 152292 20972 455980 21028
rect 456036 20972 456046 21028
rect 182242 20860 182252 20916
rect 182308 20860 350364 20916
rect 350420 20860 350430 20916
rect 551506 20748 551516 20804
rect 551572 20748 554120 20804
rect 595560 20328 597000 20552
rect 108322 20076 108332 20132
rect 108388 20076 411628 20132
rect 411684 20076 411694 20132
rect 117954 19740 117964 19796
rect 118020 19740 137788 19796
rect 137844 19740 137854 19796
rect 37986 19628 37996 19684
rect 38052 19628 97916 19684
rect 97972 19628 97982 19684
rect 131282 19628 131292 19684
rect 131348 19628 192332 19684
rect 192388 19628 192398 19684
rect 83682 19516 83692 19572
rect 83748 19516 149884 19572
rect 149940 19516 149950 19572
rect 18946 19404 18956 19460
rect 19012 19404 79212 19460
rect 79268 19404 79278 19460
rect 81442 19404 81452 19460
rect 81508 19404 210812 19460
rect 210868 19404 210878 19460
rect 552290 19404 552300 19460
rect 552356 19404 554120 19460
rect 32274 19292 32284 19348
rect 32340 19292 163884 19348
rect 163940 19292 163950 19348
rect 103282 18396 103292 18452
rect 103348 18396 399532 18452
rect 399588 18396 399598 18452
rect 349412 18284 553980 18340
rect 554036 18284 554046 18340
rect 200722 18172 200732 18228
rect 200788 18172 343420 18228
rect 343476 18172 343486 18228
rect 349412 18116 349468 18284
rect 211250 18060 211260 18116
rect 211316 18060 346892 18116
rect 346948 18060 349468 18116
rect 552626 18060 552636 18116
rect 552692 18060 554120 18116
rect 100818 17948 100828 18004
rect 100884 17948 145292 18004
rect 145348 17948 145358 18004
rect 154130 17948 154140 18004
rect 154196 17948 185724 18004
rect 185780 17948 185790 18004
rect 22754 17836 22764 17892
rect 22820 17836 101500 17892
rect 101556 17836 101566 17892
rect 119858 17836 119868 17892
rect 119924 17836 196476 17892
rect 196532 17836 196542 17892
rect 68450 17724 68460 17780
rect 68516 17724 212492 17780
rect 212548 17724 212558 17780
rect 47506 17612 47516 17668
rect 47572 17612 159628 17668
rect 159684 17612 159694 17668
rect 176754 17612 176764 17668
rect 176820 17612 182700 17668
rect 182756 17612 349804 17668
rect 349860 17612 349870 17668
rect 176978 17500 176988 17556
rect 177044 17500 350476 17556
rect 350532 17500 350542 17556
rect 199938 16828 199948 16884
rect 200004 16828 200732 16884
rect 200788 16828 200798 16884
rect 552178 16716 552188 16772
rect 552244 16716 554120 16772
rect 106530 16268 106540 16324
rect 106596 16268 141148 16324
rect 141204 16268 141214 16324
rect 593394 16268 593404 16324
rect 593460 16268 593470 16324
rect 30370 16156 30380 16212
rect 30436 16156 99708 16212
rect 99764 16156 99774 16212
rect 102722 16156 102732 16212
rect 102788 16156 202412 16212
rect 202468 16156 202478 16212
rect 41122 16044 41132 16100
rect 41188 16044 161420 16100
rect 161476 16044 161486 16100
rect 62738 15932 62748 15988
rect 62804 15932 214172 15988
rect 214228 15932 214238 15988
rect 551842 15372 551852 15428
rect 551908 15372 554120 15428
rect 142818 14588 142828 14644
rect 142884 14588 189308 14644
rect 189364 14588 189374 14644
rect 62962 14476 62972 14532
rect 63028 14476 156268 14532
rect 156324 14476 156334 14532
rect 49410 14364 49420 14420
rect 49476 14364 217532 14420
rect 217588 14364 217598 14420
rect 15138 14252 15148 14308
rect 15204 14252 225932 14308
rect 225988 14252 225998 14308
rect 228722 14252 228732 14308
rect 228788 14252 553532 14308
rect 553588 14252 553598 14308
rect 86482 13356 86492 13412
rect 86548 13356 87164 13412
rect 87220 13356 362908 13412
rect 362964 13356 362974 13412
rect 123666 13020 123676 13076
rect 123732 13020 137340 13076
rect 137396 13020 137406 13076
rect 64642 12908 64652 12964
rect 64708 12908 91532 12964
rect 91588 12908 91598 12964
rect 136994 12908 137004 12964
rect 137060 12908 190316 12964
rect 190372 12908 190382 12964
rect 89394 12796 89404 12852
rect 89460 12796 147868 12852
rect 147924 12796 147934 12852
rect 59602 12684 59612 12740
rect 59668 12684 215852 12740
rect 215908 12684 215918 12740
rect 552514 12684 552524 12740
rect 552580 12684 554120 12740
rect 11330 12572 11340 12628
rect 11396 12572 69692 12628
rect 69748 12572 69758 12628
rect 97010 12572 97020 12628
rect 97076 12572 203532 12628
rect 203588 12572 203598 12628
rect 230514 12572 230524 12628
rect 230580 12572 551852 12628
rect 551908 12572 551918 12628
rect 34402 10892 34412 10948
rect 34468 10892 220108 10948
rect 220164 10892 220174 10948
rect 554306 10780 554316 10836
rect 554372 10780 567252 10836
rect 567196 10612 567252 10780
rect 557302 10556 557340 10612
rect 557396 10556 557406 10612
rect 557554 10556 557564 10612
rect 557620 10556 560252 10612
rect 560308 10556 560318 10612
rect 567186 10556 567196 10612
rect 567252 10556 567262 10612
rect 574466 10556 574476 10612
rect 574532 10556 574588 10612
rect 574644 10556 574654 10612
rect 585974 10556 586012 10612
rect 586068 10556 586078 10612
rect 591350 10556 591388 10612
rect 591444 10556 591454 10612
rect 557442 10444 557452 10500
rect 557508 10444 559132 10500
rect 559188 10444 559198 10500
rect 559346 10444 559356 10500
rect 559412 10444 565404 10500
rect 565460 10444 565470 10500
rect 574354 10444 574364 10500
rect 574420 10444 575596 10500
rect 575652 10444 575662 10500
rect 557106 10332 557116 10388
rect 557172 10332 558012 10388
rect 558068 10332 558078 10388
rect 559990 10332 560028 10388
rect 560084 10332 560094 10388
rect 574354 10332 574364 10388
rect 574420 10332 579964 10388
rect 580020 10332 580030 10388
rect 557666 10220 557676 10276
rect 557732 10220 563612 10276
rect 563668 10220 563678 10276
rect 554642 10108 554652 10164
rect 554708 10108 557788 10164
rect 557844 10108 557854 10164
rect 558002 10108 558012 10164
rect 558068 10108 562716 10164
rect 562772 10108 562782 10164
rect 79202 9996 79212 10052
rect 79268 9996 354508 10052
rect 354564 9996 354574 10052
rect 545122 9996 545132 10052
rect 545188 9996 588924 10052
rect 588980 9996 588990 10052
rect 556994 9884 557004 9940
rect 557060 9884 561484 9940
rect 561540 9884 561550 9940
rect 567074 9884 567084 9940
rect 567140 9884 570108 9940
rect 570164 9884 570174 9940
rect 570658 9884 570668 9940
rect 570724 9884 575372 9940
rect 575428 9884 575438 9940
rect 556434 9772 556444 9828
rect 556500 9772 586348 9828
rect 586404 9772 586414 9828
rect 556882 9660 556892 9716
rect 556948 9660 564508 9716
rect 564564 9660 564574 9716
rect 568978 9660 568988 9716
rect 569044 9660 584668 9716
rect 584724 9660 584734 9716
rect 572562 9548 572572 9604
rect 572628 9548 574588 9604
rect 574644 9548 574654 9604
rect 581298 9548 581308 9604
rect 581364 9548 581374 9604
rect 581308 9492 581364 9548
rect 114370 9436 114380 9492
rect 114436 9436 198268 9492
rect 198324 9436 198334 9492
rect 573458 9436 573468 9492
rect 573524 9436 581364 9492
rect 36306 9324 36316 9380
rect 36372 9324 106652 9380
rect 106708 9324 106718 9380
rect 108658 9324 108668 9380
rect 108724 9324 200060 9380
rect 200116 9324 200126 9380
rect 571666 9324 571676 9380
rect 571732 9324 576268 9380
rect 576324 9324 576334 9380
rect 85810 9212 85820 9268
rect 85876 9212 207452 9268
rect 207508 9212 207518 9268
rect 226930 9212 226940 9268
rect 226996 9212 562940 9268
rect 562996 9212 563006 9268
rect 570770 9212 570780 9268
rect 570836 9212 579852 9268
rect 579908 9212 579918 9268
rect 549042 9100 549052 9156
rect 549108 9100 586908 9156
rect 586964 9100 586974 9156
rect 392 8792 4172 8820
rect -960 8764 4172 8792
rect 4228 8764 4238 8820
rect -960 8568 480 8764
rect 568082 8316 568092 8372
rect 568148 8316 572908 8372
rect 572964 8316 572974 8372
rect 575026 8316 575036 8372
rect 575092 8316 583324 8372
rect 583380 8316 583390 8372
rect 575036 8260 575092 8316
rect 85362 8204 85372 8260
rect 85428 8204 568988 8260
rect 569044 8204 569054 8260
rect 569202 8204 569212 8260
rect 569268 8204 575092 8260
rect 577014 8204 577052 8260
rect 577108 8204 577118 8260
rect 577612 8204 582428 8260
rect 582484 8204 582494 8260
rect 577612 8148 577668 8204
rect 571218 8092 571228 8148
rect 571284 8092 577668 8148
rect 577910 8092 577948 8148
rect 578004 8092 578014 8148
rect 578806 8092 578844 8148
rect 578900 8092 578910 8148
rect 579814 8092 579852 8148
rect 579908 8092 579918 8148
rect 196242 7980 196252 8036
rect 196308 7980 549052 8036
rect 549108 7980 549118 8036
rect 569986 7980 569996 8036
rect 570052 7980 581532 8036
rect 581588 7980 581598 8036
rect 190530 7868 190540 7924
rect 190596 7868 551068 7924
rect 551124 7868 551134 7924
rect 571106 7868 571116 7924
rect 571172 7868 580636 7924
rect 580692 7868 580702 7924
rect 51538 7756 51548 7812
rect 51604 7756 103292 7812
rect 103348 7756 103358 7812
rect 174626 7756 174636 7812
rect 174692 7756 556444 7812
rect 556500 7756 556510 7812
rect 564386 7756 564396 7812
rect 564452 7756 588700 7812
rect 588756 7756 588766 7812
rect 28690 7644 28700 7700
rect 28756 7644 108332 7700
rect 108388 7644 108398 7700
rect 165778 7644 165788 7700
rect 165844 7644 182252 7700
rect 182308 7644 182318 7700
rect 184818 7644 184828 7700
rect 184884 7644 569884 7700
rect 569940 7644 570164 7700
rect 571330 7644 571340 7700
rect 571396 7644 578620 7700
rect 578676 7644 578686 7700
rect 584612 7644 585116 7700
rect 585172 7644 585182 7700
rect 21970 7532 21980 7588
rect 22036 7532 80668 7588
rect 80724 7532 80734 7588
rect 83570 7532 83580 7588
rect 83636 7532 87500 7588
rect 87556 7532 569884 7588
rect 569940 7532 569950 7588
rect 570108 7476 570164 7644
rect 584612 7476 584668 7644
rect 570108 7420 584668 7476
rect 566962 7308 566972 7364
rect 567028 7308 572908 7364
rect 578946 7308 578956 7364
rect 579012 7308 590492 7364
rect 590548 7308 590558 7364
rect 559458 7196 559468 7252
rect 559524 7196 571340 7252
rect 571396 7196 571406 7252
rect 572852 7140 572908 7308
rect 578610 7196 578620 7252
rect 578676 7196 587804 7252
rect 587860 7196 587870 7252
rect 572852 7084 573244 7140
rect 573300 7084 584220 7140
rect 584276 7084 584286 7140
rect 595560 7112 597000 7336
rect 567970 6972 567980 7028
rect 568036 6972 569996 7028
rect 570052 6972 570062 7028
rect 574466 6860 574476 6916
rect 574532 6860 574588 6916
rect 574644 6860 574654 6916
rect 82002 6748 82012 6804
rect 82068 6748 85372 6804
rect 85428 6748 85438 6804
rect 569436 6748 571228 6804
rect 571284 6748 571294 6804
rect 577154 6748 577164 6804
rect 577220 6748 578732 6804
rect 578788 6748 578798 6804
rect 17266 6524 17276 6580
rect 17332 6524 174636 6580
rect 174692 6524 174702 6580
rect 173394 6412 173404 6468
rect 173460 6412 569212 6468
rect 569268 6412 569278 6468
rect 569436 6356 569492 6748
rect 167682 6300 167692 6356
rect 167748 6300 569492 6356
rect 112466 6188 112476 6244
rect 112532 6188 139580 6244
rect 139636 6188 139646 6244
rect 156146 6188 156156 6244
rect 156212 6188 571116 6244
rect 571172 6188 571182 6244
rect 76290 6076 76300 6132
rect 76356 6076 86492 6132
rect 86548 6076 86558 6132
rect 133410 6076 133420 6132
rect 133476 6076 572796 6132
rect 572852 6076 572862 6132
rect 70466 5964 70476 6020
rect 70532 5964 88956 6020
rect 89012 5964 89022 6020
rect 127586 5964 127596 6020
rect 127652 5964 574364 6020
rect 574420 5964 574430 6020
rect 43922 5852 43932 5908
rect 43988 5852 104188 5908
rect 104244 5852 104254 5908
rect 121986 5852 121996 5908
rect 122052 5852 574476 5908
rect 574532 5852 574542 5908
rect 74386 4956 74396 5012
rect 74452 4956 81452 5012
rect 81508 4956 81518 5012
rect 525812 4956 550956 5012
rect 551012 4956 564396 5012
rect 564452 4956 564462 5012
rect 525812 4340 525868 4956
rect 553522 4396 553532 4452
rect 553588 4396 582540 4452
rect 582596 4396 582606 4452
rect 24882 4284 24892 4340
rect 24948 4284 27692 4340
rect 27748 4284 27758 4340
rect 207666 4284 207676 4340
rect 207732 4284 525868 4340
rect 551842 4284 551852 4340
rect 551908 4284 584444 4340
rect 584500 4284 584510 4340
rect 26786 4172 26796 4228
rect 26852 4172 27916 4228
rect 27972 4172 27982 4228
rect 40114 4172 40124 4228
rect 40180 4172 41132 4228
rect 41188 4172 41198 4228
rect 57250 4172 57260 4228
rect 57316 4172 59612 4228
rect 59668 4172 59678 4228
rect 61058 4172 61068 4228
rect 61124 4172 62972 4228
rect 63028 4172 63038 4228
rect 80098 4172 80108 4228
rect 80164 4172 89852 4228
rect 89908 4172 89918 4228
rect 201954 4172 201964 4228
rect 202020 4172 559468 4228
rect 559524 4172 559534 4228
rect 562930 4172 562940 4228
rect 562996 4172 580636 4228
rect 580692 4172 580702 4228
rect 179106 3052 179116 3108
rect 179172 3052 566972 3108
rect 567028 3052 567038 3108
rect 116274 2940 116284 2996
rect 116340 2940 574364 2996
rect 574420 2940 574430 2996
rect 110562 2828 110572 2884
rect 110628 2828 573468 2884
rect 573524 2828 573534 2884
rect 104850 2716 104860 2772
rect 104916 2716 572572 2772
rect 572628 2716 572638 2772
rect 99026 2604 99036 2660
rect 99092 2604 571676 2660
rect 571732 2604 571742 2660
rect 93426 2492 93436 2548
rect 93492 2492 570780 2548
rect 570836 2492 570846 2548
rect 162642 364 162652 420
rect 162708 364 567980 420
rect 568036 364 568046 420
rect 150658 252 150668 308
rect 150724 252 571004 308
rect 571060 252 571070 308
rect 144946 140 144956 196
rect 145012 140 572684 196
rect 572740 140 572750 196
rect 139234 28 139244 84
rect 139300 28 572572 84
rect 572628 28 572638 84
<< via3 >>
rect 77308 589708 77364 589764
rect 408380 589708 408436 589764
rect 474572 589708 474628 589764
rect 540764 589708 540820 589764
rect 474572 589260 474628 589316
rect 540764 589260 540820 589316
rect 77308 588812 77364 588868
rect 408380 588812 408436 588868
rect 37772 587132 37828 587188
rect 27692 573020 27748 573076
rect 36092 558908 36148 558964
rect 5852 544796 5908 544852
rect 22652 530684 22708 530740
rect 34412 516572 34468 516628
rect 12572 502460 12628 502516
rect 4172 488348 4228 488404
rect 5964 474236 6020 474292
rect 560252 465388 560308 465444
rect 549276 462700 549332 462756
rect 14252 460124 14308 460180
rect 553532 460012 553588 460068
rect 560028 457324 560084 457380
rect 554540 454636 554596 454692
rect 554652 451948 554708 452004
rect 19292 446012 19348 446068
rect 559804 443884 559860 443940
rect 554428 441196 554484 441252
rect 559692 438508 559748 438564
rect 31052 431900 31108 431956
rect 555212 427756 555268 427812
rect 555324 419692 555380 419748
rect 15932 417788 15988 417844
rect 4284 403676 4340 403732
rect 556892 400876 556948 400932
rect 559356 395500 559412 395556
rect 550172 392812 550228 392868
rect 550284 390124 550340 390180
rect 9212 389564 9268 389620
rect 557004 387436 557060 387492
rect 557116 384748 557172 384804
rect 584668 377804 584724 377860
rect 586460 377580 586516 377636
rect 550956 377468 551012 377524
rect 552636 377356 552692 377412
rect 573244 377356 573300 377412
rect 549052 377244 549108 377300
rect 574812 377244 574868 377300
rect 557676 377132 557732 377188
rect 579964 376908 580020 376964
rect 571340 376796 571396 376852
rect 581308 376796 581364 376852
rect 571228 376684 571284 376740
rect 577052 376684 577108 376740
rect 569884 376572 569940 376628
rect 571116 376572 571172 376628
rect 572684 376572 572740 376628
rect 574364 376572 574420 376628
rect 574588 376572 574644 376628
rect 579852 376572 579908 376628
rect 584892 376572 584948 376628
rect 564396 376460 564452 376516
rect 569996 376460 570052 376516
rect 571004 376460 571060 376516
rect 572572 376460 572628 376516
rect 572796 376460 572852 376516
rect 574476 376460 574532 376516
rect 576268 376460 576324 376516
rect 577948 376460 578004 376516
rect 581532 376460 581588 376516
rect 582092 376460 582148 376516
rect 584780 376460 584836 376516
rect 586348 376460 586404 376516
rect 575372 376348 575428 376404
rect 573692 376236 573748 376292
rect 566972 375564 567028 375620
rect 17612 375452 17668 375508
rect 37884 361340 37940 361396
rect 29372 347228 29428 347284
rect 19404 333116 19460 333172
rect 36204 319004 36260 319060
rect 32732 304892 32788 304948
rect 22764 290780 22820 290836
rect 34524 276668 34580 276724
rect 591276 271404 591332 271460
rect 6076 262556 6132 262612
rect 27804 248444 27860 248500
rect 591164 244972 591220 245028
rect 44492 234332 44548 234388
rect 592956 231868 593012 231924
rect 80892 229404 80948 229460
rect 552748 229404 552804 229460
rect 63868 229292 63924 229348
rect 193228 229292 193284 229348
rect 80892 227836 80948 227892
rect 193228 227724 193284 227780
rect 63868 227612 63924 227668
rect 551852 226828 551908 226884
rect 552860 224364 552916 224420
rect 243068 220668 243124 220724
rect 4396 220220 4452 220276
rect 246092 218652 246148 218708
rect 243068 217756 243124 217812
rect 274652 217756 274708 217812
rect 549388 217644 549444 217700
rect 551852 216972 551908 217028
rect 266252 216636 266308 216692
rect 552524 216524 552580 216580
rect 252812 214620 252868 214676
rect 549388 214284 549444 214340
rect 242956 212604 243012 212660
rect 251132 210588 251188 210644
rect 242732 208572 242788 208628
rect 243068 206556 243124 206612
rect 29484 206108 29540 206164
rect 244412 205772 244468 205828
rect 591052 205324 591108 205380
rect 242844 204540 242900 204596
rect 243180 202524 243236 202580
rect 264572 200508 264628 200564
rect 552076 199836 552132 199892
rect 271292 198492 271348 198548
rect 261212 196476 261268 196532
rect 269612 194460 269668 194516
rect 552300 193228 552356 193284
rect 262892 192444 262948 192500
rect 41132 191996 41188 192052
rect 37772 190876 37828 190932
rect 257852 190428 257908 190484
rect 551628 189756 551684 189812
rect 243180 188972 243236 189028
rect 276332 188972 276388 189028
rect 247772 188412 247828 188468
rect 27692 187068 27748 187124
rect 267932 186396 267988 186452
rect 243068 185612 243124 185668
rect 276444 185612 276500 185668
rect 249452 184380 249508 184436
rect 347676 183596 347732 183652
rect 36092 183260 36148 183316
rect 264684 182364 264740 182420
rect 251244 180348 251300 180404
rect 5852 179452 5908 179508
rect 252924 178332 252980 178388
rect 347564 178220 347620 178276
rect 9324 177884 9380 177940
rect 274764 176316 274820 176372
rect 22652 175644 22708 175700
rect 242956 175532 243012 175588
rect 276556 175532 276612 175588
rect 246204 174300 246260 174356
rect 347452 172844 347508 172900
rect 241948 172284 242004 172340
rect 34412 171836 34468 171892
rect 241948 170492 242004 170548
rect 266364 170492 266420 170548
rect 271404 170268 271460 170324
rect 261324 168252 261380 168308
rect 12572 168028 12628 168084
rect 346892 167468 346948 167524
rect 247884 166236 247940 166292
rect 274652 165228 274708 165284
rect 4172 164220 4228 164276
rect 263004 164220 263060 164276
rect 246092 164108 246148 164164
rect 12572 163772 12628 163828
rect 266252 162988 266308 163044
rect 244524 162204 244580 162260
rect 347340 162092 347396 162148
rect 252812 161868 252868 161924
rect 276556 160748 276612 160804
rect 5964 160412 6020 160468
rect 269724 160188 269780 160244
rect 251132 159628 251188 159684
rect 242732 158508 242788 158564
rect 257964 158172 258020 158228
rect 276444 157388 276500 157444
rect 14252 156604 14308 156660
rect 242844 156268 242900 156324
rect 274652 156156 274708 156212
rect 264572 155372 264628 155428
rect 275548 155372 275604 155428
rect 276332 155148 276388 155204
rect 241948 154140 242004 154196
rect 275548 154028 275604 154084
rect 271292 152908 271348 152964
rect 19292 152796 19348 152852
rect 264572 152124 264628 152180
rect 261212 151788 261268 151844
rect 269612 150668 269668 150724
rect 31052 150332 31108 150388
rect 55468 150332 55524 150388
rect 241948 150332 242004 150388
rect 268044 150332 268100 150388
rect 243068 150108 243124 150164
rect 10892 149660 10948 149716
rect 262892 149548 262948 149604
rect 55468 148988 55524 149044
rect 257852 148428 257908 148484
rect 242732 148092 242788 148148
rect 247772 147308 247828 147364
rect 267932 146188 267988 146244
rect 242844 146076 242900 146132
rect 243068 145292 243124 145348
rect 249676 145292 249732 145348
rect 15932 145180 15988 145236
rect 249452 145068 249508 145124
rect 552860 144620 552916 144676
rect 243068 144060 243124 144116
rect 264684 143948 264740 144004
rect 251244 142828 251300 142884
rect 242956 142044 243012 142100
rect 252924 141708 252980 141764
rect 4284 141372 4340 141428
rect 274764 140588 274820 140644
rect 563612 140252 563668 140308
rect 243180 140028 243236 140084
rect 246204 139468 246260 139524
rect 261324 138572 261380 138628
rect 275548 138572 275604 138628
rect 266364 138348 266420 138404
rect 243404 138012 243460 138068
rect 9212 137564 9268 137620
rect 271404 137228 271460 137284
rect 275548 136108 275604 136164
rect 248108 135996 248164 136052
rect 4172 135548 4228 135604
rect 247884 134988 247940 135044
rect 552748 134764 552804 134820
rect 252812 133980 252868 134036
rect 263004 133868 263060 133924
rect 17612 133756 17668 133812
rect 244524 132748 244580 132804
rect 258188 131964 258244 132020
rect 37884 131852 37940 131908
rect 57036 131852 57092 131908
rect 257964 131852 258020 131908
rect 275548 131852 275604 131908
rect 269724 131628 269780 131684
rect 275548 130508 275604 130564
rect 57036 129948 57092 130004
rect 244524 129948 244580 130004
rect 274652 129388 274708 129444
rect 268044 128268 268100 128324
rect 268268 127932 268324 127988
rect 264572 127148 264628 127204
rect 29372 126140 29428 126196
rect 249676 126028 249732 126084
rect 243292 125916 243348 125972
rect 242732 124908 242788 124964
rect 549388 124908 549444 124964
rect 347228 124460 347284 124516
rect 246092 123900 246148 123956
rect 242844 123788 242900 123844
rect 243068 122668 243124 122724
rect 19404 122332 19460 122388
rect 242732 121884 242788 121940
rect 248108 121772 248164 121828
rect 275548 121772 275604 121828
rect 242956 121548 243012 121604
rect 14252 121436 14308 121492
rect 243180 120428 243236 120484
rect 36204 120092 36260 120148
rect 57036 120092 57092 120148
rect 242956 119868 243012 119924
rect 243404 119308 243460 119364
rect 347116 119084 347172 119140
rect 57036 118524 57092 118580
rect 275548 118188 275604 118244
rect 243068 117852 243124 117908
rect 252812 117068 252868 117124
rect 258188 115948 258244 116004
rect 243516 115836 243572 115892
rect 553308 115052 553364 115108
rect 244524 114828 244580 114884
rect 32732 114716 32788 114772
rect 242172 113820 242228 113876
rect 268268 113708 268324 113764
rect 347004 113708 347060 113764
rect 22764 113372 22820 113428
rect 57036 113372 57092 113428
rect 246092 113372 246148 113428
rect 275548 113372 275604 113428
rect 243292 112588 243348 112644
rect 242060 111804 242116 111860
rect 275548 111468 275604 111524
rect 57036 110908 57092 110964
rect 242732 110348 242788 110404
rect 242284 109788 242340 109844
rect 242956 109228 243012 109284
rect 243068 108108 243124 108164
rect 241948 107772 242004 107828
rect 4284 107324 4340 107380
rect 34524 107100 34580 107156
rect 243516 106988 243572 107044
rect 242172 105868 242228 105924
rect 243068 105756 243124 105812
rect 553420 105196 553476 105252
rect 242060 104748 242116 104804
rect 243628 103740 243684 103796
rect 242284 103628 242340 103684
rect 6076 103292 6132 103348
rect 346780 102956 346836 103012
rect 241948 102508 242004 102564
rect 273868 101724 273924 101780
rect 27804 101612 27860 101668
rect 57036 101612 57092 101668
rect 243628 101612 243684 101668
rect 275548 101612 275604 101668
rect 243068 101388 243124 101444
rect 275548 100268 275604 100324
rect 241948 99708 242004 99764
rect 57036 99484 57092 99540
rect 273868 99148 273924 99204
rect 241948 98028 242004 98084
rect 44492 96572 44548 96628
rect 57036 96572 57092 96628
rect 57036 95676 57092 95732
rect 552972 95340 553028 95396
rect 241948 93548 242004 93604
rect 5852 93212 5908 93268
rect 243180 92428 243236 92484
rect 4396 91868 4452 91924
rect 241948 91644 242004 91700
rect 243068 91308 243124 91364
rect 242060 90188 242116 90244
rect 41132 89852 41188 89908
rect 57036 89852 57092 89908
rect 243180 89628 243236 89684
rect 241948 89068 242004 89124
rect 29484 88060 29540 88116
rect 242172 87948 242228 88004
rect 243068 87612 243124 87668
rect 242284 86828 242340 86884
rect 242732 85708 242788 85764
rect 242060 85596 242116 85652
rect 553084 85484 553140 85540
rect 12572 84812 12628 84868
rect 56252 84812 56308 84868
rect 244524 84588 244580 84644
rect 57036 84252 57092 84308
rect 241948 83580 242004 83636
rect 274764 83468 274820 83524
rect 243180 82348 243236 82404
rect 242172 81564 242228 81620
rect 243292 81228 243348 81284
rect 9324 80444 9380 80500
rect 243068 80108 243124 80164
rect 242284 79548 242340 79604
rect 4396 79100 4452 79156
rect 242844 78988 242900 79044
rect 242956 77868 243012 77924
rect 242732 77532 242788 77588
rect 275548 76748 275604 76804
rect 56252 76636 56308 76692
rect 274652 75628 274708 75684
rect 549500 75628 549556 75684
rect 244524 75516 244580 75572
rect 242732 74508 242788 74564
rect 274764 73500 274820 73556
rect 244524 73052 244580 73108
rect 275548 73052 275604 73108
rect 10892 72828 10948 72884
rect 243180 71484 243236 71540
rect 243292 69468 243348 69524
rect 4172 69020 4228 69076
rect 14252 68012 14308 68068
rect 55468 68012 55524 68068
rect 243068 67452 243124 67508
rect 553196 65772 553252 65828
rect 349916 65548 349972 65604
rect 242844 65436 242900 65492
rect 55468 65212 55524 65268
rect 4172 64988 4228 65044
rect 242956 63420 243012 63476
rect 4284 61404 4340 61460
rect 244524 61404 244580 61460
rect 591052 60396 591108 60452
rect 593404 60396 593460 60452
rect 591164 60284 591220 60340
rect 593516 60284 593572 60340
rect 591388 60172 591444 60228
rect 550060 59948 550116 60004
rect 5852 59612 5908 59668
rect 57036 59612 57092 59668
rect 274652 59388 274708 59444
rect 57036 57596 57092 57652
rect 242732 57372 242788 57428
rect 552748 55916 552804 55972
rect 343980 55356 344036 55412
rect 549388 54348 549444 54404
rect 4396 53788 4452 53844
rect 350588 53340 350644 53396
rect 593292 53228 593348 53284
rect 350476 51996 350532 52052
rect 549388 51660 549444 51716
rect 350140 51324 350196 51380
rect 5068 50876 5124 50932
rect 4172 49980 4228 50036
rect 549388 49756 549444 49812
rect 242956 49308 243012 49364
rect 549276 48636 549332 48692
rect 350364 48412 350420 48468
rect 5068 47852 5124 47908
rect 57036 47852 57092 47908
rect 343532 47292 343588 47348
rect 57036 46172 57092 46228
rect 349916 45388 349972 45444
rect 349580 45276 349636 45332
rect 241948 43260 242004 43316
rect 4172 42364 4228 42420
rect 548940 42252 548996 42308
rect 549276 42252 549332 42308
rect 551068 42252 551124 42308
rect 496300 41468 496356 41524
rect 483868 41244 483924 41300
rect 488236 41244 488292 41300
rect 553980 41244 554036 41300
rect 480172 41132 480228 41188
rect 593516 40908 593572 40964
rect 431788 40684 431844 40740
rect 436268 40460 436324 40516
rect 554428 40460 554484 40516
rect 461132 40348 461188 40404
rect 554652 40236 554708 40292
rect 553532 39900 553588 39956
rect 419692 39676 419748 39732
rect 480172 39676 480228 39732
rect 483868 39676 483924 39732
rect 488236 39676 488292 39732
rect 496300 39676 496356 39732
rect 516460 39676 516516 39732
rect 532700 39676 532756 39732
rect 347004 39452 347060 39508
rect 451948 39452 452004 39508
rect 460012 39340 460068 39396
rect 437612 39228 437668 39284
rect 554652 39228 554708 39284
rect 4284 38556 4340 38612
rect 524524 38556 524580 38612
rect 524972 38556 525028 38612
rect 548828 38332 548884 38388
rect 347004 38220 347060 38276
rect 532588 37996 532644 38052
rect 550844 37996 550900 38052
rect 546028 37884 546084 37940
rect 354508 37660 354564 37716
rect 478828 37660 478884 37716
rect 483868 37660 483924 37716
rect 487228 37660 487284 37716
rect 554540 37548 554596 37604
rect 463708 37324 463764 37380
rect 362908 36988 362964 37044
rect 383852 36988 383908 37044
rect 500332 36988 500388 37044
rect 504812 36988 504868 37044
rect 512428 36988 512484 37044
rect 528556 36988 528612 37044
rect 4172 36876 4228 36932
rect 347228 36876 347284 36932
rect 241948 36764 242004 36820
rect 549500 36764 549556 36820
rect 242956 36652 243012 36708
rect 549612 36652 549668 36708
rect 343532 36540 343588 36596
rect 552972 36540 553028 36596
rect 343980 36428 344036 36484
rect 349580 36316 349636 36372
rect 553084 36316 553140 36372
rect 554316 36204 554372 36260
rect 423388 35308 423444 35364
rect 350140 35196 350196 35252
rect 553196 35196 553252 35252
rect 350588 34972 350644 35028
rect 552748 34972 552804 35028
rect 349916 34860 349972 34916
rect 4172 34748 4228 34804
rect 437612 34748 437668 34804
rect 553420 34748 553476 34804
rect 461132 34636 461188 34692
rect 553308 34636 553364 34692
rect 519148 34524 519204 34580
rect 528556 34412 528612 34468
rect 550172 34412 550228 34468
rect 350364 33516 350420 33572
rect 105084 32956 105140 33012
rect 81788 32844 81844 32900
rect 151676 32732 151732 32788
rect 223580 32620 223636 32676
rect 191100 32508 191156 32564
rect 194124 32396 194180 32452
rect 209916 31500 209972 31556
rect 200060 31388 200116 31444
rect 223580 31388 223636 31444
rect 198268 31276 198324 31332
rect 196476 31164 196532 31220
rect 188412 30828 188468 30884
rect 139132 30716 139188 30772
rect 140924 30716 140980 30772
rect 142716 30716 142772 30772
rect 149884 30716 149940 30772
rect 151676 30604 151732 30660
rect 153468 30604 153524 30660
rect 158844 30604 158900 30660
rect 160636 30604 160692 30660
rect 162428 30604 162484 30660
rect 191100 30604 191156 30660
rect 196476 30604 196532 30660
rect 198268 30604 198324 30660
rect 200060 30604 200116 30660
rect 105084 30268 105140 30324
rect 81788 30044 81844 30100
rect 554540 30044 554596 30100
rect 147868 29708 147924 29764
rect 157052 29708 157108 29764
rect 188412 29708 188468 29764
rect 221564 29596 221620 29652
rect 394828 29596 394884 29652
rect 371308 28588 371364 28644
rect 593292 28588 593348 28644
rect 110460 28476 110516 28532
rect 112252 28476 112308 28532
rect 137788 28476 137844 28532
rect 139132 28476 139188 28532
rect 139580 28476 139636 28532
rect 140924 28476 140980 28532
rect 141148 28476 141204 28532
rect 142716 28476 142772 28532
rect 194124 28476 194180 28532
rect 209916 28476 209972 28532
rect 215852 28476 215908 28532
rect 219884 28476 219940 28532
rect 220108 28476 220164 28532
rect 221564 28476 221620 28532
rect 346108 28476 346164 28532
rect 347676 28476 347732 28532
rect 140812 28364 140868 28420
rect 347452 28364 347508 28420
rect 155260 28252 155316 28308
rect 347564 28252 347620 28308
rect 346108 28140 346164 28196
rect 158844 27916 158900 27972
rect 186508 27916 186564 27972
rect 346892 27804 346948 27860
rect 552300 27692 552356 27748
rect 203308 27580 203364 27636
rect 238476 27580 238532 27636
rect 80668 27356 80724 27412
rect 104188 27356 104244 27412
rect 159628 27356 159684 27412
rect 161420 27356 161476 27412
rect 347340 27356 347396 27412
rect 551516 27020 551572 27076
rect 73836 26908 73892 26964
rect 147868 26908 147924 26964
rect 156268 26908 156324 26964
rect 551292 26908 551348 26964
rect 552076 26908 552132 26964
rect 144508 26572 144564 26628
rect 346780 26348 346836 26404
rect 554540 26348 554596 26404
rect 347116 26236 347172 26292
rect 144508 26012 144564 26068
rect 554428 25788 554484 25844
rect 554540 25452 554596 25508
rect 155260 24556 155316 24612
rect 349916 24556 349972 24612
rect 347004 24444 347060 24500
rect 548604 23100 548660 23156
rect 4284 22876 4340 22932
rect 350476 21644 350532 21700
rect 548940 21644 548996 21700
rect 209356 21532 209412 21588
rect 548716 21420 548772 21476
rect 158844 21308 158900 21364
rect 548492 21308 548548 21364
rect 218428 21196 218484 21252
rect 350364 20860 350420 20916
rect 137788 19740 137844 19796
rect 149884 19516 149940 19572
rect 159628 17612 159684 17668
rect 350476 17500 350532 17556
rect 141148 16268 141204 16324
rect 593404 16268 593460 16324
rect 161420 16044 161476 16100
rect 551852 15372 551908 15428
rect 156268 14476 156324 14532
rect 147868 12796 147924 12852
rect 215852 12684 215908 12740
rect 552524 12684 552580 12740
rect 220108 10892 220164 10948
rect 557340 10556 557396 10612
rect 557564 10556 557620 10612
rect 574476 10556 574532 10612
rect 586012 10556 586068 10612
rect 591388 10556 591444 10612
rect 557452 10444 557508 10500
rect 559356 10444 559412 10500
rect 574364 10444 574420 10500
rect 557116 10332 557172 10388
rect 558012 10332 558068 10388
rect 560028 10332 560084 10388
rect 579964 10332 580020 10388
rect 557676 10220 557732 10276
rect 554652 10108 554708 10164
rect 558012 10108 558068 10164
rect 557004 9884 557060 9940
rect 570108 9884 570164 9940
rect 575372 9884 575428 9940
rect 586348 9772 586404 9828
rect 556892 9660 556948 9716
rect 584668 9660 584724 9716
rect 574588 9548 574644 9604
rect 581308 9548 581364 9604
rect 576268 9324 576324 9380
rect 579852 9212 579908 9268
rect 549052 9100 549108 9156
rect 4172 8764 4228 8820
rect 572908 8316 572964 8372
rect 575036 8316 575092 8372
rect 577052 8204 577108 8260
rect 571228 8092 571284 8148
rect 577948 8092 578004 8148
rect 578844 8092 578900 8148
rect 579852 8092 579908 8148
rect 549052 7980 549108 8036
rect 569996 7980 570052 8036
rect 551068 7868 551124 7924
rect 571116 7868 571172 7924
rect 569884 7644 569940 7700
rect 571340 7644 571396 7700
rect 80668 7532 80724 7588
rect 571340 7196 571396 7252
rect 573244 7084 573300 7140
rect 569996 6972 570052 7028
rect 574476 6860 574532 6916
rect 571228 6748 571284 6804
rect 577164 6748 577220 6804
rect 139580 6188 139636 6244
rect 571116 6188 571172 6244
rect 572796 6076 572852 6132
rect 574364 5964 574420 6020
rect 104188 5852 104244 5908
rect 574476 5852 574532 5908
rect 550956 4956 551012 5012
rect 571004 252 571060 308
rect 572684 140 572740 196
rect 572572 28 572628 84
<< metal4 >>
rect -1916 598172 -1296 598268
rect -1916 598116 -1820 598172
rect -1764 598116 -1696 598172
rect -1640 598116 -1572 598172
rect -1516 598116 -1448 598172
rect -1392 598116 -1296 598172
rect -1916 598048 -1296 598116
rect -1916 597992 -1820 598048
rect -1764 597992 -1696 598048
rect -1640 597992 -1572 598048
rect -1516 597992 -1448 598048
rect -1392 597992 -1296 598048
rect -1916 597924 -1296 597992
rect -1916 597868 -1820 597924
rect -1764 597868 -1696 597924
rect -1640 597868 -1572 597924
rect -1516 597868 -1448 597924
rect -1392 597868 -1296 597924
rect -1916 597800 -1296 597868
rect -1916 597744 -1820 597800
rect -1764 597744 -1696 597800
rect -1640 597744 -1572 597800
rect -1516 597744 -1448 597800
rect -1392 597744 -1296 597800
rect -1916 586350 -1296 597744
rect -1916 586294 -1820 586350
rect -1764 586294 -1696 586350
rect -1640 586294 -1572 586350
rect -1516 586294 -1448 586350
rect -1392 586294 -1296 586350
rect -1916 586226 -1296 586294
rect -1916 586170 -1820 586226
rect -1764 586170 -1696 586226
rect -1640 586170 -1572 586226
rect -1516 586170 -1448 586226
rect -1392 586170 -1296 586226
rect -1916 586102 -1296 586170
rect -1916 586046 -1820 586102
rect -1764 586046 -1696 586102
rect -1640 586046 -1572 586102
rect -1516 586046 -1448 586102
rect -1392 586046 -1296 586102
rect -1916 585978 -1296 586046
rect -1916 585922 -1820 585978
rect -1764 585922 -1696 585978
rect -1640 585922 -1572 585978
rect -1516 585922 -1448 585978
rect -1392 585922 -1296 585978
rect -1916 568350 -1296 585922
rect -1916 568294 -1820 568350
rect -1764 568294 -1696 568350
rect -1640 568294 -1572 568350
rect -1516 568294 -1448 568350
rect -1392 568294 -1296 568350
rect -1916 568226 -1296 568294
rect -1916 568170 -1820 568226
rect -1764 568170 -1696 568226
rect -1640 568170 -1572 568226
rect -1516 568170 -1448 568226
rect -1392 568170 -1296 568226
rect -1916 568102 -1296 568170
rect -1916 568046 -1820 568102
rect -1764 568046 -1696 568102
rect -1640 568046 -1572 568102
rect -1516 568046 -1448 568102
rect -1392 568046 -1296 568102
rect -1916 567978 -1296 568046
rect -1916 567922 -1820 567978
rect -1764 567922 -1696 567978
rect -1640 567922 -1572 567978
rect -1516 567922 -1448 567978
rect -1392 567922 -1296 567978
rect -1916 550350 -1296 567922
rect -1916 550294 -1820 550350
rect -1764 550294 -1696 550350
rect -1640 550294 -1572 550350
rect -1516 550294 -1448 550350
rect -1392 550294 -1296 550350
rect -1916 550226 -1296 550294
rect -1916 550170 -1820 550226
rect -1764 550170 -1696 550226
rect -1640 550170 -1572 550226
rect -1516 550170 -1448 550226
rect -1392 550170 -1296 550226
rect -1916 550102 -1296 550170
rect -1916 550046 -1820 550102
rect -1764 550046 -1696 550102
rect -1640 550046 -1572 550102
rect -1516 550046 -1448 550102
rect -1392 550046 -1296 550102
rect -1916 549978 -1296 550046
rect -1916 549922 -1820 549978
rect -1764 549922 -1696 549978
rect -1640 549922 -1572 549978
rect -1516 549922 -1448 549978
rect -1392 549922 -1296 549978
rect -1916 532350 -1296 549922
rect -1916 532294 -1820 532350
rect -1764 532294 -1696 532350
rect -1640 532294 -1572 532350
rect -1516 532294 -1448 532350
rect -1392 532294 -1296 532350
rect -1916 532226 -1296 532294
rect -1916 532170 -1820 532226
rect -1764 532170 -1696 532226
rect -1640 532170 -1572 532226
rect -1516 532170 -1448 532226
rect -1392 532170 -1296 532226
rect -1916 532102 -1296 532170
rect -1916 532046 -1820 532102
rect -1764 532046 -1696 532102
rect -1640 532046 -1572 532102
rect -1516 532046 -1448 532102
rect -1392 532046 -1296 532102
rect -1916 531978 -1296 532046
rect -1916 531922 -1820 531978
rect -1764 531922 -1696 531978
rect -1640 531922 -1572 531978
rect -1516 531922 -1448 531978
rect -1392 531922 -1296 531978
rect -1916 514350 -1296 531922
rect -1916 514294 -1820 514350
rect -1764 514294 -1696 514350
rect -1640 514294 -1572 514350
rect -1516 514294 -1448 514350
rect -1392 514294 -1296 514350
rect -1916 514226 -1296 514294
rect -1916 514170 -1820 514226
rect -1764 514170 -1696 514226
rect -1640 514170 -1572 514226
rect -1516 514170 -1448 514226
rect -1392 514170 -1296 514226
rect -1916 514102 -1296 514170
rect -1916 514046 -1820 514102
rect -1764 514046 -1696 514102
rect -1640 514046 -1572 514102
rect -1516 514046 -1448 514102
rect -1392 514046 -1296 514102
rect -1916 513978 -1296 514046
rect -1916 513922 -1820 513978
rect -1764 513922 -1696 513978
rect -1640 513922 -1572 513978
rect -1516 513922 -1448 513978
rect -1392 513922 -1296 513978
rect -1916 496350 -1296 513922
rect -1916 496294 -1820 496350
rect -1764 496294 -1696 496350
rect -1640 496294 -1572 496350
rect -1516 496294 -1448 496350
rect -1392 496294 -1296 496350
rect -1916 496226 -1296 496294
rect -1916 496170 -1820 496226
rect -1764 496170 -1696 496226
rect -1640 496170 -1572 496226
rect -1516 496170 -1448 496226
rect -1392 496170 -1296 496226
rect -1916 496102 -1296 496170
rect -1916 496046 -1820 496102
rect -1764 496046 -1696 496102
rect -1640 496046 -1572 496102
rect -1516 496046 -1448 496102
rect -1392 496046 -1296 496102
rect -1916 495978 -1296 496046
rect -1916 495922 -1820 495978
rect -1764 495922 -1696 495978
rect -1640 495922 -1572 495978
rect -1516 495922 -1448 495978
rect -1392 495922 -1296 495978
rect -1916 478350 -1296 495922
rect -1916 478294 -1820 478350
rect -1764 478294 -1696 478350
rect -1640 478294 -1572 478350
rect -1516 478294 -1448 478350
rect -1392 478294 -1296 478350
rect -1916 478226 -1296 478294
rect -1916 478170 -1820 478226
rect -1764 478170 -1696 478226
rect -1640 478170 -1572 478226
rect -1516 478170 -1448 478226
rect -1392 478170 -1296 478226
rect -1916 478102 -1296 478170
rect -1916 478046 -1820 478102
rect -1764 478046 -1696 478102
rect -1640 478046 -1572 478102
rect -1516 478046 -1448 478102
rect -1392 478046 -1296 478102
rect -1916 477978 -1296 478046
rect -1916 477922 -1820 477978
rect -1764 477922 -1696 477978
rect -1640 477922 -1572 477978
rect -1516 477922 -1448 477978
rect -1392 477922 -1296 477978
rect -1916 460350 -1296 477922
rect -1916 460294 -1820 460350
rect -1764 460294 -1696 460350
rect -1640 460294 -1572 460350
rect -1516 460294 -1448 460350
rect -1392 460294 -1296 460350
rect -1916 460226 -1296 460294
rect -1916 460170 -1820 460226
rect -1764 460170 -1696 460226
rect -1640 460170 -1572 460226
rect -1516 460170 -1448 460226
rect -1392 460170 -1296 460226
rect -1916 460102 -1296 460170
rect -1916 460046 -1820 460102
rect -1764 460046 -1696 460102
rect -1640 460046 -1572 460102
rect -1516 460046 -1448 460102
rect -1392 460046 -1296 460102
rect -1916 459978 -1296 460046
rect -1916 459922 -1820 459978
rect -1764 459922 -1696 459978
rect -1640 459922 -1572 459978
rect -1516 459922 -1448 459978
rect -1392 459922 -1296 459978
rect -1916 442350 -1296 459922
rect -1916 442294 -1820 442350
rect -1764 442294 -1696 442350
rect -1640 442294 -1572 442350
rect -1516 442294 -1448 442350
rect -1392 442294 -1296 442350
rect -1916 442226 -1296 442294
rect -1916 442170 -1820 442226
rect -1764 442170 -1696 442226
rect -1640 442170 -1572 442226
rect -1516 442170 -1448 442226
rect -1392 442170 -1296 442226
rect -1916 442102 -1296 442170
rect -1916 442046 -1820 442102
rect -1764 442046 -1696 442102
rect -1640 442046 -1572 442102
rect -1516 442046 -1448 442102
rect -1392 442046 -1296 442102
rect -1916 441978 -1296 442046
rect -1916 441922 -1820 441978
rect -1764 441922 -1696 441978
rect -1640 441922 -1572 441978
rect -1516 441922 -1448 441978
rect -1392 441922 -1296 441978
rect -1916 424350 -1296 441922
rect -1916 424294 -1820 424350
rect -1764 424294 -1696 424350
rect -1640 424294 -1572 424350
rect -1516 424294 -1448 424350
rect -1392 424294 -1296 424350
rect -1916 424226 -1296 424294
rect -1916 424170 -1820 424226
rect -1764 424170 -1696 424226
rect -1640 424170 -1572 424226
rect -1516 424170 -1448 424226
rect -1392 424170 -1296 424226
rect -1916 424102 -1296 424170
rect -1916 424046 -1820 424102
rect -1764 424046 -1696 424102
rect -1640 424046 -1572 424102
rect -1516 424046 -1448 424102
rect -1392 424046 -1296 424102
rect -1916 423978 -1296 424046
rect -1916 423922 -1820 423978
rect -1764 423922 -1696 423978
rect -1640 423922 -1572 423978
rect -1516 423922 -1448 423978
rect -1392 423922 -1296 423978
rect -1916 406350 -1296 423922
rect -1916 406294 -1820 406350
rect -1764 406294 -1696 406350
rect -1640 406294 -1572 406350
rect -1516 406294 -1448 406350
rect -1392 406294 -1296 406350
rect -1916 406226 -1296 406294
rect -1916 406170 -1820 406226
rect -1764 406170 -1696 406226
rect -1640 406170 -1572 406226
rect -1516 406170 -1448 406226
rect -1392 406170 -1296 406226
rect -1916 406102 -1296 406170
rect -1916 406046 -1820 406102
rect -1764 406046 -1696 406102
rect -1640 406046 -1572 406102
rect -1516 406046 -1448 406102
rect -1392 406046 -1296 406102
rect -1916 405978 -1296 406046
rect -1916 405922 -1820 405978
rect -1764 405922 -1696 405978
rect -1640 405922 -1572 405978
rect -1516 405922 -1448 405978
rect -1392 405922 -1296 405978
rect -1916 388350 -1296 405922
rect -1916 388294 -1820 388350
rect -1764 388294 -1696 388350
rect -1640 388294 -1572 388350
rect -1516 388294 -1448 388350
rect -1392 388294 -1296 388350
rect -1916 388226 -1296 388294
rect -1916 388170 -1820 388226
rect -1764 388170 -1696 388226
rect -1640 388170 -1572 388226
rect -1516 388170 -1448 388226
rect -1392 388170 -1296 388226
rect -1916 388102 -1296 388170
rect -1916 388046 -1820 388102
rect -1764 388046 -1696 388102
rect -1640 388046 -1572 388102
rect -1516 388046 -1448 388102
rect -1392 388046 -1296 388102
rect -1916 387978 -1296 388046
rect -1916 387922 -1820 387978
rect -1764 387922 -1696 387978
rect -1640 387922 -1572 387978
rect -1516 387922 -1448 387978
rect -1392 387922 -1296 387978
rect -1916 370350 -1296 387922
rect -1916 370294 -1820 370350
rect -1764 370294 -1696 370350
rect -1640 370294 -1572 370350
rect -1516 370294 -1448 370350
rect -1392 370294 -1296 370350
rect -1916 370226 -1296 370294
rect -1916 370170 -1820 370226
rect -1764 370170 -1696 370226
rect -1640 370170 -1572 370226
rect -1516 370170 -1448 370226
rect -1392 370170 -1296 370226
rect -1916 370102 -1296 370170
rect -1916 370046 -1820 370102
rect -1764 370046 -1696 370102
rect -1640 370046 -1572 370102
rect -1516 370046 -1448 370102
rect -1392 370046 -1296 370102
rect -1916 369978 -1296 370046
rect -1916 369922 -1820 369978
rect -1764 369922 -1696 369978
rect -1640 369922 -1572 369978
rect -1516 369922 -1448 369978
rect -1392 369922 -1296 369978
rect -1916 352350 -1296 369922
rect -1916 352294 -1820 352350
rect -1764 352294 -1696 352350
rect -1640 352294 -1572 352350
rect -1516 352294 -1448 352350
rect -1392 352294 -1296 352350
rect -1916 352226 -1296 352294
rect -1916 352170 -1820 352226
rect -1764 352170 -1696 352226
rect -1640 352170 -1572 352226
rect -1516 352170 -1448 352226
rect -1392 352170 -1296 352226
rect -1916 352102 -1296 352170
rect -1916 352046 -1820 352102
rect -1764 352046 -1696 352102
rect -1640 352046 -1572 352102
rect -1516 352046 -1448 352102
rect -1392 352046 -1296 352102
rect -1916 351978 -1296 352046
rect -1916 351922 -1820 351978
rect -1764 351922 -1696 351978
rect -1640 351922 -1572 351978
rect -1516 351922 -1448 351978
rect -1392 351922 -1296 351978
rect -1916 334350 -1296 351922
rect -1916 334294 -1820 334350
rect -1764 334294 -1696 334350
rect -1640 334294 -1572 334350
rect -1516 334294 -1448 334350
rect -1392 334294 -1296 334350
rect -1916 334226 -1296 334294
rect -1916 334170 -1820 334226
rect -1764 334170 -1696 334226
rect -1640 334170 -1572 334226
rect -1516 334170 -1448 334226
rect -1392 334170 -1296 334226
rect -1916 334102 -1296 334170
rect -1916 334046 -1820 334102
rect -1764 334046 -1696 334102
rect -1640 334046 -1572 334102
rect -1516 334046 -1448 334102
rect -1392 334046 -1296 334102
rect -1916 333978 -1296 334046
rect -1916 333922 -1820 333978
rect -1764 333922 -1696 333978
rect -1640 333922 -1572 333978
rect -1516 333922 -1448 333978
rect -1392 333922 -1296 333978
rect -1916 316350 -1296 333922
rect -1916 316294 -1820 316350
rect -1764 316294 -1696 316350
rect -1640 316294 -1572 316350
rect -1516 316294 -1448 316350
rect -1392 316294 -1296 316350
rect -1916 316226 -1296 316294
rect -1916 316170 -1820 316226
rect -1764 316170 -1696 316226
rect -1640 316170 -1572 316226
rect -1516 316170 -1448 316226
rect -1392 316170 -1296 316226
rect -1916 316102 -1296 316170
rect -1916 316046 -1820 316102
rect -1764 316046 -1696 316102
rect -1640 316046 -1572 316102
rect -1516 316046 -1448 316102
rect -1392 316046 -1296 316102
rect -1916 315978 -1296 316046
rect -1916 315922 -1820 315978
rect -1764 315922 -1696 315978
rect -1640 315922 -1572 315978
rect -1516 315922 -1448 315978
rect -1392 315922 -1296 315978
rect -1916 298350 -1296 315922
rect -1916 298294 -1820 298350
rect -1764 298294 -1696 298350
rect -1640 298294 -1572 298350
rect -1516 298294 -1448 298350
rect -1392 298294 -1296 298350
rect -1916 298226 -1296 298294
rect -1916 298170 -1820 298226
rect -1764 298170 -1696 298226
rect -1640 298170 -1572 298226
rect -1516 298170 -1448 298226
rect -1392 298170 -1296 298226
rect -1916 298102 -1296 298170
rect -1916 298046 -1820 298102
rect -1764 298046 -1696 298102
rect -1640 298046 -1572 298102
rect -1516 298046 -1448 298102
rect -1392 298046 -1296 298102
rect -1916 297978 -1296 298046
rect -1916 297922 -1820 297978
rect -1764 297922 -1696 297978
rect -1640 297922 -1572 297978
rect -1516 297922 -1448 297978
rect -1392 297922 -1296 297978
rect -1916 280350 -1296 297922
rect -1916 280294 -1820 280350
rect -1764 280294 -1696 280350
rect -1640 280294 -1572 280350
rect -1516 280294 -1448 280350
rect -1392 280294 -1296 280350
rect -1916 280226 -1296 280294
rect -1916 280170 -1820 280226
rect -1764 280170 -1696 280226
rect -1640 280170 -1572 280226
rect -1516 280170 -1448 280226
rect -1392 280170 -1296 280226
rect -1916 280102 -1296 280170
rect -1916 280046 -1820 280102
rect -1764 280046 -1696 280102
rect -1640 280046 -1572 280102
rect -1516 280046 -1448 280102
rect -1392 280046 -1296 280102
rect -1916 279978 -1296 280046
rect -1916 279922 -1820 279978
rect -1764 279922 -1696 279978
rect -1640 279922 -1572 279978
rect -1516 279922 -1448 279978
rect -1392 279922 -1296 279978
rect -1916 262350 -1296 279922
rect -1916 262294 -1820 262350
rect -1764 262294 -1696 262350
rect -1640 262294 -1572 262350
rect -1516 262294 -1448 262350
rect -1392 262294 -1296 262350
rect -1916 262226 -1296 262294
rect -1916 262170 -1820 262226
rect -1764 262170 -1696 262226
rect -1640 262170 -1572 262226
rect -1516 262170 -1448 262226
rect -1392 262170 -1296 262226
rect -1916 262102 -1296 262170
rect -1916 262046 -1820 262102
rect -1764 262046 -1696 262102
rect -1640 262046 -1572 262102
rect -1516 262046 -1448 262102
rect -1392 262046 -1296 262102
rect -1916 261978 -1296 262046
rect -1916 261922 -1820 261978
rect -1764 261922 -1696 261978
rect -1640 261922 -1572 261978
rect -1516 261922 -1448 261978
rect -1392 261922 -1296 261978
rect -1916 244350 -1296 261922
rect -1916 244294 -1820 244350
rect -1764 244294 -1696 244350
rect -1640 244294 -1572 244350
rect -1516 244294 -1448 244350
rect -1392 244294 -1296 244350
rect -1916 244226 -1296 244294
rect -1916 244170 -1820 244226
rect -1764 244170 -1696 244226
rect -1640 244170 -1572 244226
rect -1516 244170 -1448 244226
rect -1392 244170 -1296 244226
rect -1916 244102 -1296 244170
rect -1916 244046 -1820 244102
rect -1764 244046 -1696 244102
rect -1640 244046 -1572 244102
rect -1516 244046 -1448 244102
rect -1392 244046 -1296 244102
rect -1916 243978 -1296 244046
rect -1916 243922 -1820 243978
rect -1764 243922 -1696 243978
rect -1640 243922 -1572 243978
rect -1516 243922 -1448 243978
rect -1392 243922 -1296 243978
rect -1916 226350 -1296 243922
rect -1916 226294 -1820 226350
rect -1764 226294 -1696 226350
rect -1640 226294 -1572 226350
rect -1516 226294 -1448 226350
rect -1392 226294 -1296 226350
rect -1916 226226 -1296 226294
rect -1916 226170 -1820 226226
rect -1764 226170 -1696 226226
rect -1640 226170 -1572 226226
rect -1516 226170 -1448 226226
rect -1392 226170 -1296 226226
rect -1916 226102 -1296 226170
rect -1916 226046 -1820 226102
rect -1764 226046 -1696 226102
rect -1640 226046 -1572 226102
rect -1516 226046 -1448 226102
rect -1392 226046 -1296 226102
rect -1916 225978 -1296 226046
rect -1916 225922 -1820 225978
rect -1764 225922 -1696 225978
rect -1640 225922 -1572 225978
rect -1516 225922 -1448 225978
rect -1392 225922 -1296 225978
rect -1916 208350 -1296 225922
rect -1916 208294 -1820 208350
rect -1764 208294 -1696 208350
rect -1640 208294 -1572 208350
rect -1516 208294 -1448 208350
rect -1392 208294 -1296 208350
rect -1916 208226 -1296 208294
rect -1916 208170 -1820 208226
rect -1764 208170 -1696 208226
rect -1640 208170 -1572 208226
rect -1516 208170 -1448 208226
rect -1392 208170 -1296 208226
rect -1916 208102 -1296 208170
rect -1916 208046 -1820 208102
rect -1764 208046 -1696 208102
rect -1640 208046 -1572 208102
rect -1516 208046 -1448 208102
rect -1392 208046 -1296 208102
rect -1916 207978 -1296 208046
rect -1916 207922 -1820 207978
rect -1764 207922 -1696 207978
rect -1640 207922 -1572 207978
rect -1516 207922 -1448 207978
rect -1392 207922 -1296 207978
rect -1916 190350 -1296 207922
rect -1916 190294 -1820 190350
rect -1764 190294 -1696 190350
rect -1640 190294 -1572 190350
rect -1516 190294 -1448 190350
rect -1392 190294 -1296 190350
rect -1916 190226 -1296 190294
rect -1916 190170 -1820 190226
rect -1764 190170 -1696 190226
rect -1640 190170 -1572 190226
rect -1516 190170 -1448 190226
rect -1392 190170 -1296 190226
rect -1916 190102 -1296 190170
rect -1916 190046 -1820 190102
rect -1764 190046 -1696 190102
rect -1640 190046 -1572 190102
rect -1516 190046 -1448 190102
rect -1392 190046 -1296 190102
rect -1916 189978 -1296 190046
rect -1916 189922 -1820 189978
rect -1764 189922 -1696 189978
rect -1640 189922 -1572 189978
rect -1516 189922 -1448 189978
rect -1392 189922 -1296 189978
rect -1916 172350 -1296 189922
rect -1916 172294 -1820 172350
rect -1764 172294 -1696 172350
rect -1640 172294 -1572 172350
rect -1516 172294 -1448 172350
rect -1392 172294 -1296 172350
rect -1916 172226 -1296 172294
rect -1916 172170 -1820 172226
rect -1764 172170 -1696 172226
rect -1640 172170 -1572 172226
rect -1516 172170 -1448 172226
rect -1392 172170 -1296 172226
rect -1916 172102 -1296 172170
rect -1916 172046 -1820 172102
rect -1764 172046 -1696 172102
rect -1640 172046 -1572 172102
rect -1516 172046 -1448 172102
rect -1392 172046 -1296 172102
rect -1916 171978 -1296 172046
rect -1916 171922 -1820 171978
rect -1764 171922 -1696 171978
rect -1640 171922 -1572 171978
rect -1516 171922 -1448 171978
rect -1392 171922 -1296 171978
rect -1916 154350 -1296 171922
rect -1916 154294 -1820 154350
rect -1764 154294 -1696 154350
rect -1640 154294 -1572 154350
rect -1516 154294 -1448 154350
rect -1392 154294 -1296 154350
rect -1916 154226 -1296 154294
rect -1916 154170 -1820 154226
rect -1764 154170 -1696 154226
rect -1640 154170 -1572 154226
rect -1516 154170 -1448 154226
rect -1392 154170 -1296 154226
rect -1916 154102 -1296 154170
rect -1916 154046 -1820 154102
rect -1764 154046 -1696 154102
rect -1640 154046 -1572 154102
rect -1516 154046 -1448 154102
rect -1392 154046 -1296 154102
rect -1916 153978 -1296 154046
rect -1916 153922 -1820 153978
rect -1764 153922 -1696 153978
rect -1640 153922 -1572 153978
rect -1516 153922 -1448 153978
rect -1392 153922 -1296 153978
rect -1916 136350 -1296 153922
rect -1916 136294 -1820 136350
rect -1764 136294 -1696 136350
rect -1640 136294 -1572 136350
rect -1516 136294 -1448 136350
rect -1392 136294 -1296 136350
rect -1916 136226 -1296 136294
rect -1916 136170 -1820 136226
rect -1764 136170 -1696 136226
rect -1640 136170 -1572 136226
rect -1516 136170 -1448 136226
rect -1392 136170 -1296 136226
rect -1916 136102 -1296 136170
rect -1916 136046 -1820 136102
rect -1764 136046 -1696 136102
rect -1640 136046 -1572 136102
rect -1516 136046 -1448 136102
rect -1392 136046 -1296 136102
rect -1916 135978 -1296 136046
rect -1916 135922 -1820 135978
rect -1764 135922 -1696 135978
rect -1640 135922 -1572 135978
rect -1516 135922 -1448 135978
rect -1392 135922 -1296 135978
rect -1916 118350 -1296 135922
rect -1916 118294 -1820 118350
rect -1764 118294 -1696 118350
rect -1640 118294 -1572 118350
rect -1516 118294 -1448 118350
rect -1392 118294 -1296 118350
rect -1916 118226 -1296 118294
rect -1916 118170 -1820 118226
rect -1764 118170 -1696 118226
rect -1640 118170 -1572 118226
rect -1516 118170 -1448 118226
rect -1392 118170 -1296 118226
rect -1916 118102 -1296 118170
rect -1916 118046 -1820 118102
rect -1764 118046 -1696 118102
rect -1640 118046 -1572 118102
rect -1516 118046 -1448 118102
rect -1392 118046 -1296 118102
rect -1916 117978 -1296 118046
rect -1916 117922 -1820 117978
rect -1764 117922 -1696 117978
rect -1640 117922 -1572 117978
rect -1516 117922 -1448 117978
rect -1392 117922 -1296 117978
rect -1916 100350 -1296 117922
rect -1916 100294 -1820 100350
rect -1764 100294 -1696 100350
rect -1640 100294 -1572 100350
rect -1516 100294 -1448 100350
rect -1392 100294 -1296 100350
rect -1916 100226 -1296 100294
rect -1916 100170 -1820 100226
rect -1764 100170 -1696 100226
rect -1640 100170 -1572 100226
rect -1516 100170 -1448 100226
rect -1392 100170 -1296 100226
rect -1916 100102 -1296 100170
rect -1916 100046 -1820 100102
rect -1764 100046 -1696 100102
rect -1640 100046 -1572 100102
rect -1516 100046 -1448 100102
rect -1392 100046 -1296 100102
rect -1916 99978 -1296 100046
rect -1916 99922 -1820 99978
rect -1764 99922 -1696 99978
rect -1640 99922 -1572 99978
rect -1516 99922 -1448 99978
rect -1392 99922 -1296 99978
rect -1916 82350 -1296 99922
rect -1916 82294 -1820 82350
rect -1764 82294 -1696 82350
rect -1640 82294 -1572 82350
rect -1516 82294 -1448 82350
rect -1392 82294 -1296 82350
rect -1916 82226 -1296 82294
rect -1916 82170 -1820 82226
rect -1764 82170 -1696 82226
rect -1640 82170 -1572 82226
rect -1516 82170 -1448 82226
rect -1392 82170 -1296 82226
rect -1916 82102 -1296 82170
rect -1916 82046 -1820 82102
rect -1764 82046 -1696 82102
rect -1640 82046 -1572 82102
rect -1516 82046 -1448 82102
rect -1392 82046 -1296 82102
rect -1916 81978 -1296 82046
rect -1916 81922 -1820 81978
rect -1764 81922 -1696 81978
rect -1640 81922 -1572 81978
rect -1516 81922 -1448 81978
rect -1392 81922 -1296 81978
rect -1916 64350 -1296 81922
rect -1916 64294 -1820 64350
rect -1764 64294 -1696 64350
rect -1640 64294 -1572 64350
rect -1516 64294 -1448 64350
rect -1392 64294 -1296 64350
rect -1916 64226 -1296 64294
rect -1916 64170 -1820 64226
rect -1764 64170 -1696 64226
rect -1640 64170 -1572 64226
rect -1516 64170 -1448 64226
rect -1392 64170 -1296 64226
rect -1916 64102 -1296 64170
rect -1916 64046 -1820 64102
rect -1764 64046 -1696 64102
rect -1640 64046 -1572 64102
rect -1516 64046 -1448 64102
rect -1392 64046 -1296 64102
rect -1916 63978 -1296 64046
rect -1916 63922 -1820 63978
rect -1764 63922 -1696 63978
rect -1640 63922 -1572 63978
rect -1516 63922 -1448 63978
rect -1392 63922 -1296 63978
rect -1916 46350 -1296 63922
rect -1916 46294 -1820 46350
rect -1764 46294 -1696 46350
rect -1640 46294 -1572 46350
rect -1516 46294 -1448 46350
rect -1392 46294 -1296 46350
rect -1916 46226 -1296 46294
rect -1916 46170 -1820 46226
rect -1764 46170 -1696 46226
rect -1640 46170 -1572 46226
rect -1516 46170 -1448 46226
rect -1392 46170 -1296 46226
rect -1916 46102 -1296 46170
rect -1916 46046 -1820 46102
rect -1764 46046 -1696 46102
rect -1640 46046 -1572 46102
rect -1516 46046 -1448 46102
rect -1392 46046 -1296 46102
rect -1916 45978 -1296 46046
rect -1916 45922 -1820 45978
rect -1764 45922 -1696 45978
rect -1640 45922 -1572 45978
rect -1516 45922 -1448 45978
rect -1392 45922 -1296 45978
rect -1916 28350 -1296 45922
rect -1916 28294 -1820 28350
rect -1764 28294 -1696 28350
rect -1640 28294 -1572 28350
rect -1516 28294 -1448 28350
rect -1392 28294 -1296 28350
rect -1916 28226 -1296 28294
rect -1916 28170 -1820 28226
rect -1764 28170 -1696 28226
rect -1640 28170 -1572 28226
rect -1516 28170 -1448 28226
rect -1392 28170 -1296 28226
rect -1916 28102 -1296 28170
rect -1916 28046 -1820 28102
rect -1764 28046 -1696 28102
rect -1640 28046 -1572 28102
rect -1516 28046 -1448 28102
rect -1392 28046 -1296 28102
rect -1916 27978 -1296 28046
rect -1916 27922 -1820 27978
rect -1764 27922 -1696 27978
rect -1640 27922 -1572 27978
rect -1516 27922 -1448 27978
rect -1392 27922 -1296 27978
rect -1916 10350 -1296 27922
rect -1916 10294 -1820 10350
rect -1764 10294 -1696 10350
rect -1640 10294 -1572 10350
rect -1516 10294 -1448 10350
rect -1392 10294 -1296 10350
rect -1916 10226 -1296 10294
rect -1916 10170 -1820 10226
rect -1764 10170 -1696 10226
rect -1640 10170 -1572 10226
rect -1516 10170 -1448 10226
rect -1392 10170 -1296 10226
rect -1916 10102 -1296 10170
rect -1916 10046 -1820 10102
rect -1764 10046 -1696 10102
rect -1640 10046 -1572 10102
rect -1516 10046 -1448 10102
rect -1392 10046 -1296 10102
rect -1916 9978 -1296 10046
rect -1916 9922 -1820 9978
rect -1764 9922 -1696 9978
rect -1640 9922 -1572 9978
rect -1516 9922 -1448 9978
rect -1392 9922 -1296 9978
rect -1916 -1120 -1296 9922
rect -956 597212 -336 597308
rect -956 597156 -860 597212
rect -804 597156 -736 597212
rect -680 597156 -612 597212
rect -556 597156 -488 597212
rect -432 597156 -336 597212
rect -956 597088 -336 597156
rect -956 597032 -860 597088
rect -804 597032 -736 597088
rect -680 597032 -612 597088
rect -556 597032 -488 597088
rect -432 597032 -336 597088
rect -956 596964 -336 597032
rect -956 596908 -860 596964
rect -804 596908 -736 596964
rect -680 596908 -612 596964
rect -556 596908 -488 596964
rect -432 596908 -336 596964
rect -956 596840 -336 596908
rect -956 596784 -860 596840
rect -804 596784 -736 596840
rect -680 596784 -612 596840
rect -556 596784 -488 596840
rect -432 596784 -336 596840
rect -956 580350 -336 596784
rect -956 580294 -860 580350
rect -804 580294 -736 580350
rect -680 580294 -612 580350
rect -556 580294 -488 580350
rect -432 580294 -336 580350
rect -956 580226 -336 580294
rect -956 580170 -860 580226
rect -804 580170 -736 580226
rect -680 580170 -612 580226
rect -556 580170 -488 580226
rect -432 580170 -336 580226
rect -956 580102 -336 580170
rect -956 580046 -860 580102
rect -804 580046 -736 580102
rect -680 580046 -612 580102
rect -556 580046 -488 580102
rect -432 580046 -336 580102
rect -956 579978 -336 580046
rect -956 579922 -860 579978
rect -804 579922 -736 579978
rect -680 579922 -612 579978
rect -556 579922 -488 579978
rect -432 579922 -336 579978
rect -956 562350 -336 579922
rect -956 562294 -860 562350
rect -804 562294 -736 562350
rect -680 562294 -612 562350
rect -556 562294 -488 562350
rect -432 562294 -336 562350
rect -956 562226 -336 562294
rect -956 562170 -860 562226
rect -804 562170 -736 562226
rect -680 562170 -612 562226
rect -556 562170 -488 562226
rect -432 562170 -336 562226
rect -956 562102 -336 562170
rect -956 562046 -860 562102
rect -804 562046 -736 562102
rect -680 562046 -612 562102
rect -556 562046 -488 562102
rect -432 562046 -336 562102
rect -956 561978 -336 562046
rect -956 561922 -860 561978
rect -804 561922 -736 561978
rect -680 561922 -612 561978
rect -556 561922 -488 561978
rect -432 561922 -336 561978
rect -956 544350 -336 561922
rect -956 544294 -860 544350
rect -804 544294 -736 544350
rect -680 544294 -612 544350
rect -556 544294 -488 544350
rect -432 544294 -336 544350
rect -956 544226 -336 544294
rect -956 544170 -860 544226
rect -804 544170 -736 544226
rect -680 544170 -612 544226
rect -556 544170 -488 544226
rect -432 544170 -336 544226
rect -956 544102 -336 544170
rect -956 544046 -860 544102
rect -804 544046 -736 544102
rect -680 544046 -612 544102
rect -556 544046 -488 544102
rect -432 544046 -336 544102
rect -956 543978 -336 544046
rect -956 543922 -860 543978
rect -804 543922 -736 543978
rect -680 543922 -612 543978
rect -556 543922 -488 543978
rect -432 543922 -336 543978
rect -956 526350 -336 543922
rect -956 526294 -860 526350
rect -804 526294 -736 526350
rect -680 526294 -612 526350
rect -556 526294 -488 526350
rect -432 526294 -336 526350
rect -956 526226 -336 526294
rect -956 526170 -860 526226
rect -804 526170 -736 526226
rect -680 526170 -612 526226
rect -556 526170 -488 526226
rect -432 526170 -336 526226
rect -956 526102 -336 526170
rect -956 526046 -860 526102
rect -804 526046 -736 526102
rect -680 526046 -612 526102
rect -556 526046 -488 526102
rect -432 526046 -336 526102
rect -956 525978 -336 526046
rect -956 525922 -860 525978
rect -804 525922 -736 525978
rect -680 525922 -612 525978
rect -556 525922 -488 525978
rect -432 525922 -336 525978
rect -956 508350 -336 525922
rect -956 508294 -860 508350
rect -804 508294 -736 508350
rect -680 508294 -612 508350
rect -556 508294 -488 508350
rect -432 508294 -336 508350
rect -956 508226 -336 508294
rect -956 508170 -860 508226
rect -804 508170 -736 508226
rect -680 508170 -612 508226
rect -556 508170 -488 508226
rect -432 508170 -336 508226
rect -956 508102 -336 508170
rect -956 508046 -860 508102
rect -804 508046 -736 508102
rect -680 508046 -612 508102
rect -556 508046 -488 508102
rect -432 508046 -336 508102
rect -956 507978 -336 508046
rect -956 507922 -860 507978
rect -804 507922 -736 507978
rect -680 507922 -612 507978
rect -556 507922 -488 507978
rect -432 507922 -336 507978
rect -956 490350 -336 507922
rect -956 490294 -860 490350
rect -804 490294 -736 490350
rect -680 490294 -612 490350
rect -556 490294 -488 490350
rect -432 490294 -336 490350
rect -956 490226 -336 490294
rect -956 490170 -860 490226
rect -804 490170 -736 490226
rect -680 490170 -612 490226
rect -556 490170 -488 490226
rect -432 490170 -336 490226
rect -956 490102 -336 490170
rect -956 490046 -860 490102
rect -804 490046 -736 490102
rect -680 490046 -612 490102
rect -556 490046 -488 490102
rect -432 490046 -336 490102
rect -956 489978 -336 490046
rect -956 489922 -860 489978
rect -804 489922 -736 489978
rect -680 489922 -612 489978
rect -556 489922 -488 489978
rect -432 489922 -336 489978
rect -956 472350 -336 489922
rect -956 472294 -860 472350
rect -804 472294 -736 472350
rect -680 472294 -612 472350
rect -556 472294 -488 472350
rect -432 472294 -336 472350
rect -956 472226 -336 472294
rect -956 472170 -860 472226
rect -804 472170 -736 472226
rect -680 472170 -612 472226
rect -556 472170 -488 472226
rect -432 472170 -336 472226
rect -956 472102 -336 472170
rect -956 472046 -860 472102
rect -804 472046 -736 472102
rect -680 472046 -612 472102
rect -556 472046 -488 472102
rect -432 472046 -336 472102
rect -956 471978 -336 472046
rect -956 471922 -860 471978
rect -804 471922 -736 471978
rect -680 471922 -612 471978
rect -556 471922 -488 471978
rect -432 471922 -336 471978
rect -956 454350 -336 471922
rect -956 454294 -860 454350
rect -804 454294 -736 454350
rect -680 454294 -612 454350
rect -556 454294 -488 454350
rect -432 454294 -336 454350
rect -956 454226 -336 454294
rect -956 454170 -860 454226
rect -804 454170 -736 454226
rect -680 454170 -612 454226
rect -556 454170 -488 454226
rect -432 454170 -336 454226
rect -956 454102 -336 454170
rect -956 454046 -860 454102
rect -804 454046 -736 454102
rect -680 454046 -612 454102
rect -556 454046 -488 454102
rect -432 454046 -336 454102
rect -956 453978 -336 454046
rect -956 453922 -860 453978
rect -804 453922 -736 453978
rect -680 453922 -612 453978
rect -556 453922 -488 453978
rect -432 453922 -336 453978
rect -956 436350 -336 453922
rect -956 436294 -860 436350
rect -804 436294 -736 436350
rect -680 436294 -612 436350
rect -556 436294 -488 436350
rect -432 436294 -336 436350
rect -956 436226 -336 436294
rect -956 436170 -860 436226
rect -804 436170 -736 436226
rect -680 436170 -612 436226
rect -556 436170 -488 436226
rect -432 436170 -336 436226
rect -956 436102 -336 436170
rect -956 436046 -860 436102
rect -804 436046 -736 436102
rect -680 436046 -612 436102
rect -556 436046 -488 436102
rect -432 436046 -336 436102
rect -956 435978 -336 436046
rect -956 435922 -860 435978
rect -804 435922 -736 435978
rect -680 435922 -612 435978
rect -556 435922 -488 435978
rect -432 435922 -336 435978
rect -956 418350 -336 435922
rect -956 418294 -860 418350
rect -804 418294 -736 418350
rect -680 418294 -612 418350
rect -556 418294 -488 418350
rect -432 418294 -336 418350
rect -956 418226 -336 418294
rect -956 418170 -860 418226
rect -804 418170 -736 418226
rect -680 418170 -612 418226
rect -556 418170 -488 418226
rect -432 418170 -336 418226
rect -956 418102 -336 418170
rect -956 418046 -860 418102
rect -804 418046 -736 418102
rect -680 418046 -612 418102
rect -556 418046 -488 418102
rect -432 418046 -336 418102
rect -956 417978 -336 418046
rect -956 417922 -860 417978
rect -804 417922 -736 417978
rect -680 417922 -612 417978
rect -556 417922 -488 417978
rect -432 417922 -336 417978
rect -956 400350 -336 417922
rect -956 400294 -860 400350
rect -804 400294 -736 400350
rect -680 400294 -612 400350
rect -556 400294 -488 400350
rect -432 400294 -336 400350
rect -956 400226 -336 400294
rect -956 400170 -860 400226
rect -804 400170 -736 400226
rect -680 400170 -612 400226
rect -556 400170 -488 400226
rect -432 400170 -336 400226
rect -956 400102 -336 400170
rect -956 400046 -860 400102
rect -804 400046 -736 400102
rect -680 400046 -612 400102
rect -556 400046 -488 400102
rect -432 400046 -336 400102
rect -956 399978 -336 400046
rect -956 399922 -860 399978
rect -804 399922 -736 399978
rect -680 399922 -612 399978
rect -556 399922 -488 399978
rect -432 399922 -336 399978
rect -956 382350 -336 399922
rect -956 382294 -860 382350
rect -804 382294 -736 382350
rect -680 382294 -612 382350
rect -556 382294 -488 382350
rect -432 382294 -336 382350
rect -956 382226 -336 382294
rect -956 382170 -860 382226
rect -804 382170 -736 382226
rect -680 382170 -612 382226
rect -556 382170 -488 382226
rect -432 382170 -336 382226
rect -956 382102 -336 382170
rect -956 382046 -860 382102
rect -804 382046 -736 382102
rect -680 382046 -612 382102
rect -556 382046 -488 382102
rect -432 382046 -336 382102
rect -956 381978 -336 382046
rect -956 381922 -860 381978
rect -804 381922 -736 381978
rect -680 381922 -612 381978
rect -556 381922 -488 381978
rect -432 381922 -336 381978
rect -956 364350 -336 381922
rect -956 364294 -860 364350
rect -804 364294 -736 364350
rect -680 364294 -612 364350
rect -556 364294 -488 364350
rect -432 364294 -336 364350
rect -956 364226 -336 364294
rect -956 364170 -860 364226
rect -804 364170 -736 364226
rect -680 364170 -612 364226
rect -556 364170 -488 364226
rect -432 364170 -336 364226
rect -956 364102 -336 364170
rect -956 364046 -860 364102
rect -804 364046 -736 364102
rect -680 364046 -612 364102
rect -556 364046 -488 364102
rect -432 364046 -336 364102
rect -956 363978 -336 364046
rect -956 363922 -860 363978
rect -804 363922 -736 363978
rect -680 363922 -612 363978
rect -556 363922 -488 363978
rect -432 363922 -336 363978
rect -956 346350 -336 363922
rect -956 346294 -860 346350
rect -804 346294 -736 346350
rect -680 346294 -612 346350
rect -556 346294 -488 346350
rect -432 346294 -336 346350
rect -956 346226 -336 346294
rect -956 346170 -860 346226
rect -804 346170 -736 346226
rect -680 346170 -612 346226
rect -556 346170 -488 346226
rect -432 346170 -336 346226
rect -956 346102 -336 346170
rect -956 346046 -860 346102
rect -804 346046 -736 346102
rect -680 346046 -612 346102
rect -556 346046 -488 346102
rect -432 346046 -336 346102
rect -956 345978 -336 346046
rect -956 345922 -860 345978
rect -804 345922 -736 345978
rect -680 345922 -612 345978
rect -556 345922 -488 345978
rect -432 345922 -336 345978
rect -956 328350 -336 345922
rect -956 328294 -860 328350
rect -804 328294 -736 328350
rect -680 328294 -612 328350
rect -556 328294 -488 328350
rect -432 328294 -336 328350
rect -956 328226 -336 328294
rect -956 328170 -860 328226
rect -804 328170 -736 328226
rect -680 328170 -612 328226
rect -556 328170 -488 328226
rect -432 328170 -336 328226
rect -956 328102 -336 328170
rect -956 328046 -860 328102
rect -804 328046 -736 328102
rect -680 328046 -612 328102
rect -556 328046 -488 328102
rect -432 328046 -336 328102
rect -956 327978 -336 328046
rect -956 327922 -860 327978
rect -804 327922 -736 327978
rect -680 327922 -612 327978
rect -556 327922 -488 327978
rect -432 327922 -336 327978
rect -956 310350 -336 327922
rect -956 310294 -860 310350
rect -804 310294 -736 310350
rect -680 310294 -612 310350
rect -556 310294 -488 310350
rect -432 310294 -336 310350
rect -956 310226 -336 310294
rect -956 310170 -860 310226
rect -804 310170 -736 310226
rect -680 310170 -612 310226
rect -556 310170 -488 310226
rect -432 310170 -336 310226
rect -956 310102 -336 310170
rect -956 310046 -860 310102
rect -804 310046 -736 310102
rect -680 310046 -612 310102
rect -556 310046 -488 310102
rect -432 310046 -336 310102
rect -956 309978 -336 310046
rect -956 309922 -860 309978
rect -804 309922 -736 309978
rect -680 309922 -612 309978
rect -556 309922 -488 309978
rect -432 309922 -336 309978
rect -956 292350 -336 309922
rect -956 292294 -860 292350
rect -804 292294 -736 292350
rect -680 292294 -612 292350
rect -556 292294 -488 292350
rect -432 292294 -336 292350
rect -956 292226 -336 292294
rect -956 292170 -860 292226
rect -804 292170 -736 292226
rect -680 292170 -612 292226
rect -556 292170 -488 292226
rect -432 292170 -336 292226
rect -956 292102 -336 292170
rect -956 292046 -860 292102
rect -804 292046 -736 292102
rect -680 292046 -612 292102
rect -556 292046 -488 292102
rect -432 292046 -336 292102
rect -956 291978 -336 292046
rect -956 291922 -860 291978
rect -804 291922 -736 291978
rect -680 291922 -612 291978
rect -556 291922 -488 291978
rect -432 291922 -336 291978
rect -956 274350 -336 291922
rect -956 274294 -860 274350
rect -804 274294 -736 274350
rect -680 274294 -612 274350
rect -556 274294 -488 274350
rect -432 274294 -336 274350
rect -956 274226 -336 274294
rect -956 274170 -860 274226
rect -804 274170 -736 274226
rect -680 274170 -612 274226
rect -556 274170 -488 274226
rect -432 274170 -336 274226
rect -956 274102 -336 274170
rect -956 274046 -860 274102
rect -804 274046 -736 274102
rect -680 274046 -612 274102
rect -556 274046 -488 274102
rect -432 274046 -336 274102
rect -956 273978 -336 274046
rect -956 273922 -860 273978
rect -804 273922 -736 273978
rect -680 273922 -612 273978
rect -556 273922 -488 273978
rect -432 273922 -336 273978
rect -956 256350 -336 273922
rect -956 256294 -860 256350
rect -804 256294 -736 256350
rect -680 256294 -612 256350
rect -556 256294 -488 256350
rect -432 256294 -336 256350
rect -956 256226 -336 256294
rect -956 256170 -860 256226
rect -804 256170 -736 256226
rect -680 256170 -612 256226
rect -556 256170 -488 256226
rect -432 256170 -336 256226
rect -956 256102 -336 256170
rect -956 256046 -860 256102
rect -804 256046 -736 256102
rect -680 256046 -612 256102
rect -556 256046 -488 256102
rect -432 256046 -336 256102
rect -956 255978 -336 256046
rect -956 255922 -860 255978
rect -804 255922 -736 255978
rect -680 255922 -612 255978
rect -556 255922 -488 255978
rect -432 255922 -336 255978
rect -956 238350 -336 255922
rect -956 238294 -860 238350
rect -804 238294 -736 238350
rect -680 238294 -612 238350
rect -556 238294 -488 238350
rect -432 238294 -336 238350
rect -956 238226 -336 238294
rect -956 238170 -860 238226
rect -804 238170 -736 238226
rect -680 238170 -612 238226
rect -556 238170 -488 238226
rect -432 238170 -336 238226
rect -956 238102 -336 238170
rect -956 238046 -860 238102
rect -804 238046 -736 238102
rect -680 238046 -612 238102
rect -556 238046 -488 238102
rect -432 238046 -336 238102
rect -956 237978 -336 238046
rect -956 237922 -860 237978
rect -804 237922 -736 237978
rect -680 237922 -612 237978
rect -556 237922 -488 237978
rect -432 237922 -336 237978
rect -956 220350 -336 237922
rect -956 220294 -860 220350
rect -804 220294 -736 220350
rect -680 220294 -612 220350
rect -556 220294 -488 220350
rect -432 220294 -336 220350
rect -956 220226 -336 220294
rect -956 220170 -860 220226
rect -804 220170 -736 220226
rect -680 220170 -612 220226
rect -556 220170 -488 220226
rect -432 220170 -336 220226
rect -956 220102 -336 220170
rect -956 220046 -860 220102
rect -804 220046 -736 220102
rect -680 220046 -612 220102
rect -556 220046 -488 220102
rect -432 220046 -336 220102
rect -956 219978 -336 220046
rect -956 219922 -860 219978
rect -804 219922 -736 219978
rect -680 219922 -612 219978
rect -556 219922 -488 219978
rect -432 219922 -336 219978
rect -956 202350 -336 219922
rect -956 202294 -860 202350
rect -804 202294 -736 202350
rect -680 202294 -612 202350
rect -556 202294 -488 202350
rect -432 202294 -336 202350
rect -956 202226 -336 202294
rect -956 202170 -860 202226
rect -804 202170 -736 202226
rect -680 202170 -612 202226
rect -556 202170 -488 202226
rect -432 202170 -336 202226
rect -956 202102 -336 202170
rect -956 202046 -860 202102
rect -804 202046 -736 202102
rect -680 202046 -612 202102
rect -556 202046 -488 202102
rect -432 202046 -336 202102
rect -956 201978 -336 202046
rect -956 201922 -860 201978
rect -804 201922 -736 201978
rect -680 201922 -612 201978
rect -556 201922 -488 201978
rect -432 201922 -336 201978
rect -956 184350 -336 201922
rect -956 184294 -860 184350
rect -804 184294 -736 184350
rect -680 184294 -612 184350
rect -556 184294 -488 184350
rect -432 184294 -336 184350
rect -956 184226 -336 184294
rect -956 184170 -860 184226
rect -804 184170 -736 184226
rect -680 184170 -612 184226
rect -556 184170 -488 184226
rect -432 184170 -336 184226
rect -956 184102 -336 184170
rect -956 184046 -860 184102
rect -804 184046 -736 184102
rect -680 184046 -612 184102
rect -556 184046 -488 184102
rect -432 184046 -336 184102
rect -956 183978 -336 184046
rect -956 183922 -860 183978
rect -804 183922 -736 183978
rect -680 183922 -612 183978
rect -556 183922 -488 183978
rect -432 183922 -336 183978
rect -956 166350 -336 183922
rect -956 166294 -860 166350
rect -804 166294 -736 166350
rect -680 166294 -612 166350
rect -556 166294 -488 166350
rect -432 166294 -336 166350
rect -956 166226 -336 166294
rect -956 166170 -860 166226
rect -804 166170 -736 166226
rect -680 166170 -612 166226
rect -556 166170 -488 166226
rect -432 166170 -336 166226
rect -956 166102 -336 166170
rect -956 166046 -860 166102
rect -804 166046 -736 166102
rect -680 166046 -612 166102
rect -556 166046 -488 166102
rect -432 166046 -336 166102
rect -956 165978 -336 166046
rect -956 165922 -860 165978
rect -804 165922 -736 165978
rect -680 165922 -612 165978
rect -556 165922 -488 165978
rect -432 165922 -336 165978
rect -956 148350 -336 165922
rect -956 148294 -860 148350
rect -804 148294 -736 148350
rect -680 148294 -612 148350
rect -556 148294 -488 148350
rect -432 148294 -336 148350
rect -956 148226 -336 148294
rect -956 148170 -860 148226
rect -804 148170 -736 148226
rect -680 148170 -612 148226
rect -556 148170 -488 148226
rect -432 148170 -336 148226
rect -956 148102 -336 148170
rect -956 148046 -860 148102
rect -804 148046 -736 148102
rect -680 148046 -612 148102
rect -556 148046 -488 148102
rect -432 148046 -336 148102
rect -956 147978 -336 148046
rect -956 147922 -860 147978
rect -804 147922 -736 147978
rect -680 147922 -612 147978
rect -556 147922 -488 147978
rect -432 147922 -336 147978
rect -956 130350 -336 147922
rect -956 130294 -860 130350
rect -804 130294 -736 130350
rect -680 130294 -612 130350
rect -556 130294 -488 130350
rect -432 130294 -336 130350
rect -956 130226 -336 130294
rect -956 130170 -860 130226
rect -804 130170 -736 130226
rect -680 130170 -612 130226
rect -556 130170 -488 130226
rect -432 130170 -336 130226
rect -956 130102 -336 130170
rect -956 130046 -860 130102
rect -804 130046 -736 130102
rect -680 130046 -612 130102
rect -556 130046 -488 130102
rect -432 130046 -336 130102
rect -956 129978 -336 130046
rect -956 129922 -860 129978
rect -804 129922 -736 129978
rect -680 129922 -612 129978
rect -556 129922 -488 129978
rect -432 129922 -336 129978
rect -956 112350 -336 129922
rect -956 112294 -860 112350
rect -804 112294 -736 112350
rect -680 112294 -612 112350
rect -556 112294 -488 112350
rect -432 112294 -336 112350
rect -956 112226 -336 112294
rect -956 112170 -860 112226
rect -804 112170 -736 112226
rect -680 112170 -612 112226
rect -556 112170 -488 112226
rect -432 112170 -336 112226
rect -956 112102 -336 112170
rect -956 112046 -860 112102
rect -804 112046 -736 112102
rect -680 112046 -612 112102
rect -556 112046 -488 112102
rect -432 112046 -336 112102
rect -956 111978 -336 112046
rect -956 111922 -860 111978
rect -804 111922 -736 111978
rect -680 111922 -612 111978
rect -556 111922 -488 111978
rect -432 111922 -336 111978
rect -956 94350 -336 111922
rect -956 94294 -860 94350
rect -804 94294 -736 94350
rect -680 94294 -612 94350
rect -556 94294 -488 94350
rect -432 94294 -336 94350
rect -956 94226 -336 94294
rect -956 94170 -860 94226
rect -804 94170 -736 94226
rect -680 94170 -612 94226
rect -556 94170 -488 94226
rect -432 94170 -336 94226
rect -956 94102 -336 94170
rect -956 94046 -860 94102
rect -804 94046 -736 94102
rect -680 94046 -612 94102
rect -556 94046 -488 94102
rect -432 94046 -336 94102
rect -956 93978 -336 94046
rect -956 93922 -860 93978
rect -804 93922 -736 93978
rect -680 93922 -612 93978
rect -556 93922 -488 93978
rect -432 93922 -336 93978
rect -956 76350 -336 93922
rect -956 76294 -860 76350
rect -804 76294 -736 76350
rect -680 76294 -612 76350
rect -556 76294 -488 76350
rect -432 76294 -336 76350
rect -956 76226 -336 76294
rect -956 76170 -860 76226
rect -804 76170 -736 76226
rect -680 76170 -612 76226
rect -556 76170 -488 76226
rect -432 76170 -336 76226
rect -956 76102 -336 76170
rect -956 76046 -860 76102
rect -804 76046 -736 76102
rect -680 76046 -612 76102
rect -556 76046 -488 76102
rect -432 76046 -336 76102
rect -956 75978 -336 76046
rect -956 75922 -860 75978
rect -804 75922 -736 75978
rect -680 75922 -612 75978
rect -556 75922 -488 75978
rect -432 75922 -336 75978
rect -956 58350 -336 75922
rect -956 58294 -860 58350
rect -804 58294 -736 58350
rect -680 58294 -612 58350
rect -556 58294 -488 58350
rect -432 58294 -336 58350
rect -956 58226 -336 58294
rect -956 58170 -860 58226
rect -804 58170 -736 58226
rect -680 58170 -612 58226
rect -556 58170 -488 58226
rect -432 58170 -336 58226
rect -956 58102 -336 58170
rect -956 58046 -860 58102
rect -804 58046 -736 58102
rect -680 58046 -612 58102
rect -556 58046 -488 58102
rect -432 58046 -336 58102
rect -956 57978 -336 58046
rect -956 57922 -860 57978
rect -804 57922 -736 57978
rect -680 57922 -612 57978
rect -556 57922 -488 57978
rect -432 57922 -336 57978
rect -956 40350 -336 57922
rect -956 40294 -860 40350
rect -804 40294 -736 40350
rect -680 40294 -612 40350
rect -556 40294 -488 40350
rect -432 40294 -336 40350
rect -956 40226 -336 40294
rect -956 40170 -860 40226
rect -804 40170 -736 40226
rect -680 40170 -612 40226
rect -556 40170 -488 40226
rect -432 40170 -336 40226
rect -956 40102 -336 40170
rect -956 40046 -860 40102
rect -804 40046 -736 40102
rect -680 40046 -612 40102
rect -556 40046 -488 40102
rect -432 40046 -336 40102
rect -956 39978 -336 40046
rect -956 39922 -860 39978
rect -804 39922 -736 39978
rect -680 39922 -612 39978
rect -556 39922 -488 39978
rect -432 39922 -336 39978
rect -956 22350 -336 39922
rect -956 22294 -860 22350
rect -804 22294 -736 22350
rect -680 22294 -612 22350
rect -556 22294 -488 22350
rect -432 22294 -336 22350
rect -956 22226 -336 22294
rect -956 22170 -860 22226
rect -804 22170 -736 22226
rect -680 22170 -612 22226
rect -556 22170 -488 22226
rect -432 22170 -336 22226
rect -956 22102 -336 22170
rect -956 22046 -860 22102
rect -804 22046 -736 22102
rect -680 22046 -612 22102
rect -556 22046 -488 22102
rect -432 22046 -336 22102
rect -956 21978 -336 22046
rect -956 21922 -860 21978
rect -804 21922 -736 21978
rect -680 21922 -612 21978
rect -556 21922 -488 21978
rect -432 21922 -336 21978
rect -956 4350 -336 21922
rect -956 4294 -860 4350
rect -804 4294 -736 4350
rect -680 4294 -612 4350
rect -556 4294 -488 4350
rect -432 4294 -336 4350
rect -956 4226 -336 4294
rect -956 4170 -860 4226
rect -804 4170 -736 4226
rect -680 4170 -612 4226
rect -556 4170 -488 4226
rect -432 4170 -336 4226
rect -956 4102 -336 4170
rect -956 4046 -860 4102
rect -804 4046 -736 4102
rect -680 4046 -612 4102
rect -556 4046 -488 4102
rect -432 4046 -336 4102
rect -956 3978 -336 4046
rect -956 3922 -860 3978
rect -804 3922 -736 3978
rect -680 3922 -612 3978
rect -556 3922 -488 3978
rect -432 3922 -336 3978
rect -956 -160 -336 3922
rect -956 -216 -860 -160
rect -804 -216 -736 -160
rect -680 -216 -612 -160
rect -556 -216 -488 -160
rect -432 -216 -336 -160
rect -956 -284 -336 -216
rect -956 -340 -860 -284
rect -804 -340 -736 -284
rect -680 -340 -612 -284
rect -556 -340 -488 -284
rect -432 -340 -336 -284
rect -956 -408 -336 -340
rect -956 -464 -860 -408
rect -804 -464 -736 -408
rect -680 -464 -612 -408
rect -556 -464 -488 -408
rect -432 -464 -336 -408
rect -956 -532 -336 -464
rect -956 -588 -860 -532
rect -804 -588 -736 -532
rect -680 -588 -612 -532
rect -556 -588 -488 -532
rect -432 -588 -336 -532
rect -956 -684 -336 -588
rect 3154 597212 3774 598268
rect 3154 597156 3250 597212
rect 3306 597156 3374 597212
rect 3430 597156 3498 597212
rect 3554 597156 3622 597212
rect 3678 597156 3774 597212
rect 3154 597088 3774 597156
rect 3154 597032 3250 597088
rect 3306 597032 3374 597088
rect 3430 597032 3498 597088
rect 3554 597032 3622 597088
rect 3678 597032 3774 597088
rect 3154 596964 3774 597032
rect 3154 596908 3250 596964
rect 3306 596908 3374 596964
rect 3430 596908 3498 596964
rect 3554 596908 3622 596964
rect 3678 596908 3774 596964
rect 3154 596840 3774 596908
rect 3154 596784 3250 596840
rect 3306 596784 3374 596840
rect 3430 596784 3498 596840
rect 3554 596784 3622 596840
rect 3678 596784 3774 596840
rect 3154 580350 3774 596784
rect 3154 580294 3250 580350
rect 3306 580294 3374 580350
rect 3430 580294 3498 580350
rect 3554 580294 3622 580350
rect 3678 580294 3774 580350
rect 3154 580226 3774 580294
rect 3154 580170 3250 580226
rect 3306 580170 3374 580226
rect 3430 580170 3498 580226
rect 3554 580170 3622 580226
rect 3678 580170 3774 580226
rect 3154 580102 3774 580170
rect 3154 580046 3250 580102
rect 3306 580046 3374 580102
rect 3430 580046 3498 580102
rect 3554 580046 3622 580102
rect 3678 580046 3774 580102
rect 3154 579978 3774 580046
rect 3154 579922 3250 579978
rect 3306 579922 3374 579978
rect 3430 579922 3498 579978
rect 3554 579922 3622 579978
rect 3678 579922 3774 579978
rect 3154 562350 3774 579922
rect 3154 562294 3250 562350
rect 3306 562294 3374 562350
rect 3430 562294 3498 562350
rect 3554 562294 3622 562350
rect 3678 562294 3774 562350
rect 3154 562226 3774 562294
rect 3154 562170 3250 562226
rect 3306 562170 3374 562226
rect 3430 562170 3498 562226
rect 3554 562170 3622 562226
rect 3678 562170 3774 562226
rect 3154 562102 3774 562170
rect 3154 562046 3250 562102
rect 3306 562046 3374 562102
rect 3430 562046 3498 562102
rect 3554 562046 3622 562102
rect 3678 562046 3774 562102
rect 3154 561978 3774 562046
rect 3154 561922 3250 561978
rect 3306 561922 3374 561978
rect 3430 561922 3498 561978
rect 3554 561922 3622 561978
rect 3678 561922 3774 561978
rect 3154 544350 3774 561922
rect 6874 598172 7494 598268
rect 6874 598116 6970 598172
rect 7026 598116 7094 598172
rect 7150 598116 7218 598172
rect 7274 598116 7342 598172
rect 7398 598116 7494 598172
rect 6874 598048 7494 598116
rect 6874 597992 6970 598048
rect 7026 597992 7094 598048
rect 7150 597992 7218 598048
rect 7274 597992 7342 598048
rect 7398 597992 7494 598048
rect 6874 597924 7494 597992
rect 6874 597868 6970 597924
rect 7026 597868 7094 597924
rect 7150 597868 7218 597924
rect 7274 597868 7342 597924
rect 7398 597868 7494 597924
rect 6874 597800 7494 597868
rect 6874 597744 6970 597800
rect 7026 597744 7094 597800
rect 7150 597744 7218 597800
rect 7274 597744 7342 597800
rect 7398 597744 7494 597800
rect 6874 586350 7494 597744
rect 6874 586294 6970 586350
rect 7026 586294 7094 586350
rect 7150 586294 7218 586350
rect 7274 586294 7342 586350
rect 7398 586294 7494 586350
rect 6874 586226 7494 586294
rect 6874 586170 6970 586226
rect 7026 586170 7094 586226
rect 7150 586170 7218 586226
rect 7274 586170 7342 586226
rect 7398 586170 7494 586226
rect 6874 586102 7494 586170
rect 6874 586046 6970 586102
rect 7026 586046 7094 586102
rect 7150 586046 7218 586102
rect 7274 586046 7342 586102
rect 7398 586046 7494 586102
rect 6874 585978 7494 586046
rect 6874 585922 6970 585978
rect 7026 585922 7094 585978
rect 7150 585922 7218 585978
rect 7274 585922 7342 585978
rect 7398 585922 7494 585978
rect 6874 568350 7494 585922
rect 6874 568294 6970 568350
rect 7026 568294 7094 568350
rect 7150 568294 7218 568350
rect 7274 568294 7342 568350
rect 7398 568294 7494 568350
rect 6874 568226 7494 568294
rect 6874 568170 6970 568226
rect 7026 568170 7094 568226
rect 7150 568170 7218 568226
rect 7274 568170 7342 568226
rect 7398 568170 7494 568226
rect 6874 568102 7494 568170
rect 6874 568046 6970 568102
rect 7026 568046 7094 568102
rect 7150 568046 7218 568102
rect 7274 568046 7342 568102
rect 7398 568046 7494 568102
rect 6874 567978 7494 568046
rect 6874 567922 6970 567978
rect 7026 567922 7094 567978
rect 7150 567922 7218 567978
rect 7274 567922 7342 567978
rect 7398 567922 7494 567978
rect 6874 550350 7494 567922
rect 6874 550294 6970 550350
rect 7026 550294 7094 550350
rect 7150 550294 7218 550350
rect 7274 550294 7342 550350
rect 7398 550294 7494 550350
rect 6874 550226 7494 550294
rect 6874 550170 6970 550226
rect 7026 550170 7094 550226
rect 7150 550170 7218 550226
rect 7274 550170 7342 550226
rect 7398 550170 7494 550226
rect 6874 550102 7494 550170
rect 6874 550046 6970 550102
rect 7026 550046 7094 550102
rect 7150 550046 7218 550102
rect 7274 550046 7342 550102
rect 7398 550046 7494 550102
rect 6874 549978 7494 550046
rect 6874 549922 6970 549978
rect 7026 549922 7094 549978
rect 7150 549922 7218 549978
rect 7274 549922 7342 549978
rect 7398 549922 7494 549978
rect 3154 544294 3250 544350
rect 3306 544294 3374 544350
rect 3430 544294 3498 544350
rect 3554 544294 3622 544350
rect 3678 544294 3774 544350
rect 3154 544226 3774 544294
rect 3154 544170 3250 544226
rect 3306 544170 3374 544226
rect 3430 544170 3498 544226
rect 3554 544170 3622 544226
rect 3678 544170 3774 544226
rect 3154 544102 3774 544170
rect 3154 544046 3250 544102
rect 3306 544046 3374 544102
rect 3430 544046 3498 544102
rect 3554 544046 3622 544102
rect 3678 544046 3774 544102
rect 3154 543978 3774 544046
rect 3154 543922 3250 543978
rect 3306 543922 3374 543978
rect 3430 543922 3498 543978
rect 3554 543922 3622 543978
rect 3678 543922 3774 543978
rect 3154 526350 3774 543922
rect 3154 526294 3250 526350
rect 3306 526294 3374 526350
rect 3430 526294 3498 526350
rect 3554 526294 3622 526350
rect 3678 526294 3774 526350
rect 3154 526226 3774 526294
rect 3154 526170 3250 526226
rect 3306 526170 3374 526226
rect 3430 526170 3498 526226
rect 3554 526170 3622 526226
rect 3678 526170 3774 526226
rect 3154 526102 3774 526170
rect 3154 526046 3250 526102
rect 3306 526046 3374 526102
rect 3430 526046 3498 526102
rect 3554 526046 3622 526102
rect 3678 526046 3774 526102
rect 3154 525978 3774 526046
rect 3154 525922 3250 525978
rect 3306 525922 3374 525978
rect 3430 525922 3498 525978
rect 3554 525922 3622 525978
rect 3678 525922 3774 525978
rect 3154 508350 3774 525922
rect 3154 508294 3250 508350
rect 3306 508294 3374 508350
rect 3430 508294 3498 508350
rect 3554 508294 3622 508350
rect 3678 508294 3774 508350
rect 3154 508226 3774 508294
rect 3154 508170 3250 508226
rect 3306 508170 3374 508226
rect 3430 508170 3498 508226
rect 3554 508170 3622 508226
rect 3678 508170 3774 508226
rect 3154 508102 3774 508170
rect 3154 508046 3250 508102
rect 3306 508046 3374 508102
rect 3430 508046 3498 508102
rect 3554 508046 3622 508102
rect 3678 508046 3774 508102
rect 3154 507978 3774 508046
rect 3154 507922 3250 507978
rect 3306 507922 3374 507978
rect 3430 507922 3498 507978
rect 3554 507922 3622 507978
rect 3678 507922 3774 507978
rect 3154 490350 3774 507922
rect 3154 490294 3250 490350
rect 3306 490294 3374 490350
rect 3430 490294 3498 490350
rect 3554 490294 3622 490350
rect 3678 490294 3774 490350
rect 3154 490226 3774 490294
rect 3154 490170 3250 490226
rect 3306 490170 3374 490226
rect 3430 490170 3498 490226
rect 3554 490170 3622 490226
rect 3678 490170 3774 490226
rect 3154 490102 3774 490170
rect 3154 490046 3250 490102
rect 3306 490046 3374 490102
rect 3430 490046 3498 490102
rect 3554 490046 3622 490102
rect 3678 490046 3774 490102
rect 3154 489978 3774 490046
rect 3154 489922 3250 489978
rect 3306 489922 3374 489978
rect 3430 489922 3498 489978
rect 3554 489922 3622 489978
rect 3678 489922 3774 489978
rect 3154 472350 3774 489922
rect 5852 544852 5908 544862
rect 3154 472294 3250 472350
rect 3306 472294 3374 472350
rect 3430 472294 3498 472350
rect 3554 472294 3622 472350
rect 3678 472294 3774 472350
rect 3154 472226 3774 472294
rect 3154 472170 3250 472226
rect 3306 472170 3374 472226
rect 3430 472170 3498 472226
rect 3554 472170 3622 472226
rect 3678 472170 3774 472226
rect 3154 472102 3774 472170
rect 3154 472046 3250 472102
rect 3306 472046 3374 472102
rect 3430 472046 3498 472102
rect 3554 472046 3622 472102
rect 3678 472046 3774 472102
rect 3154 471978 3774 472046
rect 3154 471922 3250 471978
rect 3306 471922 3374 471978
rect 3430 471922 3498 471978
rect 3554 471922 3622 471978
rect 3678 471922 3774 471978
rect 3154 454350 3774 471922
rect 3154 454294 3250 454350
rect 3306 454294 3374 454350
rect 3430 454294 3498 454350
rect 3554 454294 3622 454350
rect 3678 454294 3774 454350
rect 3154 454226 3774 454294
rect 3154 454170 3250 454226
rect 3306 454170 3374 454226
rect 3430 454170 3498 454226
rect 3554 454170 3622 454226
rect 3678 454170 3774 454226
rect 3154 454102 3774 454170
rect 3154 454046 3250 454102
rect 3306 454046 3374 454102
rect 3430 454046 3498 454102
rect 3554 454046 3622 454102
rect 3678 454046 3774 454102
rect 3154 453978 3774 454046
rect 3154 453922 3250 453978
rect 3306 453922 3374 453978
rect 3430 453922 3498 453978
rect 3554 453922 3622 453978
rect 3678 453922 3774 453978
rect 3154 436350 3774 453922
rect 3154 436294 3250 436350
rect 3306 436294 3374 436350
rect 3430 436294 3498 436350
rect 3554 436294 3622 436350
rect 3678 436294 3774 436350
rect 3154 436226 3774 436294
rect 3154 436170 3250 436226
rect 3306 436170 3374 436226
rect 3430 436170 3498 436226
rect 3554 436170 3622 436226
rect 3678 436170 3774 436226
rect 3154 436102 3774 436170
rect 3154 436046 3250 436102
rect 3306 436046 3374 436102
rect 3430 436046 3498 436102
rect 3554 436046 3622 436102
rect 3678 436046 3774 436102
rect 3154 435978 3774 436046
rect 3154 435922 3250 435978
rect 3306 435922 3374 435978
rect 3430 435922 3498 435978
rect 3554 435922 3622 435978
rect 3678 435922 3774 435978
rect 3154 418350 3774 435922
rect 3154 418294 3250 418350
rect 3306 418294 3374 418350
rect 3430 418294 3498 418350
rect 3554 418294 3622 418350
rect 3678 418294 3774 418350
rect 3154 418226 3774 418294
rect 3154 418170 3250 418226
rect 3306 418170 3374 418226
rect 3430 418170 3498 418226
rect 3554 418170 3622 418226
rect 3678 418170 3774 418226
rect 3154 418102 3774 418170
rect 3154 418046 3250 418102
rect 3306 418046 3374 418102
rect 3430 418046 3498 418102
rect 3554 418046 3622 418102
rect 3678 418046 3774 418102
rect 3154 417978 3774 418046
rect 3154 417922 3250 417978
rect 3306 417922 3374 417978
rect 3430 417922 3498 417978
rect 3554 417922 3622 417978
rect 3678 417922 3774 417978
rect 3154 400350 3774 417922
rect 3154 400294 3250 400350
rect 3306 400294 3374 400350
rect 3430 400294 3498 400350
rect 3554 400294 3622 400350
rect 3678 400294 3774 400350
rect 3154 400226 3774 400294
rect 3154 400170 3250 400226
rect 3306 400170 3374 400226
rect 3430 400170 3498 400226
rect 3554 400170 3622 400226
rect 3678 400170 3774 400226
rect 3154 400102 3774 400170
rect 3154 400046 3250 400102
rect 3306 400046 3374 400102
rect 3430 400046 3498 400102
rect 3554 400046 3622 400102
rect 3678 400046 3774 400102
rect 3154 399978 3774 400046
rect 3154 399922 3250 399978
rect 3306 399922 3374 399978
rect 3430 399922 3498 399978
rect 3554 399922 3622 399978
rect 3678 399922 3774 399978
rect 3154 382350 3774 399922
rect 3154 382294 3250 382350
rect 3306 382294 3374 382350
rect 3430 382294 3498 382350
rect 3554 382294 3622 382350
rect 3678 382294 3774 382350
rect 3154 382226 3774 382294
rect 3154 382170 3250 382226
rect 3306 382170 3374 382226
rect 3430 382170 3498 382226
rect 3554 382170 3622 382226
rect 3678 382170 3774 382226
rect 3154 382102 3774 382170
rect 3154 382046 3250 382102
rect 3306 382046 3374 382102
rect 3430 382046 3498 382102
rect 3554 382046 3622 382102
rect 3678 382046 3774 382102
rect 3154 381978 3774 382046
rect 3154 381922 3250 381978
rect 3306 381922 3374 381978
rect 3430 381922 3498 381978
rect 3554 381922 3622 381978
rect 3678 381922 3774 381978
rect 3154 364350 3774 381922
rect 3154 364294 3250 364350
rect 3306 364294 3374 364350
rect 3430 364294 3498 364350
rect 3554 364294 3622 364350
rect 3678 364294 3774 364350
rect 3154 364226 3774 364294
rect 3154 364170 3250 364226
rect 3306 364170 3374 364226
rect 3430 364170 3498 364226
rect 3554 364170 3622 364226
rect 3678 364170 3774 364226
rect 3154 364102 3774 364170
rect 3154 364046 3250 364102
rect 3306 364046 3374 364102
rect 3430 364046 3498 364102
rect 3554 364046 3622 364102
rect 3678 364046 3774 364102
rect 3154 363978 3774 364046
rect 3154 363922 3250 363978
rect 3306 363922 3374 363978
rect 3430 363922 3498 363978
rect 3554 363922 3622 363978
rect 3678 363922 3774 363978
rect 3154 346350 3774 363922
rect 3154 346294 3250 346350
rect 3306 346294 3374 346350
rect 3430 346294 3498 346350
rect 3554 346294 3622 346350
rect 3678 346294 3774 346350
rect 3154 346226 3774 346294
rect 3154 346170 3250 346226
rect 3306 346170 3374 346226
rect 3430 346170 3498 346226
rect 3554 346170 3622 346226
rect 3678 346170 3774 346226
rect 3154 346102 3774 346170
rect 3154 346046 3250 346102
rect 3306 346046 3374 346102
rect 3430 346046 3498 346102
rect 3554 346046 3622 346102
rect 3678 346046 3774 346102
rect 3154 345978 3774 346046
rect 3154 345922 3250 345978
rect 3306 345922 3374 345978
rect 3430 345922 3498 345978
rect 3554 345922 3622 345978
rect 3678 345922 3774 345978
rect 3154 328350 3774 345922
rect 3154 328294 3250 328350
rect 3306 328294 3374 328350
rect 3430 328294 3498 328350
rect 3554 328294 3622 328350
rect 3678 328294 3774 328350
rect 3154 328226 3774 328294
rect 3154 328170 3250 328226
rect 3306 328170 3374 328226
rect 3430 328170 3498 328226
rect 3554 328170 3622 328226
rect 3678 328170 3774 328226
rect 3154 328102 3774 328170
rect 3154 328046 3250 328102
rect 3306 328046 3374 328102
rect 3430 328046 3498 328102
rect 3554 328046 3622 328102
rect 3678 328046 3774 328102
rect 3154 327978 3774 328046
rect 3154 327922 3250 327978
rect 3306 327922 3374 327978
rect 3430 327922 3498 327978
rect 3554 327922 3622 327978
rect 3678 327922 3774 327978
rect 3154 310350 3774 327922
rect 3154 310294 3250 310350
rect 3306 310294 3374 310350
rect 3430 310294 3498 310350
rect 3554 310294 3622 310350
rect 3678 310294 3774 310350
rect 3154 310226 3774 310294
rect 3154 310170 3250 310226
rect 3306 310170 3374 310226
rect 3430 310170 3498 310226
rect 3554 310170 3622 310226
rect 3678 310170 3774 310226
rect 3154 310102 3774 310170
rect 3154 310046 3250 310102
rect 3306 310046 3374 310102
rect 3430 310046 3498 310102
rect 3554 310046 3622 310102
rect 3678 310046 3774 310102
rect 3154 309978 3774 310046
rect 3154 309922 3250 309978
rect 3306 309922 3374 309978
rect 3430 309922 3498 309978
rect 3554 309922 3622 309978
rect 3678 309922 3774 309978
rect 3154 292350 3774 309922
rect 3154 292294 3250 292350
rect 3306 292294 3374 292350
rect 3430 292294 3498 292350
rect 3554 292294 3622 292350
rect 3678 292294 3774 292350
rect 3154 292226 3774 292294
rect 3154 292170 3250 292226
rect 3306 292170 3374 292226
rect 3430 292170 3498 292226
rect 3554 292170 3622 292226
rect 3678 292170 3774 292226
rect 3154 292102 3774 292170
rect 3154 292046 3250 292102
rect 3306 292046 3374 292102
rect 3430 292046 3498 292102
rect 3554 292046 3622 292102
rect 3678 292046 3774 292102
rect 3154 291978 3774 292046
rect 3154 291922 3250 291978
rect 3306 291922 3374 291978
rect 3430 291922 3498 291978
rect 3554 291922 3622 291978
rect 3678 291922 3774 291978
rect 3154 274350 3774 291922
rect 3154 274294 3250 274350
rect 3306 274294 3374 274350
rect 3430 274294 3498 274350
rect 3554 274294 3622 274350
rect 3678 274294 3774 274350
rect 3154 274226 3774 274294
rect 3154 274170 3250 274226
rect 3306 274170 3374 274226
rect 3430 274170 3498 274226
rect 3554 274170 3622 274226
rect 3678 274170 3774 274226
rect 3154 274102 3774 274170
rect 3154 274046 3250 274102
rect 3306 274046 3374 274102
rect 3430 274046 3498 274102
rect 3554 274046 3622 274102
rect 3678 274046 3774 274102
rect 3154 273978 3774 274046
rect 3154 273922 3250 273978
rect 3306 273922 3374 273978
rect 3430 273922 3498 273978
rect 3554 273922 3622 273978
rect 3678 273922 3774 273978
rect 3154 256350 3774 273922
rect 3154 256294 3250 256350
rect 3306 256294 3374 256350
rect 3430 256294 3498 256350
rect 3554 256294 3622 256350
rect 3678 256294 3774 256350
rect 3154 256226 3774 256294
rect 3154 256170 3250 256226
rect 3306 256170 3374 256226
rect 3430 256170 3498 256226
rect 3554 256170 3622 256226
rect 3678 256170 3774 256226
rect 3154 256102 3774 256170
rect 3154 256046 3250 256102
rect 3306 256046 3374 256102
rect 3430 256046 3498 256102
rect 3554 256046 3622 256102
rect 3678 256046 3774 256102
rect 3154 255978 3774 256046
rect 3154 255922 3250 255978
rect 3306 255922 3374 255978
rect 3430 255922 3498 255978
rect 3554 255922 3622 255978
rect 3678 255922 3774 255978
rect 3154 238350 3774 255922
rect 3154 238294 3250 238350
rect 3306 238294 3374 238350
rect 3430 238294 3498 238350
rect 3554 238294 3622 238350
rect 3678 238294 3774 238350
rect 3154 238226 3774 238294
rect 3154 238170 3250 238226
rect 3306 238170 3374 238226
rect 3430 238170 3498 238226
rect 3554 238170 3622 238226
rect 3678 238170 3774 238226
rect 3154 238102 3774 238170
rect 3154 238046 3250 238102
rect 3306 238046 3374 238102
rect 3430 238046 3498 238102
rect 3554 238046 3622 238102
rect 3678 238046 3774 238102
rect 3154 237978 3774 238046
rect 3154 237922 3250 237978
rect 3306 237922 3374 237978
rect 3430 237922 3498 237978
rect 3554 237922 3622 237978
rect 3678 237922 3774 237978
rect 3154 220350 3774 237922
rect 3154 220294 3250 220350
rect 3306 220294 3374 220350
rect 3430 220294 3498 220350
rect 3554 220294 3622 220350
rect 3678 220294 3774 220350
rect 3154 220226 3774 220294
rect 3154 220170 3250 220226
rect 3306 220170 3374 220226
rect 3430 220170 3498 220226
rect 3554 220170 3622 220226
rect 3678 220170 3774 220226
rect 3154 220102 3774 220170
rect 3154 220046 3250 220102
rect 3306 220046 3374 220102
rect 3430 220046 3498 220102
rect 3554 220046 3622 220102
rect 3678 220046 3774 220102
rect 3154 219978 3774 220046
rect 3154 219922 3250 219978
rect 3306 219922 3374 219978
rect 3430 219922 3498 219978
rect 3554 219922 3622 219978
rect 3678 219922 3774 219978
rect 3154 202350 3774 219922
rect 3154 202294 3250 202350
rect 3306 202294 3374 202350
rect 3430 202294 3498 202350
rect 3554 202294 3622 202350
rect 3678 202294 3774 202350
rect 3154 202226 3774 202294
rect 3154 202170 3250 202226
rect 3306 202170 3374 202226
rect 3430 202170 3498 202226
rect 3554 202170 3622 202226
rect 3678 202170 3774 202226
rect 3154 202102 3774 202170
rect 3154 202046 3250 202102
rect 3306 202046 3374 202102
rect 3430 202046 3498 202102
rect 3554 202046 3622 202102
rect 3678 202046 3774 202102
rect 3154 201978 3774 202046
rect 3154 201922 3250 201978
rect 3306 201922 3374 201978
rect 3430 201922 3498 201978
rect 3554 201922 3622 201978
rect 3678 201922 3774 201978
rect 3154 184350 3774 201922
rect 3154 184294 3250 184350
rect 3306 184294 3374 184350
rect 3430 184294 3498 184350
rect 3554 184294 3622 184350
rect 3678 184294 3774 184350
rect 3154 184226 3774 184294
rect 3154 184170 3250 184226
rect 3306 184170 3374 184226
rect 3430 184170 3498 184226
rect 3554 184170 3622 184226
rect 3678 184170 3774 184226
rect 3154 184102 3774 184170
rect 3154 184046 3250 184102
rect 3306 184046 3374 184102
rect 3430 184046 3498 184102
rect 3554 184046 3622 184102
rect 3678 184046 3774 184102
rect 3154 183978 3774 184046
rect 3154 183922 3250 183978
rect 3306 183922 3374 183978
rect 3430 183922 3498 183978
rect 3554 183922 3622 183978
rect 3678 183922 3774 183978
rect 3154 166350 3774 183922
rect 3154 166294 3250 166350
rect 3306 166294 3374 166350
rect 3430 166294 3498 166350
rect 3554 166294 3622 166350
rect 3678 166294 3774 166350
rect 3154 166226 3774 166294
rect 3154 166170 3250 166226
rect 3306 166170 3374 166226
rect 3430 166170 3498 166226
rect 3554 166170 3622 166226
rect 3678 166170 3774 166226
rect 3154 166102 3774 166170
rect 3154 166046 3250 166102
rect 3306 166046 3374 166102
rect 3430 166046 3498 166102
rect 3554 166046 3622 166102
rect 3678 166046 3774 166102
rect 3154 165978 3774 166046
rect 3154 165922 3250 165978
rect 3306 165922 3374 165978
rect 3430 165922 3498 165978
rect 3554 165922 3622 165978
rect 3678 165922 3774 165978
rect 3154 148350 3774 165922
rect 4172 488404 4228 488414
rect 4172 164276 4228 488348
rect 4172 164210 4228 164220
rect 4284 403732 4340 403742
rect 3154 148294 3250 148350
rect 3306 148294 3374 148350
rect 3430 148294 3498 148350
rect 3554 148294 3622 148350
rect 3678 148294 3774 148350
rect 3154 148226 3774 148294
rect 3154 148170 3250 148226
rect 3306 148170 3374 148226
rect 3430 148170 3498 148226
rect 3554 148170 3622 148226
rect 3678 148170 3774 148226
rect 3154 148102 3774 148170
rect 3154 148046 3250 148102
rect 3306 148046 3374 148102
rect 3430 148046 3498 148102
rect 3554 148046 3622 148102
rect 3678 148046 3774 148102
rect 3154 147978 3774 148046
rect 3154 147922 3250 147978
rect 3306 147922 3374 147978
rect 3430 147922 3498 147978
rect 3554 147922 3622 147978
rect 3678 147922 3774 147978
rect 3154 130350 3774 147922
rect 4284 141428 4340 403676
rect 4284 141362 4340 141372
rect 4396 220276 4452 220286
rect 3154 130294 3250 130350
rect 3306 130294 3374 130350
rect 3430 130294 3498 130350
rect 3554 130294 3622 130350
rect 3678 130294 3774 130350
rect 3154 130226 3774 130294
rect 3154 130170 3250 130226
rect 3306 130170 3374 130226
rect 3430 130170 3498 130226
rect 3554 130170 3622 130226
rect 3678 130170 3774 130226
rect 3154 130102 3774 130170
rect 3154 130046 3250 130102
rect 3306 130046 3374 130102
rect 3430 130046 3498 130102
rect 3554 130046 3622 130102
rect 3678 130046 3774 130102
rect 3154 129978 3774 130046
rect 3154 129922 3250 129978
rect 3306 129922 3374 129978
rect 3430 129922 3498 129978
rect 3554 129922 3622 129978
rect 3678 129922 3774 129978
rect 3154 112350 3774 129922
rect 3154 112294 3250 112350
rect 3306 112294 3374 112350
rect 3430 112294 3498 112350
rect 3554 112294 3622 112350
rect 3678 112294 3774 112350
rect 3154 112226 3774 112294
rect 3154 112170 3250 112226
rect 3306 112170 3374 112226
rect 3430 112170 3498 112226
rect 3554 112170 3622 112226
rect 3678 112170 3774 112226
rect 3154 112102 3774 112170
rect 3154 112046 3250 112102
rect 3306 112046 3374 112102
rect 3430 112046 3498 112102
rect 3554 112046 3622 112102
rect 3678 112046 3774 112102
rect 3154 111978 3774 112046
rect 3154 111922 3250 111978
rect 3306 111922 3374 111978
rect 3430 111922 3498 111978
rect 3554 111922 3622 111978
rect 3678 111922 3774 111978
rect 3154 94350 3774 111922
rect 3154 94294 3250 94350
rect 3306 94294 3374 94350
rect 3430 94294 3498 94350
rect 3554 94294 3622 94350
rect 3678 94294 3774 94350
rect 3154 94226 3774 94294
rect 3154 94170 3250 94226
rect 3306 94170 3374 94226
rect 3430 94170 3498 94226
rect 3554 94170 3622 94226
rect 3678 94170 3774 94226
rect 3154 94102 3774 94170
rect 3154 94046 3250 94102
rect 3306 94046 3374 94102
rect 3430 94046 3498 94102
rect 3554 94046 3622 94102
rect 3678 94046 3774 94102
rect 3154 93978 3774 94046
rect 3154 93922 3250 93978
rect 3306 93922 3374 93978
rect 3430 93922 3498 93978
rect 3554 93922 3622 93978
rect 3678 93922 3774 93978
rect 3154 76350 3774 93922
rect 3154 76294 3250 76350
rect 3306 76294 3374 76350
rect 3430 76294 3498 76350
rect 3554 76294 3622 76350
rect 3678 76294 3774 76350
rect 3154 76226 3774 76294
rect 3154 76170 3250 76226
rect 3306 76170 3374 76226
rect 3430 76170 3498 76226
rect 3554 76170 3622 76226
rect 3678 76170 3774 76226
rect 3154 76102 3774 76170
rect 3154 76046 3250 76102
rect 3306 76046 3374 76102
rect 3430 76046 3498 76102
rect 3554 76046 3622 76102
rect 3678 76046 3774 76102
rect 3154 75978 3774 76046
rect 3154 75922 3250 75978
rect 3306 75922 3374 75978
rect 3430 75922 3498 75978
rect 3554 75922 3622 75978
rect 3678 75922 3774 75978
rect 3154 58350 3774 75922
rect 4172 135604 4228 135614
rect 4172 69076 4228 135548
rect 4172 69010 4228 69020
rect 4284 107380 4340 107390
rect 3154 58294 3250 58350
rect 3306 58294 3374 58350
rect 3430 58294 3498 58350
rect 3554 58294 3622 58350
rect 3678 58294 3774 58350
rect 3154 58226 3774 58294
rect 3154 58170 3250 58226
rect 3306 58170 3374 58226
rect 3430 58170 3498 58226
rect 3554 58170 3622 58226
rect 3678 58170 3774 58226
rect 3154 58102 3774 58170
rect 3154 58046 3250 58102
rect 3306 58046 3374 58102
rect 3430 58046 3498 58102
rect 3554 58046 3622 58102
rect 3678 58046 3774 58102
rect 3154 57978 3774 58046
rect 3154 57922 3250 57978
rect 3306 57922 3374 57978
rect 3430 57922 3498 57978
rect 3554 57922 3622 57978
rect 3678 57922 3774 57978
rect 3154 40350 3774 57922
rect 4172 65044 4228 65054
rect 4172 50036 4228 64988
rect 4284 61460 4340 107324
rect 4396 91924 4452 220220
rect 5852 179508 5908 544796
rect 6874 532350 7494 549922
rect 6874 532294 6970 532350
rect 7026 532294 7094 532350
rect 7150 532294 7218 532350
rect 7274 532294 7342 532350
rect 7398 532294 7494 532350
rect 6874 532226 7494 532294
rect 6874 532170 6970 532226
rect 7026 532170 7094 532226
rect 7150 532170 7218 532226
rect 7274 532170 7342 532226
rect 7398 532170 7494 532226
rect 6874 532102 7494 532170
rect 6874 532046 6970 532102
rect 7026 532046 7094 532102
rect 7150 532046 7218 532102
rect 7274 532046 7342 532102
rect 7398 532046 7494 532102
rect 6874 531978 7494 532046
rect 6874 531922 6970 531978
rect 7026 531922 7094 531978
rect 7150 531922 7218 531978
rect 7274 531922 7342 531978
rect 7398 531922 7494 531978
rect 6874 514350 7494 531922
rect 6874 514294 6970 514350
rect 7026 514294 7094 514350
rect 7150 514294 7218 514350
rect 7274 514294 7342 514350
rect 7398 514294 7494 514350
rect 6874 514226 7494 514294
rect 6874 514170 6970 514226
rect 7026 514170 7094 514226
rect 7150 514170 7218 514226
rect 7274 514170 7342 514226
rect 7398 514170 7494 514226
rect 6874 514102 7494 514170
rect 6874 514046 6970 514102
rect 7026 514046 7094 514102
rect 7150 514046 7218 514102
rect 7274 514046 7342 514102
rect 7398 514046 7494 514102
rect 6874 513978 7494 514046
rect 6874 513922 6970 513978
rect 7026 513922 7094 513978
rect 7150 513922 7218 513978
rect 7274 513922 7342 513978
rect 7398 513922 7494 513978
rect 6874 496350 7494 513922
rect 21154 597212 21774 598268
rect 21154 597156 21250 597212
rect 21306 597156 21374 597212
rect 21430 597156 21498 597212
rect 21554 597156 21622 597212
rect 21678 597156 21774 597212
rect 21154 597088 21774 597156
rect 21154 597032 21250 597088
rect 21306 597032 21374 597088
rect 21430 597032 21498 597088
rect 21554 597032 21622 597088
rect 21678 597032 21774 597088
rect 21154 596964 21774 597032
rect 21154 596908 21250 596964
rect 21306 596908 21374 596964
rect 21430 596908 21498 596964
rect 21554 596908 21622 596964
rect 21678 596908 21774 596964
rect 21154 596840 21774 596908
rect 21154 596784 21250 596840
rect 21306 596784 21374 596840
rect 21430 596784 21498 596840
rect 21554 596784 21622 596840
rect 21678 596784 21774 596840
rect 21154 580350 21774 596784
rect 21154 580294 21250 580350
rect 21306 580294 21374 580350
rect 21430 580294 21498 580350
rect 21554 580294 21622 580350
rect 21678 580294 21774 580350
rect 21154 580226 21774 580294
rect 21154 580170 21250 580226
rect 21306 580170 21374 580226
rect 21430 580170 21498 580226
rect 21554 580170 21622 580226
rect 21678 580170 21774 580226
rect 21154 580102 21774 580170
rect 21154 580046 21250 580102
rect 21306 580046 21374 580102
rect 21430 580046 21498 580102
rect 21554 580046 21622 580102
rect 21678 580046 21774 580102
rect 21154 579978 21774 580046
rect 21154 579922 21250 579978
rect 21306 579922 21374 579978
rect 21430 579922 21498 579978
rect 21554 579922 21622 579978
rect 21678 579922 21774 579978
rect 21154 562350 21774 579922
rect 21154 562294 21250 562350
rect 21306 562294 21374 562350
rect 21430 562294 21498 562350
rect 21554 562294 21622 562350
rect 21678 562294 21774 562350
rect 21154 562226 21774 562294
rect 21154 562170 21250 562226
rect 21306 562170 21374 562226
rect 21430 562170 21498 562226
rect 21554 562170 21622 562226
rect 21678 562170 21774 562226
rect 21154 562102 21774 562170
rect 21154 562046 21250 562102
rect 21306 562046 21374 562102
rect 21430 562046 21498 562102
rect 21554 562046 21622 562102
rect 21678 562046 21774 562102
rect 21154 561978 21774 562046
rect 21154 561922 21250 561978
rect 21306 561922 21374 561978
rect 21430 561922 21498 561978
rect 21554 561922 21622 561978
rect 21678 561922 21774 561978
rect 21154 544350 21774 561922
rect 21154 544294 21250 544350
rect 21306 544294 21374 544350
rect 21430 544294 21498 544350
rect 21554 544294 21622 544350
rect 21678 544294 21774 544350
rect 21154 544226 21774 544294
rect 21154 544170 21250 544226
rect 21306 544170 21374 544226
rect 21430 544170 21498 544226
rect 21554 544170 21622 544226
rect 21678 544170 21774 544226
rect 21154 544102 21774 544170
rect 21154 544046 21250 544102
rect 21306 544046 21374 544102
rect 21430 544046 21498 544102
rect 21554 544046 21622 544102
rect 21678 544046 21774 544102
rect 21154 543978 21774 544046
rect 21154 543922 21250 543978
rect 21306 543922 21374 543978
rect 21430 543922 21498 543978
rect 21554 543922 21622 543978
rect 21678 543922 21774 543978
rect 21154 526350 21774 543922
rect 24874 598172 25494 598268
rect 24874 598116 24970 598172
rect 25026 598116 25094 598172
rect 25150 598116 25218 598172
rect 25274 598116 25342 598172
rect 25398 598116 25494 598172
rect 24874 598048 25494 598116
rect 24874 597992 24970 598048
rect 25026 597992 25094 598048
rect 25150 597992 25218 598048
rect 25274 597992 25342 598048
rect 25398 597992 25494 598048
rect 24874 597924 25494 597992
rect 24874 597868 24970 597924
rect 25026 597868 25094 597924
rect 25150 597868 25218 597924
rect 25274 597868 25342 597924
rect 25398 597868 25494 597924
rect 24874 597800 25494 597868
rect 24874 597744 24970 597800
rect 25026 597744 25094 597800
rect 25150 597744 25218 597800
rect 25274 597744 25342 597800
rect 25398 597744 25494 597800
rect 24874 586350 25494 597744
rect 39154 597212 39774 598268
rect 39154 597156 39250 597212
rect 39306 597156 39374 597212
rect 39430 597156 39498 597212
rect 39554 597156 39622 597212
rect 39678 597156 39774 597212
rect 39154 597088 39774 597156
rect 39154 597032 39250 597088
rect 39306 597032 39374 597088
rect 39430 597032 39498 597088
rect 39554 597032 39622 597088
rect 39678 597032 39774 597088
rect 39154 596964 39774 597032
rect 39154 596908 39250 596964
rect 39306 596908 39374 596964
rect 39430 596908 39498 596964
rect 39554 596908 39622 596964
rect 39678 596908 39774 596964
rect 39154 596840 39774 596908
rect 39154 596784 39250 596840
rect 39306 596784 39374 596840
rect 39430 596784 39498 596840
rect 39554 596784 39622 596840
rect 39678 596784 39774 596840
rect 24874 586294 24970 586350
rect 25026 586294 25094 586350
rect 25150 586294 25218 586350
rect 25274 586294 25342 586350
rect 25398 586294 25494 586350
rect 24874 586226 25494 586294
rect 24874 586170 24970 586226
rect 25026 586170 25094 586226
rect 25150 586170 25218 586226
rect 25274 586170 25342 586226
rect 25398 586170 25494 586226
rect 24874 586102 25494 586170
rect 24874 586046 24970 586102
rect 25026 586046 25094 586102
rect 25150 586046 25218 586102
rect 25274 586046 25342 586102
rect 25398 586046 25494 586102
rect 24874 585978 25494 586046
rect 24874 585922 24970 585978
rect 25026 585922 25094 585978
rect 25150 585922 25218 585978
rect 25274 585922 25342 585978
rect 25398 585922 25494 585978
rect 24874 568350 25494 585922
rect 37772 587188 37828 587198
rect 24874 568294 24970 568350
rect 25026 568294 25094 568350
rect 25150 568294 25218 568350
rect 25274 568294 25342 568350
rect 25398 568294 25494 568350
rect 24874 568226 25494 568294
rect 24874 568170 24970 568226
rect 25026 568170 25094 568226
rect 25150 568170 25218 568226
rect 25274 568170 25342 568226
rect 25398 568170 25494 568226
rect 24874 568102 25494 568170
rect 24874 568046 24970 568102
rect 25026 568046 25094 568102
rect 25150 568046 25218 568102
rect 25274 568046 25342 568102
rect 25398 568046 25494 568102
rect 24874 567978 25494 568046
rect 24874 567922 24970 567978
rect 25026 567922 25094 567978
rect 25150 567922 25218 567978
rect 25274 567922 25342 567978
rect 25398 567922 25494 567978
rect 24874 550350 25494 567922
rect 24874 550294 24970 550350
rect 25026 550294 25094 550350
rect 25150 550294 25218 550350
rect 25274 550294 25342 550350
rect 25398 550294 25494 550350
rect 24874 550226 25494 550294
rect 24874 550170 24970 550226
rect 25026 550170 25094 550226
rect 25150 550170 25218 550226
rect 25274 550170 25342 550226
rect 25398 550170 25494 550226
rect 24874 550102 25494 550170
rect 24874 550046 24970 550102
rect 25026 550046 25094 550102
rect 25150 550046 25218 550102
rect 25274 550046 25342 550102
rect 25398 550046 25494 550102
rect 24874 549978 25494 550046
rect 24874 549922 24970 549978
rect 25026 549922 25094 549978
rect 25150 549922 25218 549978
rect 25274 549922 25342 549978
rect 25398 549922 25494 549978
rect 24874 532350 25494 549922
rect 24874 532294 24970 532350
rect 25026 532294 25094 532350
rect 25150 532294 25218 532350
rect 25274 532294 25342 532350
rect 25398 532294 25494 532350
rect 24874 532226 25494 532294
rect 24874 532170 24970 532226
rect 25026 532170 25094 532226
rect 25150 532170 25218 532226
rect 25274 532170 25342 532226
rect 25398 532170 25494 532226
rect 24874 532102 25494 532170
rect 24874 532046 24970 532102
rect 25026 532046 25094 532102
rect 25150 532046 25218 532102
rect 25274 532046 25342 532102
rect 25398 532046 25494 532102
rect 24874 531978 25494 532046
rect 24874 531922 24970 531978
rect 25026 531922 25094 531978
rect 25150 531922 25218 531978
rect 25274 531922 25342 531978
rect 25398 531922 25494 531978
rect 21154 526294 21250 526350
rect 21306 526294 21374 526350
rect 21430 526294 21498 526350
rect 21554 526294 21622 526350
rect 21678 526294 21774 526350
rect 21154 526226 21774 526294
rect 21154 526170 21250 526226
rect 21306 526170 21374 526226
rect 21430 526170 21498 526226
rect 21554 526170 21622 526226
rect 21678 526170 21774 526226
rect 21154 526102 21774 526170
rect 21154 526046 21250 526102
rect 21306 526046 21374 526102
rect 21430 526046 21498 526102
rect 21554 526046 21622 526102
rect 21678 526046 21774 526102
rect 21154 525978 21774 526046
rect 21154 525922 21250 525978
rect 21306 525922 21374 525978
rect 21430 525922 21498 525978
rect 21554 525922 21622 525978
rect 21678 525922 21774 525978
rect 21154 508350 21774 525922
rect 21154 508294 21250 508350
rect 21306 508294 21374 508350
rect 21430 508294 21498 508350
rect 21554 508294 21622 508350
rect 21678 508294 21774 508350
rect 21154 508226 21774 508294
rect 21154 508170 21250 508226
rect 21306 508170 21374 508226
rect 21430 508170 21498 508226
rect 21554 508170 21622 508226
rect 21678 508170 21774 508226
rect 21154 508102 21774 508170
rect 21154 508046 21250 508102
rect 21306 508046 21374 508102
rect 21430 508046 21498 508102
rect 21554 508046 21622 508102
rect 21678 508046 21774 508102
rect 21154 507978 21774 508046
rect 21154 507922 21250 507978
rect 21306 507922 21374 507978
rect 21430 507922 21498 507978
rect 21554 507922 21622 507978
rect 21678 507922 21774 507978
rect 6874 496294 6970 496350
rect 7026 496294 7094 496350
rect 7150 496294 7218 496350
rect 7274 496294 7342 496350
rect 7398 496294 7494 496350
rect 6874 496226 7494 496294
rect 6874 496170 6970 496226
rect 7026 496170 7094 496226
rect 7150 496170 7218 496226
rect 7274 496170 7342 496226
rect 7398 496170 7494 496226
rect 6874 496102 7494 496170
rect 6874 496046 6970 496102
rect 7026 496046 7094 496102
rect 7150 496046 7218 496102
rect 7274 496046 7342 496102
rect 7398 496046 7494 496102
rect 6874 495978 7494 496046
rect 6874 495922 6970 495978
rect 7026 495922 7094 495978
rect 7150 495922 7218 495978
rect 7274 495922 7342 495978
rect 7398 495922 7494 495978
rect 6874 478350 7494 495922
rect 6874 478294 6970 478350
rect 7026 478294 7094 478350
rect 7150 478294 7218 478350
rect 7274 478294 7342 478350
rect 7398 478294 7494 478350
rect 6874 478226 7494 478294
rect 6874 478170 6970 478226
rect 7026 478170 7094 478226
rect 7150 478170 7218 478226
rect 7274 478170 7342 478226
rect 7398 478170 7494 478226
rect 6874 478102 7494 478170
rect 6874 478046 6970 478102
rect 7026 478046 7094 478102
rect 7150 478046 7218 478102
rect 7274 478046 7342 478102
rect 7398 478046 7494 478102
rect 6874 477978 7494 478046
rect 6874 477922 6970 477978
rect 7026 477922 7094 477978
rect 7150 477922 7218 477978
rect 7274 477922 7342 477978
rect 7398 477922 7494 477978
rect 5852 179442 5908 179452
rect 5964 474292 6020 474302
rect 5964 160468 6020 474236
rect 6874 460350 7494 477922
rect 6874 460294 6970 460350
rect 7026 460294 7094 460350
rect 7150 460294 7218 460350
rect 7274 460294 7342 460350
rect 7398 460294 7494 460350
rect 6874 460226 7494 460294
rect 6874 460170 6970 460226
rect 7026 460170 7094 460226
rect 7150 460170 7218 460226
rect 7274 460170 7342 460226
rect 7398 460170 7494 460226
rect 6874 460102 7494 460170
rect 6874 460046 6970 460102
rect 7026 460046 7094 460102
rect 7150 460046 7218 460102
rect 7274 460046 7342 460102
rect 7398 460046 7494 460102
rect 6874 459978 7494 460046
rect 6874 459922 6970 459978
rect 7026 459922 7094 459978
rect 7150 459922 7218 459978
rect 7274 459922 7342 459978
rect 7398 459922 7494 459978
rect 6874 442350 7494 459922
rect 6874 442294 6970 442350
rect 7026 442294 7094 442350
rect 7150 442294 7218 442350
rect 7274 442294 7342 442350
rect 7398 442294 7494 442350
rect 6874 442226 7494 442294
rect 6874 442170 6970 442226
rect 7026 442170 7094 442226
rect 7150 442170 7218 442226
rect 7274 442170 7342 442226
rect 7398 442170 7494 442226
rect 6874 442102 7494 442170
rect 6874 442046 6970 442102
rect 7026 442046 7094 442102
rect 7150 442046 7218 442102
rect 7274 442046 7342 442102
rect 7398 442046 7494 442102
rect 6874 441978 7494 442046
rect 6874 441922 6970 441978
rect 7026 441922 7094 441978
rect 7150 441922 7218 441978
rect 7274 441922 7342 441978
rect 7398 441922 7494 441978
rect 6874 424350 7494 441922
rect 6874 424294 6970 424350
rect 7026 424294 7094 424350
rect 7150 424294 7218 424350
rect 7274 424294 7342 424350
rect 7398 424294 7494 424350
rect 6874 424226 7494 424294
rect 6874 424170 6970 424226
rect 7026 424170 7094 424226
rect 7150 424170 7218 424226
rect 7274 424170 7342 424226
rect 7398 424170 7494 424226
rect 6874 424102 7494 424170
rect 6874 424046 6970 424102
rect 7026 424046 7094 424102
rect 7150 424046 7218 424102
rect 7274 424046 7342 424102
rect 7398 424046 7494 424102
rect 6874 423978 7494 424046
rect 6874 423922 6970 423978
rect 7026 423922 7094 423978
rect 7150 423922 7218 423978
rect 7274 423922 7342 423978
rect 7398 423922 7494 423978
rect 6874 406350 7494 423922
rect 6874 406294 6970 406350
rect 7026 406294 7094 406350
rect 7150 406294 7218 406350
rect 7274 406294 7342 406350
rect 7398 406294 7494 406350
rect 6874 406226 7494 406294
rect 6874 406170 6970 406226
rect 7026 406170 7094 406226
rect 7150 406170 7218 406226
rect 7274 406170 7342 406226
rect 7398 406170 7494 406226
rect 6874 406102 7494 406170
rect 6874 406046 6970 406102
rect 7026 406046 7094 406102
rect 7150 406046 7218 406102
rect 7274 406046 7342 406102
rect 7398 406046 7494 406102
rect 6874 405978 7494 406046
rect 6874 405922 6970 405978
rect 7026 405922 7094 405978
rect 7150 405922 7218 405978
rect 7274 405922 7342 405978
rect 7398 405922 7494 405978
rect 6874 388350 7494 405922
rect 12572 502516 12628 502526
rect 6874 388294 6970 388350
rect 7026 388294 7094 388350
rect 7150 388294 7218 388350
rect 7274 388294 7342 388350
rect 7398 388294 7494 388350
rect 6874 388226 7494 388294
rect 6874 388170 6970 388226
rect 7026 388170 7094 388226
rect 7150 388170 7218 388226
rect 7274 388170 7342 388226
rect 7398 388170 7494 388226
rect 6874 388102 7494 388170
rect 6874 388046 6970 388102
rect 7026 388046 7094 388102
rect 7150 388046 7218 388102
rect 7274 388046 7342 388102
rect 7398 388046 7494 388102
rect 6874 387978 7494 388046
rect 6874 387922 6970 387978
rect 7026 387922 7094 387978
rect 7150 387922 7218 387978
rect 7274 387922 7342 387978
rect 7398 387922 7494 387978
rect 6874 370350 7494 387922
rect 6874 370294 6970 370350
rect 7026 370294 7094 370350
rect 7150 370294 7218 370350
rect 7274 370294 7342 370350
rect 7398 370294 7494 370350
rect 6874 370226 7494 370294
rect 6874 370170 6970 370226
rect 7026 370170 7094 370226
rect 7150 370170 7218 370226
rect 7274 370170 7342 370226
rect 7398 370170 7494 370226
rect 6874 370102 7494 370170
rect 6874 370046 6970 370102
rect 7026 370046 7094 370102
rect 7150 370046 7218 370102
rect 7274 370046 7342 370102
rect 7398 370046 7494 370102
rect 6874 369978 7494 370046
rect 6874 369922 6970 369978
rect 7026 369922 7094 369978
rect 7150 369922 7218 369978
rect 7274 369922 7342 369978
rect 7398 369922 7494 369978
rect 6874 352350 7494 369922
rect 6874 352294 6970 352350
rect 7026 352294 7094 352350
rect 7150 352294 7218 352350
rect 7274 352294 7342 352350
rect 7398 352294 7494 352350
rect 6874 352226 7494 352294
rect 6874 352170 6970 352226
rect 7026 352170 7094 352226
rect 7150 352170 7218 352226
rect 7274 352170 7342 352226
rect 7398 352170 7494 352226
rect 6874 352102 7494 352170
rect 6874 352046 6970 352102
rect 7026 352046 7094 352102
rect 7150 352046 7218 352102
rect 7274 352046 7342 352102
rect 7398 352046 7494 352102
rect 6874 351978 7494 352046
rect 6874 351922 6970 351978
rect 7026 351922 7094 351978
rect 7150 351922 7218 351978
rect 7274 351922 7342 351978
rect 7398 351922 7494 351978
rect 6874 334350 7494 351922
rect 6874 334294 6970 334350
rect 7026 334294 7094 334350
rect 7150 334294 7218 334350
rect 7274 334294 7342 334350
rect 7398 334294 7494 334350
rect 6874 334226 7494 334294
rect 6874 334170 6970 334226
rect 7026 334170 7094 334226
rect 7150 334170 7218 334226
rect 7274 334170 7342 334226
rect 7398 334170 7494 334226
rect 6874 334102 7494 334170
rect 6874 334046 6970 334102
rect 7026 334046 7094 334102
rect 7150 334046 7218 334102
rect 7274 334046 7342 334102
rect 7398 334046 7494 334102
rect 6874 333978 7494 334046
rect 6874 333922 6970 333978
rect 7026 333922 7094 333978
rect 7150 333922 7218 333978
rect 7274 333922 7342 333978
rect 7398 333922 7494 333978
rect 6874 316350 7494 333922
rect 6874 316294 6970 316350
rect 7026 316294 7094 316350
rect 7150 316294 7218 316350
rect 7274 316294 7342 316350
rect 7398 316294 7494 316350
rect 6874 316226 7494 316294
rect 6874 316170 6970 316226
rect 7026 316170 7094 316226
rect 7150 316170 7218 316226
rect 7274 316170 7342 316226
rect 7398 316170 7494 316226
rect 6874 316102 7494 316170
rect 6874 316046 6970 316102
rect 7026 316046 7094 316102
rect 7150 316046 7218 316102
rect 7274 316046 7342 316102
rect 7398 316046 7494 316102
rect 6874 315978 7494 316046
rect 6874 315922 6970 315978
rect 7026 315922 7094 315978
rect 7150 315922 7218 315978
rect 7274 315922 7342 315978
rect 7398 315922 7494 315978
rect 6874 298350 7494 315922
rect 6874 298294 6970 298350
rect 7026 298294 7094 298350
rect 7150 298294 7218 298350
rect 7274 298294 7342 298350
rect 7398 298294 7494 298350
rect 6874 298226 7494 298294
rect 6874 298170 6970 298226
rect 7026 298170 7094 298226
rect 7150 298170 7218 298226
rect 7274 298170 7342 298226
rect 7398 298170 7494 298226
rect 6874 298102 7494 298170
rect 6874 298046 6970 298102
rect 7026 298046 7094 298102
rect 7150 298046 7218 298102
rect 7274 298046 7342 298102
rect 7398 298046 7494 298102
rect 6874 297978 7494 298046
rect 6874 297922 6970 297978
rect 7026 297922 7094 297978
rect 7150 297922 7218 297978
rect 7274 297922 7342 297978
rect 7398 297922 7494 297978
rect 6874 280350 7494 297922
rect 6874 280294 6970 280350
rect 7026 280294 7094 280350
rect 7150 280294 7218 280350
rect 7274 280294 7342 280350
rect 7398 280294 7494 280350
rect 6874 280226 7494 280294
rect 6874 280170 6970 280226
rect 7026 280170 7094 280226
rect 7150 280170 7218 280226
rect 7274 280170 7342 280226
rect 7398 280170 7494 280226
rect 6874 280102 7494 280170
rect 6874 280046 6970 280102
rect 7026 280046 7094 280102
rect 7150 280046 7218 280102
rect 7274 280046 7342 280102
rect 7398 280046 7494 280102
rect 6874 279978 7494 280046
rect 6874 279922 6970 279978
rect 7026 279922 7094 279978
rect 7150 279922 7218 279978
rect 7274 279922 7342 279978
rect 7398 279922 7494 279978
rect 5964 160402 6020 160412
rect 6076 262612 6132 262622
rect 6076 103348 6132 262556
rect 6076 103282 6132 103292
rect 6874 262350 7494 279922
rect 6874 262294 6970 262350
rect 7026 262294 7094 262350
rect 7150 262294 7218 262350
rect 7274 262294 7342 262350
rect 7398 262294 7494 262350
rect 6874 262226 7494 262294
rect 6874 262170 6970 262226
rect 7026 262170 7094 262226
rect 7150 262170 7218 262226
rect 7274 262170 7342 262226
rect 7398 262170 7494 262226
rect 6874 262102 7494 262170
rect 6874 262046 6970 262102
rect 7026 262046 7094 262102
rect 7150 262046 7218 262102
rect 7274 262046 7342 262102
rect 7398 262046 7494 262102
rect 6874 261978 7494 262046
rect 6874 261922 6970 261978
rect 7026 261922 7094 261978
rect 7150 261922 7218 261978
rect 7274 261922 7342 261978
rect 7398 261922 7494 261978
rect 6874 244350 7494 261922
rect 6874 244294 6970 244350
rect 7026 244294 7094 244350
rect 7150 244294 7218 244350
rect 7274 244294 7342 244350
rect 7398 244294 7494 244350
rect 6874 244226 7494 244294
rect 6874 244170 6970 244226
rect 7026 244170 7094 244226
rect 7150 244170 7218 244226
rect 7274 244170 7342 244226
rect 7398 244170 7494 244226
rect 6874 244102 7494 244170
rect 6874 244046 6970 244102
rect 7026 244046 7094 244102
rect 7150 244046 7218 244102
rect 7274 244046 7342 244102
rect 7398 244046 7494 244102
rect 6874 243978 7494 244046
rect 6874 243922 6970 243978
rect 7026 243922 7094 243978
rect 7150 243922 7218 243978
rect 7274 243922 7342 243978
rect 7398 243922 7494 243978
rect 6874 226350 7494 243922
rect 6874 226294 6970 226350
rect 7026 226294 7094 226350
rect 7150 226294 7218 226350
rect 7274 226294 7342 226350
rect 7398 226294 7494 226350
rect 6874 226226 7494 226294
rect 6874 226170 6970 226226
rect 7026 226170 7094 226226
rect 7150 226170 7218 226226
rect 7274 226170 7342 226226
rect 7398 226170 7494 226226
rect 6874 226102 7494 226170
rect 6874 226046 6970 226102
rect 7026 226046 7094 226102
rect 7150 226046 7218 226102
rect 7274 226046 7342 226102
rect 7398 226046 7494 226102
rect 6874 225978 7494 226046
rect 6874 225922 6970 225978
rect 7026 225922 7094 225978
rect 7150 225922 7218 225978
rect 7274 225922 7342 225978
rect 7398 225922 7494 225978
rect 6874 208350 7494 225922
rect 6874 208294 6970 208350
rect 7026 208294 7094 208350
rect 7150 208294 7218 208350
rect 7274 208294 7342 208350
rect 7398 208294 7494 208350
rect 6874 208226 7494 208294
rect 6874 208170 6970 208226
rect 7026 208170 7094 208226
rect 7150 208170 7218 208226
rect 7274 208170 7342 208226
rect 7398 208170 7494 208226
rect 6874 208102 7494 208170
rect 6874 208046 6970 208102
rect 7026 208046 7094 208102
rect 7150 208046 7218 208102
rect 7274 208046 7342 208102
rect 7398 208046 7494 208102
rect 6874 207978 7494 208046
rect 6874 207922 6970 207978
rect 7026 207922 7094 207978
rect 7150 207922 7218 207978
rect 7274 207922 7342 207978
rect 7398 207922 7494 207978
rect 6874 190350 7494 207922
rect 6874 190294 6970 190350
rect 7026 190294 7094 190350
rect 7150 190294 7218 190350
rect 7274 190294 7342 190350
rect 7398 190294 7494 190350
rect 6874 190226 7494 190294
rect 6874 190170 6970 190226
rect 7026 190170 7094 190226
rect 7150 190170 7218 190226
rect 7274 190170 7342 190226
rect 7398 190170 7494 190226
rect 6874 190102 7494 190170
rect 6874 190046 6970 190102
rect 7026 190046 7094 190102
rect 7150 190046 7218 190102
rect 7274 190046 7342 190102
rect 7398 190046 7494 190102
rect 6874 189978 7494 190046
rect 6874 189922 6970 189978
rect 7026 189922 7094 189978
rect 7150 189922 7218 189978
rect 7274 189922 7342 189978
rect 7398 189922 7494 189978
rect 6874 172350 7494 189922
rect 6874 172294 6970 172350
rect 7026 172294 7094 172350
rect 7150 172294 7218 172350
rect 7274 172294 7342 172350
rect 7398 172294 7494 172350
rect 6874 172226 7494 172294
rect 6874 172170 6970 172226
rect 7026 172170 7094 172226
rect 7150 172170 7218 172226
rect 7274 172170 7342 172226
rect 7398 172170 7494 172226
rect 6874 172102 7494 172170
rect 6874 172046 6970 172102
rect 7026 172046 7094 172102
rect 7150 172046 7218 172102
rect 7274 172046 7342 172102
rect 7398 172046 7494 172102
rect 6874 171978 7494 172046
rect 6874 171922 6970 171978
rect 7026 171922 7094 171978
rect 7150 171922 7218 171978
rect 7274 171922 7342 171978
rect 7398 171922 7494 171978
rect 6874 154350 7494 171922
rect 6874 154294 6970 154350
rect 7026 154294 7094 154350
rect 7150 154294 7218 154350
rect 7274 154294 7342 154350
rect 7398 154294 7494 154350
rect 6874 154226 7494 154294
rect 6874 154170 6970 154226
rect 7026 154170 7094 154226
rect 7150 154170 7218 154226
rect 7274 154170 7342 154226
rect 7398 154170 7494 154226
rect 6874 154102 7494 154170
rect 6874 154046 6970 154102
rect 7026 154046 7094 154102
rect 7150 154046 7218 154102
rect 7274 154046 7342 154102
rect 7398 154046 7494 154102
rect 6874 153978 7494 154046
rect 6874 153922 6970 153978
rect 7026 153922 7094 153978
rect 7150 153922 7218 153978
rect 7274 153922 7342 153978
rect 7398 153922 7494 153978
rect 6874 136350 7494 153922
rect 9212 389620 9268 389630
rect 9212 137620 9268 389564
rect 9212 137554 9268 137564
rect 9324 177940 9380 177950
rect 6874 136294 6970 136350
rect 7026 136294 7094 136350
rect 7150 136294 7218 136350
rect 7274 136294 7342 136350
rect 7398 136294 7494 136350
rect 6874 136226 7494 136294
rect 6874 136170 6970 136226
rect 7026 136170 7094 136226
rect 7150 136170 7218 136226
rect 7274 136170 7342 136226
rect 7398 136170 7494 136226
rect 6874 136102 7494 136170
rect 6874 136046 6970 136102
rect 7026 136046 7094 136102
rect 7150 136046 7218 136102
rect 7274 136046 7342 136102
rect 7398 136046 7494 136102
rect 6874 135978 7494 136046
rect 6874 135922 6970 135978
rect 7026 135922 7094 135978
rect 7150 135922 7218 135978
rect 7274 135922 7342 135978
rect 7398 135922 7494 135978
rect 6874 118350 7494 135922
rect 6874 118294 6970 118350
rect 7026 118294 7094 118350
rect 7150 118294 7218 118350
rect 7274 118294 7342 118350
rect 7398 118294 7494 118350
rect 6874 118226 7494 118294
rect 6874 118170 6970 118226
rect 7026 118170 7094 118226
rect 7150 118170 7218 118226
rect 7274 118170 7342 118226
rect 7398 118170 7494 118226
rect 6874 118102 7494 118170
rect 6874 118046 6970 118102
rect 7026 118046 7094 118102
rect 7150 118046 7218 118102
rect 7274 118046 7342 118102
rect 7398 118046 7494 118102
rect 6874 117978 7494 118046
rect 6874 117922 6970 117978
rect 7026 117922 7094 117978
rect 7150 117922 7218 117978
rect 7274 117922 7342 117978
rect 7398 117922 7494 117978
rect 6874 100350 7494 117922
rect 6874 100294 6970 100350
rect 7026 100294 7094 100350
rect 7150 100294 7218 100350
rect 7274 100294 7342 100350
rect 7398 100294 7494 100350
rect 6874 100226 7494 100294
rect 6874 100170 6970 100226
rect 7026 100170 7094 100226
rect 7150 100170 7218 100226
rect 7274 100170 7342 100226
rect 7398 100170 7494 100226
rect 6874 100102 7494 100170
rect 6874 100046 6970 100102
rect 7026 100046 7094 100102
rect 7150 100046 7218 100102
rect 7274 100046 7342 100102
rect 7398 100046 7494 100102
rect 6874 99978 7494 100046
rect 6874 99922 6970 99978
rect 7026 99922 7094 99978
rect 7150 99922 7218 99978
rect 7274 99922 7342 99978
rect 7398 99922 7494 99978
rect 4396 91858 4452 91868
rect 5852 93268 5908 93278
rect 4284 61394 4340 61404
rect 4396 79156 4452 79166
rect 4396 53844 4452 79100
rect 5852 59668 5908 93212
rect 5852 59602 5908 59612
rect 6874 82350 7494 99922
rect 6874 82294 6970 82350
rect 7026 82294 7094 82350
rect 7150 82294 7218 82350
rect 7274 82294 7342 82350
rect 7398 82294 7494 82350
rect 6874 82226 7494 82294
rect 6874 82170 6970 82226
rect 7026 82170 7094 82226
rect 7150 82170 7218 82226
rect 7274 82170 7342 82226
rect 7398 82170 7494 82226
rect 6874 82102 7494 82170
rect 6874 82046 6970 82102
rect 7026 82046 7094 82102
rect 7150 82046 7218 82102
rect 7274 82046 7342 82102
rect 7398 82046 7494 82102
rect 6874 81978 7494 82046
rect 6874 81922 6970 81978
rect 7026 81922 7094 81978
rect 7150 81922 7218 81978
rect 7274 81922 7342 81978
rect 7398 81922 7494 81978
rect 6874 64350 7494 81922
rect 9324 80500 9380 177884
rect 12572 168084 12628 502460
rect 21154 490350 21774 507922
rect 21154 490294 21250 490350
rect 21306 490294 21374 490350
rect 21430 490294 21498 490350
rect 21554 490294 21622 490350
rect 21678 490294 21774 490350
rect 21154 490226 21774 490294
rect 21154 490170 21250 490226
rect 21306 490170 21374 490226
rect 21430 490170 21498 490226
rect 21554 490170 21622 490226
rect 21678 490170 21774 490226
rect 21154 490102 21774 490170
rect 21154 490046 21250 490102
rect 21306 490046 21374 490102
rect 21430 490046 21498 490102
rect 21554 490046 21622 490102
rect 21678 490046 21774 490102
rect 21154 489978 21774 490046
rect 21154 489922 21250 489978
rect 21306 489922 21374 489978
rect 21430 489922 21498 489978
rect 21554 489922 21622 489978
rect 21678 489922 21774 489978
rect 21154 472350 21774 489922
rect 21154 472294 21250 472350
rect 21306 472294 21374 472350
rect 21430 472294 21498 472350
rect 21554 472294 21622 472350
rect 21678 472294 21774 472350
rect 21154 472226 21774 472294
rect 21154 472170 21250 472226
rect 21306 472170 21374 472226
rect 21430 472170 21498 472226
rect 21554 472170 21622 472226
rect 21678 472170 21774 472226
rect 21154 472102 21774 472170
rect 21154 472046 21250 472102
rect 21306 472046 21374 472102
rect 21430 472046 21498 472102
rect 21554 472046 21622 472102
rect 21678 472046 21774 472102
rect 21154 471978 21774 472046
rect 21154 471922 21250 471978
rect 21306 471922 21374 471978
rect 21430 471922 21498 471978
rect 21554 471922 21622 471978
rect 21678 471922 21774 471978
rect 12572 168018 12628 168028
rect 14252 460180 14308 460190
rect 12572 163828 12628 163838
rect 9324 80434 9380 80444
rect 10892 149716 10948 149726
rect 10892 72884 10948 149660
rect 12572 84868 12628 163772
rect 14252 156660 14308 460124
rect 21154 454350 21774 471922
rect 21154 454294 21250 454350
rect 21306 454294 21374 454350
rect 21430 454294 21498 454350
rect 21554 454294 21622 454350
rect 21678 454294 21774 454350
rect 21154 454226 21774 454294
rect 21154 454170 21250 454226
rect 21306 454170 21374 454226
rect 21430 454170 21498 454226
rect 21554 454170 21622 454226
rect 21678 454170 21774 454226
rect 21154 454102 21774 454170
rect 21154 454046 21250 454102
rect 21306 454046 21374 454102
rect 21430 454046 21498 454102
rect 21554 454046 21622 454102
rect 21678 454046 21774 454102
rect 21154 453978 21774 454046
rect 21154 453922 21250 453978
rect 21306 453922 21374 453978
rect 21430 453922 21498 453978
rect 21554 453922 21622 453978
rect 21678 453922 21774 453978
rect 19292 446068 19348 446078
rect 14252 156594 14308 156604
rect 15932 417844 15988 417854
rect 15932 145236 15988 417788
rect 15932 145170 15988 145180
rect 17612 375508 17668 375518
rect 17612 133812 17668 375452
rect 19292 152852 19348 446012
rect 21154 436350 21774 453922
rect 21154 436294 21250 436350
rect 21306 436294 21374 436350
rect 21430 436294 21498 436350
rect 21554 436294 21622 436350
rect 21678 436294 21774 436350
rect 21154 436226 21774 436294
rect 21154 436170 21250 436226
rect 21306 436170 21374 436226
rect 21430 436170 21498 436226
rect 21554 436170 21622 436226
rect 21678 436170 21774 436226
rect 21154 436102 21774 436170
rect 21154 436046 21250 436102
rect 21306 436046 21374 436102
rect 21430 436046 21498 436102
rect 21554 436046 21622 436102
rect 21678 436046 21774 436102
rect 21154 435978 21774 436046
rect 21154 435922 21250 435978
rect 21306 435922 21374 435978
rect 21430 435922 21498 435978
rect 21554 435922 21622 435978
rect 21678 435922 21774 435978
rect 21154 418350 21774 435922
rect 21154 418294 21250 418350
rect 21306 418294 21374 418350
rect 21430 418294 21498 418350
rect 21554 418294 21622 418350
rect 21678 418294 21774 418350
rect 21154 418226 21774 418294
rect 21154 418170 21250 418226
rect 21306 418170 21374 418226
rect 21430 418170 21498 418226
rect 21554 418170 21622 418226
rect 21678 418170 21774 418226
rect 21154 418102 21774 418170
rect 21154 418046 21250 418102
rect 21306 418046 21374 418102
rect 21430 418046 21498 418102
rect 21554 418046 21622 418102
rect 21678 418046 21774 418102
rect 21154 417978 21774 418046
rect 21154 417922 21250 417978
rect 21306 417922 21374 417978
rect 21430 417922 21498 417978
rect 21554 417922 21622 417978
rect 21678 417922 21774 417978
rect 21154 400350 21774 417922
rect 21154 400294 21250 400350
rect 21306 400294 21374 400350
rect 21430 400294 21498 400350
rect 21554 400294 21622 400350
rect 21678 400294 21774 400350
rect 21154 400226 21774 400294
rect 21154 400170 21250 400226
rect 21306 400170 21374 400226
rect 21430 400170 21498 400226
rect 21554 400170 21622 400226
rect 21678 400170 21774 400226
rect 21154 400102 21774 400170
rect 21154 400046 21250 400102
rect 21306 400046 21374 400102
rect 21430 400046 21498 400102
rect 21554 400046 21622 400102
rect 21678 400046 21774 400102
rect 21154 399978 21774 400046
rect 21154 399922 21250 399978
rect 21306 399922 21374 399978
rect 21430 399922 21498 399978
rect 21554 399922 21622 399978
rect 21678 399922 21774 399978
rect 21154 382350 21774 399922
rect 21154 382294 21250 382350
rect 21306 382294 21374 382350
rect 21430 382294 21498 382350
rect 21554 382294 21622 382350
rect 21678 382294 21774 382350
rect 21154 382226 21774 382294
rect 21154 382170 21250 382226
rect 21306 382170 21374 382226
rect 21430 382170 21498 382226
rect 21554 382170 21622 382226
rect 21678 382170 21774 382226
rect 21154 382102 21774 382170
rect 21154 382046 21250 382102
rect 21306 382046 21374 382102
rect 21430 382046 21498 382102
rect 21554 382046 21622 382102
rect 21678 382046 21774 382102
rect 21154 381978 21774 382046
rect 21154 381922 21250 381978
rect 21306 381922 21374 381978
rect 21430 381922 21498 381978
rect 21554 381922 21622 381978
rect 21678 381922 21774 381978
rect 21154 364350 21774 381922
rect 21154 364294 21250 364350
rect 21306 364294 21374 364350
rect 21430 364294 21498 364350
rect 21554 364294 21622 364350
rect 21678 364294 21774 364350
rect 21154 364226 21774 364294
rect 21154 364170 21250 364226
rect 21306 364170 21374 364226
rect 21430 364170 21498 364226
rect 21554 364170 21622 364226
rect 21678 364170 21774 364226
rect 21154 364102 21774 364170
rect 21154 364046 21250 364102
rect 21306 364046 21374 364102
rect 21430 364046 21498 364102
rect 21554 364046 21622 364102
rect 21678 364046 21774 364102
rect 21154 363978 21774 364046
rect 21154 363922 21250 363978
rect 21306 363922 21374 363978
rect 21430 363922 21498 363978
rect 21554 363922 21622 363978
rect 21678 363922 21774 363978
rect 21154 346350 21774 363922
rect 21154 346294 21250 346350
rect 21306 346294 21374 346350
rect 21430 346294 21498 346350
rect 21554 346294 21622 346350
rect 21678 346294 21774 346350
rect 21154 346226 21774 346294
rect 21154 346170 21250 346226
rect 21306 346170 21374 346226
rect 21430 346170 21498 346226
rect 21554 346170 21622 346226
rect 21678 346170 21774 346226
rect 21154 346102 21774 346170
rect 21154 346046 21250 346102
rect 21306 346046 21374 346102
rect 21430 346046 21498 346102
rect 21554 346046 21622 346102
rect 21678 346046 21774 346102
rect 21154 345978 21774 346046
rect 21154 345922 21250 345978
rect 21306 345922 21374 345978
rect 21430 345922 21498 345978
rect 21554 345922 21622 345978
rect 21678 345922 21774 345978
rect 19292 152786 19348 152796
rect 19404 333172 19460 333182
rect 17612 133746 17668 133756
rect 19404 122388 19460 333116
rect 19404 122322 19460 122332
rect 21154 328350 21774 345922
rect 21154 328294 21250 328350
rect 21306 328294 21374 328350
rect 21430 328294 21498 328350
rect 21554 328294 21622 328350
rect 21678 328294 21774 328350
rect 21154 328226 21774 328294
rect 21154 328170 21250 328226
rect 21306 328170 21374 328226
rect 21430 328170 21498 328226
rect 21554 328170 21622 328226
rect 21678 328170 21774 328226
rect 21154 328102 21774 328170
rect 21154 328046 21250 328102
rect 21306 328046 21374 328102
rect 21430 328046 21498 328102
rect 21554 328046 21622 328102
rect 21678 328046 21774 328102
rect 21154 327978 21774 328046
rect 21154 327922 21250 327978
rect 21306 327922 21374 327978
rect 21430 327922 21498 327978
rect 21554 327922 21622 327978
rect 21678 327922 21774 327978
rect 21154 310350 21774 327922
rect 21154 310294 21250 310350
rect 21306 310294 21374 310350
rect 21430 310294 21498 310350
rect 21554 310294 21622 310350
rect 21678 310294 21774 310350
rect 21154 310226 21774 310294
rect 21154 310170 21250 310226
rect 21306 310170 21374 310226
rect 21430 310170 21498 310226
rect 21554 310170 21622 310226
rect 21678 310170 21774 310226
rect 21154 310102 21774 310170
rect 21154 310046 21250 310102
rect 21306 310046 21374 310102
rect 21430 310046 21498 310102
rect 21554 310046 21622 310102
rect 21678 310046 21774 310102
rect 21154 309978 21774 310046
rect 21154 309922 21250 309978
rect 21306 309922 21374 309978
rect 21430 309922 21498 309978
rect 21554 309922 21622 309978
rect 21678 309922 21774 309978
rect 21154 292350 21774 309922
rect 21154 292294 21250 292350
rect 21306 292294 21374 292350
rect 21430 292294 21498 292350
rect 21554 292294 21622 292350
rect 21678 292294 21774 292350
rect 21154 292226 21774 292294
rect 21154 292170 21250 292226
rect 21306 292170 21374 292226
rect 21430 292170 21498 292226
rect 21554 292170 21622 292226
rect 21678 292170 21774 292226
rect 21154 292102 21774 292170
rect 21154 292046 21250 292102
rect 21306 292046 21374 292102
rect 21430 292046 21498 292102
rect 21554 292046 21622 292102
rect 21678 292046 21774 292102
rect 21154 291978 21774 292046
rect 21154 291922 21250 291978
rect 21306 291922 21374 291978
rect 21430 291922 21498 291978
rect 21554 291922 21622 291978
rect 21678 291922 21774 291978
rect 21154 274350 21774 291922
rect 21154 274294 21250 274350
rect 21306 274294 21374 274350
rect 21430 274294 21498 274350
rect 21554 274294 21622 274350
rect 21678 274294 21774 274350
rect 21154 274226 21774 274294
rect 21154 274170 21250 274226
rect 21306 274170 21374 274226
rect 21430 274170 21498 274226
rect 21554 274170 21622 274226
rect 21678 274170 21774 274226
rect 21154 274102 21774 274170
rect 21154 274046 21250 274102
rect 21306 274046 21374 274102
rect 21430 274046 21498 274102
rect 21554 274046 21622 274102
rect 21678 274046 21774 274102
rect 21154 273978 21774 274046
rect 21154 273922 21250 273978
rect 21306 273922 21374 273978
rect 21430 273922 21498 273978
rect 21554 273922 21622 273978
rect 21678 273922 21774 273978
rect 21154 256350 21774 273922
rect 21154 256294 21250 256350
rect 21306 256294 21374 256350
rect 21430 256294 21498 256350
rect 21554 256294 21622 256350
rect 21678 256294 21774 256350
rect 21154 256226 21774 256294
rect 21154 256170 21250 256226
rect 21306 256170 21374 256226
rect 21430 256170 21498 256226
rect 21554 256170 21622 256226
rect 21678 256170 21774 256226
rect 21154 256102 21774 256170
rect 21154 256046 21250 256102
rect 21306 256046 21374 256102
rect 21430 256046 21498 256102
rect 21554 256046 21622 256102
rect 21678 256046 21774 256102
rect 21154 255978 21774 256046
rect 21154 255922 21250 255978
rect 21306 255922 21374 255978
rect 21430 255922 21498 255978
rect 21554 255922 21622 255978
rect 21678 255922 21774 255978
rect 21154 238350 21774 255922
rect 21154 238294 21250 238350
rect 21306 238294 21374 238350
rect 21430 238294 21498 238350
rect 21554 238294 21622 238350
rect 21678 238294 21774 238350
rect 21154 238226 21774 238294
rect 21154 238170 21250 238226
rect 21306 238170 21374 238226
rect 21430 238170 21498 238226
rect 21554 238170 21622 238226
rect 21678 238170 21774 238226
rect 21154 238102 21774 238170
rect 21154 238046 21250 238102
rect 21306 238046 21374 238102
rect 21430 238046 21498 238102
rect 21554 238046 21622 238102
rect 21678 238046 21774 238102
rect 21154 237978 21774 238046
rect 21154 237922 21250 237978
rect 21306 237922 21374 237978
rect 21430 237922 21498 237978
rect 21554 237922 21622 237978
rect 21678 237922 21774 237978
rect 21154 220350 21774 237922
rect 21154 220294 21250 220350
rect 21306 220294 21374 220350
rect 21430 220294 21498 220350
rect 21554 220294 21622 220350
rect 21678 220294 21774 220350
rect 21154 220226 21774 220294
rect 21154 220170 21250 220226
rect 21306 220170 21374 220226
rect 21430 220170 21498 220226
rect 21554 220170 21622 220226
rect 21678 220170 21774 220226
rect 21154 220102 21774 220170
rect 21154 220046 21250 220102
rect 21306 220046 21374 220102
rect 21430 220046 21498 220102
rect 21554 220046 21622 220102
rect 21678 220046 21774 220102
rect 21154 219978 21774 220046
rect 21154 219922 21250 219978
rect 21306 219922 21374 219978
rect 21430 219922 21498 219978
rect 21554 219922 21622 219978
rect 21678 219922 21774 219978
rect 21154 202350 21774 219922
rect 21154 202294 21250 202350
rect 21306 202294 21374 202350
rect 21430 202294 21498 202350
rect 21554 202294 21622 202350
rect 21678 202294 21774 202350
rect 21154 202226 21774 202294
rect 21154 202170 21250 202226
rect 21306 202170 21374 202226
rect 21430 202170 21498 202226
rect 21554 202170 21622 202226
rect 21678 202170 21774 202226
rect 21154 202102 21774 202170
rect 21154 202046 21250 202102
rect 21306 202046 21374 202102
rect 21430 202046 21498 202102
rect 21554 202046 21622 202102
rect 21678 202046 21774 202102
rect 21154 201978 21774 202046
rect 21154 201922 21250 201978
rect 21306 201922 21374 201978
rect 21430 201922 21498 201978
rect 21554 201922 21622 201978
rect 21678 201922 21774 201978
rect 21154 184350 21774 201922
rect 21154 184294 21250 184350
rect 21306 184294 21374 184350
rect 21430 184294 21498 184350
rect 21554 184294 21622 184350
rect 21678 184294 21774 184350
rect 21154 184226 21774 184294
rect 21154 184170 21250 184226
rect 21306 184170 21374 184226
rect 21430 184170 21498 184226
rect 21554 184170 21622 184226
rect 21678 184170 21774 184226
rect 21154 184102 21774 184170
rect 21154 184046 21250 184102
rect 21306 184046 21374 184102
rect 21430 184046 21498 184102
rect 21554 184046 21622 184102
rect 21678 184046 21774 184102
rect 21154 183978 21774 184046
rect 21154 183922 21250 183978
rect 21306 183922 21374 183978
rect 21430 183922 21498 183978
rect 21554 183922 21622 183978
rect 21678 183922 21774 183978
rect 21154 166350 21774 183922
rect 22652 530740 22708 530750
rect 22652 175700 22708 530684
rect 24874 514350 25494 531922
rect 24874 514294 24970 514350
rect 25026 514294 25094 514350
rect 25150 514294 25218 514350
rect 25274 514294 25342 514350
rect 25398 514294 25494 514350
rect 24874 514226 25494 514294
rect 24874 514170 24970 514226
rect 25026 514170 25094 514226
rect 25150 514170 25218 514226
rect 25274 514170 25342 514226
rect 25398 514170 25494 514226
rect 24874 514102 25494 514170
rect 24874 514046 24970 514102
rect 25026 514046 25094 514102
rect 25150 514046 25218 514102
rect 25274 514046 25342 514102
rect 25398 514046 25494 514102
rect 24874 513978 25494 514046
rect 24874 513922 24970 513978
rect 25026 513922 25094 513978
rect 25150 513922 25218 513978
rect 25274 513922 25342 513978
rect 25398 513922 25494 513978
rect 24874 496350 25494 513922
rect 24874 496294 24970 496350
rect 25026 496294 25094 496350
rect 25150 496294 25218 496350
rect 25274 496294 25342 496350
rect 25398 496294 25494 496350
rect 24874 496226 25494 496294
rect 24874 496170 24970 496226
rect 25026 496170 25094 496226
rect 25150 496170 25218 496226
rect 25274 496170 25342 496226
rect 25398 496170 25494 496226
rect 24874 496102 25494 496170
rect 24874 496046 24970 496102
rect 25026 496046 25094 496102
rect 25150 496046 25218 496102
rect 25274 496046 25342 496102
rect 25398 496046 25494 496102
rect 24874 495978 25494 496046
rect 24874 495922 24970 495978
rect 25026 495922 25094 495978
rect 25150 495922 25218 495978
rect 25274 495922 25342 495978
rect 25398 495922 25494 495978
rect 24874 478350 25494 495922
rect 24874 478294 24970 478350
rect 25026 478294 25094 478350
rect 25150 478294 25218 478350
rect 25274 478294 25342 478350
rect 25398 478294 25494 478350
rect 24874 478226 25494 478294
rect 24874 478170 24970 478226
rect 25026 478170 25094 478226
rect 25150 478170 25218 478226
rect 25274 478170 25342 478226
rect 25398 478170 25494 478226
rect 24874 478102 25494 478170
rect 24874 478046 24970 478102
rect 25026 478046 25094 478102
rect 25150 478046 25218 478102
rect 25274 478046 25342 478102
rect 25398 478046 25494 478102
rect 24874 477978 25494 478046
rect 24874 477922 24970 477978
rect 25026 477922 25094 477978
rect 25150 477922 25218 477978
rect 25274 477922 25342 477978
rect 25398 477922 25494 477978
rect 24874 460350 25494 477922
rect 24874 460294 24970 460350
rect 25026 460294 25094 460350
rect 25150 460294 25218 460350
rect 25274 460294 25342 460350
rect 25398 460294 25494 460350
rect 24874 460226 25494 460294
rect 24874 460170 24970 460226
rect 25026 460170 25094 460226
rect 25150 460170 25218 460226
rect 25274 460170 25342 460226
rect 25398 460170 25494 460226
rect 24874 460102 25494 460170
rect 24874 460046 24970 460102
rect 25026 460046 25094 460102
rect 25150 460046 25218 460102
rect 25274 460046 25342 460102
rect 25398 460046 25494 460102
rect 24874 459978 25494 460046
rect 24874 459922 24970 459978
rect 25026 459922 25094 459978
rect 25150 459922 25218 459978
rect 25274 459922 25342 459978
rect 25398 459922 25494 459978
rect 24874 442350 25494 459922
rect 24874 442294 24970 442350
rect 25026 442294 25094 442350
rect 25150 442294 25218 442350
rect 25274 442294 25342 442350
rect 25398 442294 25494 442350
rect 24874 442226 25494 442294
rect 24874 442170 24970 442226
rect 25026 442170 25094 442226
rect 25150 442170 25218 442226
rect 25274 442170 25342 442226
rect 25398 442170 25494 442226
rect 24874 442102 25494 442170
rect 24874 442046 24970 442102
rect 25026 442046 25094 442102
rect 25150 442046 25218 442102
rect 25274 442046 25342 442102
rect 25398 442046 25494 442102
rect 24874 441978 25494 442046
rect 24874 441922 24970 441978
rect 25026 441922 25094 441978
rect 25150 441922 25218 441978
rect 25274 441922 25342 441978
rect 25398 441922 25494 441978
rect 24874 424350 25494 441922
rect 24874 424294 24970 424350
rect 25026 424294 25094 424350
rect 25150 424294 25218 424350
rect 25274 424294 25342 424350
rect 25398 424294 25494 424350
rect 24874 424226 25494 424294
rect 24874 424170 24970 424226
rect 25026 424170 25094 424226
rect 25150 424170 25218 424226
rect 25274 424170 25342 424226
rect 25398 424170 25494 424226
rect 24874 424102 25494 424170
rect 24874 424046 24970 424102
rect 25026 424046 25094 424102
rect 25150 424046 25218 424102
rect 25274 424046 25342 424102
rect 25398 424046 25494 424102
rect 24874 423978 25494 424046
rect 24874 423922 24970 423978
rect 25026 423922 25094 423978
rect 25150 423922 25218 423978
rect 25274 423922 25342 423978
rect 25398 423922 25494 423978
rect 24874 406350 25494 423922
rect 24874 406294 24970 406350
rect 25026 406294 25094 406350
rect 25150 406294 25218 406350
rect 25274 406294 25342 406350
rect 25398 406294 25494 406350
rect 24874 406226 25494 406294
rect 24874 406170 24970 406226
rect 25026 406170 25094 406226
rect 25150 406170 25218 406226
rect 25274 406170 25342 406226
rect 25398 406170 25494 406226
rect 24874 406102 25494 406170
rect 24874 406046 24970 406102
rect 25026 406046 25094 406102
rect 25150 406046 25218 406102
rect 25274 406046 25342 406102
rect 25398 406046 25494 406102
rect 24874 405978 25494 406046
rect 24874 405922 24970 405978
rect 25026 405922 25094 405978
rect 25150 405922 25218 405978
rect 25274 405922 25342 405978
rect 25398 405922 25494 405978
rect 24874 388350 25494 405922
rect 24874 388294 24970 388350
rect 25026 388294 25094 388350
rect 25150 388294 25218 388350
rect 25274 388294 25342 388350
rect 25398 388294 25494 388350
rect 24874 388226 25494 388294
rect 24874 388170 24970 388226
rect 25026 388170 25094 388226
rect 25150 388170 25218 388226
rect 25274 388170 25342 388226
rect 25398 388170 25494 388226
rect 24874 388102 25494 388170
rect 24874 388046 24970 388102
rect 25026 388046 25094 388102
rect 25150 388046 25218 388102
rect 25274 388046 25342 388102
rect 25398 388046 25494 388102
rect 24874 387978 25494 388046
rect 24874 387922 24970 387978
rect 25026 387922 25094 387978
rect 25150 387922 25218 387978
rect 25274 387922 25342 387978
rect 25398 387922 25494 387978
rect 24874 370350 25494 387922
rect 24874 370294 24970 370350
rect 25026 370294 25094 370350
rect 25150 370294 25218 370350
rect 25274 370294 25342 370350
rect 25398 370294 25494 370350
rect 24874 370226 25494 370294
rect 24874 370170 24970 370226
rect 25026 370170 25094 370226
rect 25150 370170 25218 370226
rect 25274 370170 25342 370226
rect 25398 370170 25494 370226
rect 24874 370102 25494 370170
rect 24874 370046 24970 370102
rect 25026 370046 25094 370102
rect 25150 370046 25218 370102
rect 25274 370046 25342 370102
rect 25398 370046 25494 370102
rect 24874 369978 25494 370046
rect 24874 369922 24970 369978
rect 25026 369922 25094 369978
rect 25150 369922 25218 369978
rect 25274 369922 25342 369978
rect 25398 369922 25494 369978
rect 24874 352350 25494 369922
rect 24874 352294 24970 352350
rect 25026 352294 25094 352350
rect 25150 352294 25218 352350
rect 25274 352294 25342 352350
rect 25398 352294 25494 352350
rect 24874 352226 25494 352294
rect 24874 352170 24970 352226
rect 25026 352170 25094 352226
rect 25150 352170 25218 352226
rect 25274 352170 25342 352226
rect 25398 352170 25494 352226
rect 24874 352102 25494 352170
rect 24874 352046 24970 352102
rect 25026 352046 25094 352102
rect 25150 352046 25218 352102
rect 25274 352046 25342 352102
rect 25398 352046 25494 352102
rect 24874 351978 25494 352046
rect 24874 351922 24970 351978
rect 25026 351922 25094 351978
rect 25150 351922 25218 351978
rect 25274 351922 25342 351978
rect 25398 351922 25494 351978
rect 24874 334350 25494 351922
rect 24874 334294 24970 334350
rect 25026 334294 25094 334350
rect 25150 334294 25218 334350
rect 25274 334294 25342 334350
rect 25398 334294 25494 334350
rect 24874 334226 25494 334294
rect 24874 334170 24970 334226
rect 25026 334170 25094 334226
rect 25150 334170 25218 334226
rect 25274 334170 25342 334226
rect 25398 334170 25494 334226
rect 24874 334102 25494 334170
rect 24874 334046 24970 334102
rect 25026 334046 25094 334102
rect 25150 334046 25218 334102
rect 25274 334046 25342 334102
rect 25398 334046 25494 334102
rect 24874 333978 25494 334046
rect 24874 333922 24970 333978
rect 25026 333922 25094 333978
rect 25150 333922 25218 333978
rect 25274 333922 25342 333978
rect 25398 333922 25494 333978
rect 24874 316350 25494 333922
rect 24874 316294 24970 316350
rect 25026 316294 25094 316350
rect 25150 316294 25218 316350
rect 25274 316294 25342 316350
rect 25398 316294 25494 316350
rect 24874 316226 25494 316294
rect 24874 316170 24970 316226
rect 25026 316170 25094 316226
rect 25150 316170 25218 316226
rect 25274 316170 25342 316226
rect 25398 316170 25494 316226
rect 24874 316102 25494 316170
rect 24874 316046 24970 316102
rect 25026 316046 25094 316102
rect 25150 316046 25218 316102
rect 25274 316046 25342 316102
rect 25398 316046 25494 316102
rect 24874 315978 25494 316046
rect 24874 315922 24970 315978
rect 25026 315922 25094 315978
rect 25150 315922 25218 315978
rect 25274 315922 25342 315978
rect 25398 315922 25494 315978
rect 24874 298350 25494 315922
rect 24874 298294 24970 298350
rect 25026 298294 25094 298350
rect 25150 298294 25218 298350
rect 25274 298294 25342 298350
rect 25398 298294 25494 298350
rect 24874 298226 25494 298294
rect 24874 298170 24970 298226
rect 25026 298170 25094 298226
rect 25150 298170 25218 298226
rect 25274 298170 25342 298226
rect 25398 298170 25494 298226
rect 24874 298102 25494 298170
rect 24874 298046 24970 298102
rect 25026 298046 25094 298102
rect 25150 298046 25218 298102
rect 25274 298046 25342 298102
rect 25398 298046 25494 298102
rect 24874 297978 25494 298046
rect 24874 297922 24970 297978
rect 25026 297922 25094 297978
rect 25150 297922 25218 297978
rect 25274 297922 25342 297978
rect 25398 297922 25494 297978
rect 22652 175634 22708 175644
rect 22764 290836 22820 290846
rect 21154 166294 21250 166350
rect 21306 166294 21374 166350
rect 21430 166294 21498 166350
rect 21554 166294 21622 166350
rect 21678 166294 21774 166350
rect 21154 166226 21774 166294
rect 21154 166170 21250 166226
rect 21306 166170 21374 166226
rect 21430 166170 21498 166226
rect 21554 166170 21622 166226
rect 21678 166170 21774 166226
rect 21154 166102 21774 166170
rect 21154 166046 21250 166102
rect 21306 166046 21374 166102
rect 21430 166046 21498 166102
rect 21554 166046 21622 166102
rect 21678 166046 21774 166102
rect 21154 165978 21774 166046
rect 21154 165922 21250 165978
rect 21306 165922 21374 165978
rect 21430 165922 21498 165978
rect 21554 165922 21622 165978
rect 21678 165922 21774 165978
rect 21154 148350 21774 165922
rect 21154 148294 21250 148350
rect 21306 148294 21374 148350
rect 21430 148294 21498 148350
rect 21554 148294 21622 148350
rect 21678 148294 21774 148350
rect 21154 148226 21774 148294
rect 21154 148170 21250 148226
rect 21306 148170 21374 148226
rect 21430 148170 21498 148226
rect 21554 148170 21622 148226
rect 21678 148170 21774 148226
rect 21154 148102 21774 148170
rect 21154 148046 21250 148102
rect 21306 148046 21374 148102
rect 21430 148046 21498 148102
rect 21554 148046 21622 148102
rect 21678 148046 21774 148102
rect 21154 147978 21774 148046
rect 21154 147922 21250 147978
rect 21306 147922 21374 147978
rect 21430 147922 21498 147978
rect 21554 147922 21622 147978
rect 21678 147922 21774 147978
rect 21154 130350 21774 147922
rect 21154 130294 21250 130350
rect 21306 130294 21374 130350
rect 21430 130294 21498 130350
rect 21554 130294 21622 130350
rect 21678 130294 21774 130350
rect 21154 130226 21774 130294
rect 21154 130170 21250 130226
rect 21306 130170 21374 130226
rect 21430 130170 21498 130226
rect 21554 130170 21622 130226
rect 21678 130170 21774 130226
rect 21154 130102 21774 130170
rect 21154 130046 21250 130102
rect 21306 130046 21374 130102
rect 21430 130046 21498 130102
rect 21554 130046 21622 130102
rect 21678 130046 21774 130102
rect 21154 129978 21774 130046
rect 21154 129922 21250 129978
rect 21306 129922 21374 129978
rect 21430 129922 21498 129978
rect 21554 129922 21622 129978
rect 21678 129922 21774 129978
rect 12572 84802 12628 84812
rect 14252 121492 14308 121502
rect 10892 72818 10948 72828
rect 14252 68068 14308 121436
rect 14252 68002 14308 68012
rect 21154 112350 21774 129922
rect 22764 113428 22820 290780
rect 22764 113362 22820 113372
rect 24874 280350 25494 297922
rect 24874 280294 24970 280350
rect 25026 280294 25094 280350
rect 25150 280294 25218 280350
rect 25274 280294 25342 280350
rect 25398 280294 25494 280350
rect 24874 280226 25494 280294
rect 24874 280170 24970 280226
rect 25026 280170 25094 280226
rect 25150 280170 25218 280226
rect 25274 280170 25342 280226
rect 25398 280170 25494 280226
rect 24874 280102 25494 280170
rect 24874 280046 24970 280102
rect 25026 280046 25094 280102
rect 25150 280046 25218 280102
rect 25274 280046 25342 280102
rect 25398 280046 25494 280102
rect 24874 279978 25494 280046
rect 24874 279922 24970 279978
rect 25026 279922 25094 279978
rect 25150 279922 25218 279978
rect 25274 279922 25342 279978
rect 25398 279922 25494 279978
rect 24874 262350 25494 279922
rect 24874 262294 24970 262350
rect 25026 262294 25094 262350
rect 25150 262294 25218 262350
rect 25274 262294 25342 262350
rect 25398 262294 25494 262350
rect 24874 262226 25494 262294
rect 24874 262170 24970 262226
rect 25026 262170 25094 262226
rect 25150 262170 25218 262226
rect 25274 262170 25342 262226
rect 25398 262170 25494 262226
rect 24874 262102 25494 262170
rect 24874 262046 24970 262102
rect 25026 262046 25094 262102
rect 25150 262046 25218 262102
rect 25274 262046 25342 262102
rect 25398 262046 25494 262102
rect 24874 261978 25494 262046
rect 24874 261922 24970 261978
rect 25026 261922 25094 261978
rect 25150 261922 25218 261978
rect 25274 261922 25342 261978
rect 25398 261922 25494 261978
rect 24874 244350 25494 261922
rect 24874 244294 24970 244350
rect 25026 244294 25094 244350
rect 25150 244294 25218 244350
rect 25274 244294 25342 244350
rect 25398 244294 25494 244350
rect 24874 244226 25494 244294
rect 24874 244170 24970 244226
rect 25026 244170 25094 244226
rect 25150 244170 25218 244226
rect 25274 244170 25342 244226
rect 25398 244170 25494 244226
rect 24874 244102 25494 244170
rect 24874 244046 24970 244102
rect 25026 244046 25094 244102
rect 25150 244046 25218 244102
rect 25274 244046 25342 244102
rect 25398 244046 25494 244102
rect 24874 243978 25494 244046
rect 24874 243922 24970 243978
rect 25026 243922 25094 243978
rect 25150 243922 25218 243978
rect 25274 243922 25342 243978
rect 25398 243922 25494 243978
rect 24874 226350 25494 243922
rect 24874 226294 24970 226350
rect 25026 226294 25094 226350
rect 25150 226294 25218 226350
rect 25274 226294 25342 226350
rect 25398 226294 25494 226350
rect 24874 226226 25494 226294
rect 24874 226170 24970 226226
rect 25026 226170 25094 226226
rect 25150 226170 25218 226226
rect 25274 226170 25342 226226
rect 25398 226170 25494 226226
rect 24874 226102 25494 226170
rect 24874 226046 24970 226102
rect 25026 226046 25094 226102
rect 25150 226046 25218 226102
rect 25274 226046 25342 226102
rect 25398 226046 25494 226102
rect 24874 225978 25494 226046
rect 24874 225922 24970 225978
rect 25026 225922 25094 225978
rect 25150 225922 25218 225978
rect 25274 225922 25342 225978
rect 25398 225922 25494 225978
rect 24874 208350 25494 225922
rect 24874 208294 24970 208350
rect 25026 208294 25094 208350
rect 25150 208294 25218 208350
rect 25274 208294 25342 208350
rect 25398 208294 25494 208350
rect 24874 208226 25494 208294
rect 24874 208170 24970 208226
rect 25026 208170 25094 208226
rect 25150 208170 25218 208226
rect 25274 208170 25342 208226
rect 25398 208170 25494 208226
rect 24874 208102 25494 208170
rect 24874 208046 24970 208102
rect 25026 208046 25094 208102
rect 25150 208046 25218 208102
rect 25274 208046 25342 208102
rect 25398 208046 25494 208102
rect 24874 207978 25494 208046
rect 24874 207922 24970 207978
rect 25026 207922 25094 207978
rect 25150 207922 25218 207978
rect 25274 207922 25342 207978
rect 25398 207922 25494 207978
rect 24874 190350 25494 207922
rect 24874 190294 24970 190350
rect 25026 190294 25094 190350
rect 25150 190294 25218 190350
rect 25274 190294 25342 190350
rect 25398 190294 25494 190350
rect 24874 190226 25494 190294
rect 24874 190170 24970 190226
rect 25026 190170 25094 190226
rect 25150 190170 25218 190226
rect 25274 190170 25342 190226
rect 25398 190170 25494 190226
rect 24874 190102 25494 190170
rect 24874 190046 24970 190102
rect 25026 190046 25094 190102
rect 25150 190046 25218 190102
rect 25274 190046 25342 190102
rect 25398 190046 25494 190102
rect 24874 189978 25494 190046
rect 24874 189922 24970 189978
rect 25026 189922 25094 189978
rect 25150 189922 25218 189978
rect 25274 189922 25342 189978
rect 25398 189922 25494 189978
rect 24874 172350 25494 189922
rect 27692 573076 27748 573086
rect 27692 187124 27748 573020
rect 36092 558964 36148 558974
rect 34412 516628 34468 516638
rect 31052 431956 31108 431966
rect 29372 347284 29428 347294
rect 27692 187058 27748 187068
rect 27804 248500 27860 248510
rect 24874 172294 24970 172350
rect 25026 172294 25094 172350
rect 25150 172294 25218 172350
rect 25274 172294 25342 172350
rect 25398 172294 25494 172350
rect 24874 172226 25494 172294
rect 24874 172170 24970 172226
rect 25026 172170 25094 172226
rect 25150 172170 25218 172226
rect 25274 172170 25342 172226
rect 25398 172170 25494 172226
rect 24874 172102 25494 172170
rect 24874 172046 24970 172102
rect 25026 172046 25094 172102
rect 25150 172046 25218 172102
rect 25274 172046 25342 172102
rect 25398 172046 25494 172102
rect 24874 171978 25494 172046
rect 24874 171922 24970 171978
rect 25026 171922 25094 171978
rect 25150 171922 25218 171978
rect 25274 171922 25342 171978
rect 25398 171922 25494 171978
rect 24874 154350 25494 171922
rect 24874 154294 24970 154350
rect 25026 154294 25094 154350
rect 25150 154294 25218 154350
rect 25274 154294 25342 154350
rect 25398 154294 25494 154350
rect 24874 154226 25494 154294
rect 24874 154170 24970 154226
rect 25026 154170 25094 154226
rect 25150 154170 25218 154226
rect 25274 154170 25342 154226
rect 25398 154170 25494 154226
rect 24874 154102 25494 154170
rect 24874 154046 24970 154102
rect 25026 154046 25094 154102
rect 25150 154046 25218 154102
rect 25274 154046 25342 154102
rect 25398 154046 25494 154102
rect 24874 153978 25494 154046
rect 24874 153922 24970 153978
rect 25026 153922 25094 153978
rect 25150 153922 25218 153978
rect 25274 153922 25342 153978
rect 25398 153922 25494 153978
rect 24874 136350 25494 153922
rect 24874 136294 24970 136350
rect 25026 136294 25094 136350
rect 25150 136294 25218 136350
rect 25274 136294 25342 136350
rect 25398 136294 25494 136350
rect 24874 136226 25494 136294
rect 24874 136170 24970 136226
rect 25026 136170 25094 136226
rect 25150 136170 25218 136226
rect 25274 136170 25342 136226
rect 25398 136170 25494 136226
rect 24874 136102 25494 136170
rect 24874 136046 24970 136102
rect 25026 136046 25094 136102
rect 25150 136046 25218 136102
rect 25274 136046 25342 136102
rect 25398 136046 25494 136102
rect 24874 135978 25494 136046
rect 24874 135922 24970 135978
rect 25026 135922 25094 135978
rect 25150 135922 25218 135978
rect 25274 135922 25342 135978
rect 25398 135922 25494 135978
rect 24874 118350 25494 135922
rect 24874 118294 24970 118350
rect 25026 118294 25094 118350
rect 25150 118294 25218 118350
rect 25274 118294 25342 118350
rect 25398 118294 25494 118350
rect 24874 118226 25494 118294
rect 24874 118170 24970 118226
rect 25026 118170 25094 118226
rect 25150 118170 25218 118226
rect 25274 118170 25342 118226
rect 25398 118170 25494 118226
rect 24874 118102 25494 118170
rect 24874 118046 24970 118102
rect 25026 118046 25094 118102
rect 25150 118046 25218 118102
rect 25274 118046 25342 118102
rect 25398 118046 25494 118102
rect 24874 117978 25494 118046
rect 24874 117922 24970 117978
rect 25026 117922 25094 117978
rect 25150 117922 25218 117978
rect 25274 117922 25342 117978
rect 25398 117922 25494 117978
rect 21154 112294 21250 112350
rect 21306 112294 21374 112350
rect 21430 112294 21498 112350
rect 21554 112294 21622 112350
rect 21678 112294 21774 112350
rect 21154 112226 21774 112294
rect 21154 112170 21250 112226
rect 21306 112170 21374 112226
rect 21430 112170 21498 112226
rect 21554 112170 21622 112226
rect 21678 112170 21774 112226
rect 21154 112102 21774 112170
rect 21154 112046 21250 112102
rect 21306 112046 21374 112102
rect 21430 112046 21498 112102
rect 21554 112046 21622 112102
rect 21678 112046 21774 112102
rect 21154 111978 21774 112046
rect 21154 111922 21250 111978
rect 21306 111922 21374 111978
rect 21430 111922 21498 111978
rect 21554 111922 21622 111978
rect 21678 111922 21774 111978
rect 21154 94350 21774 111922
rect 21154 94294 21250 94350
rect 21306 94294 21374 94350
rect 21430 94294 21498 94350
rect 21554 94294 21622 94350
rect 21678 94294 21774 94350
rect 21154 94226 21774 94294
rect 21154 94170 21250 94226
rect 21306 94170 21374 94226
rect 21430 94170 21498 94226
rect 21554 94170 21622 94226
rect 21678 94170 21774 94226
rect 21154 94102 21774 94170
rect 21154 94046 21250 94102
rect 21306 94046 21374 94102
rect 21430 94046 21498 94102
rect 21554 94046 21622 94102
rect 21678 94046 21774 94102
rect 21154 93978 21774 94046
rect 21154 93922 21250 93978
rect 21306 93922 21374 93978
rect 21430 93922 21498 93978
rect 21554 93922 21622 93978
rect 21678 93922 21774 93978
rect 21154 76350 21774 93922
rect 21154 76294 21250 76350
rect 21306 76294 21374 76350
rect 21430 76294 21498 76350
rect 21554 76294 21622 76350
rect 21678 76294 21774 76350
rect 21154 76226 21774 76294
rect 21154 76170 21250 76226
rect 21306 76170 21374 76226
rect 21430 76170 21498 76226
rect 21554 76170 21622 76226
rect 21678 76170 21774 76226
rect 21154 76102 21774 76170
rect 21154 76046 21250 76102
rect 21306 76046 21374 76102
rect 21430 76046 21498 76102
rect 21554 76046 21622 76102
rect 21678 76046 21774 76102
rect 21154 75978 21774 76046
rect 21154 75922 21250 75978
rect 21306 75922 21374 75978
rect 21430 75922 21498 75978
rect 21554 75922 21622 75978
rect 21678 75922 21774 75978
rect 6874 64294 6970 64350
rect 7026 64294 7094 64350
rect 7150 64294 7218 64350
rect 7274 64294 7342 64350
rect 7398 64294 7494 64350
rect 6874 64226 7494 64294
rect 6874 64170 6970 64226
rect 7026 64170 7094 64226
rect 7150 64170 7218 64226
rect 7274 64170 7342 64226
rect 7398 64170 7494 64226
rect 6874 64102 7494 64170
rect 6874 64046 6970 64102
rect 7026 64046 7094 64102
rect 7150 64046 7218 64102
rect 7274 64046 7342 64102
rect 7398 64046 7494 64102
rect 6874 63978 7494 64046
rect 6874 63922 6970 63978
rect 7026 63922 7094 63978
rect 7150 63922 7218 63978
rect 7274 63922 7342 63978
rect 7398 63922 7494 63978
rect 4396 53778 4452 53788
rect 4172 49970 4228 49980
rect 5068 50932 5124 50942
rect 5068 47908 5124 50876
rect 5068 47842 5124 47852
rect 6874 46350 7494 63922
rect 6874 46294 6970 46350
rect 7026 46294 7094 46350
rect 7150 46294 7218 46350
rect 7274 46294 7342 46350
rect 7398 46294 7494 46350
rect 6874 46226 7494 46294
rect 6874 46170 6970 46226
rect 7026 46170 7094 46226
rect 7150 46170 7218 46226
rect 7274 46170 7342 46226
rect 7398 46170 7494 46226
rect 6874 46102 7494 46170
rect 6874 46046 6970 46102
rect 7026 46046 7094 46102
rect 7150 46046 7218 46102
rect 7274 46046 7342 46102
rect 7398 46046 7494 46102
rect 6874 45978 7494 46046
rect 6874 45922 6970 45978
rect 7026 45922 7094 45978
rect 7150 45922 7218 45978
rect 7274 45922 7342 45978
rect 7398 45922 7494 45978
rect 3154 40294 3250 40350
rect 3306 40294 3374 40350
rect 3430 40294 3498 40350
rect 3554 40294 3622 40350
rect 3678 40294 3774 40350
rect 3154 40226 3774 40294
rect 3154 40170 3250 40226
rect 3306 40170 3374 40226
rect 3430 40170 3498 40226
rect 3554 40170 3622 40226
rect 3678 40170 3774 40226
rect 3154 40102 3774 40170
rect 3154 40046 3250 40102
rect 3306 40046 3374 40102
rect 3430 40046 3498 40102
rect 3554 40046 3622 40102
rect 3678 40046 3774 40102
rect 3154 39978 3774 40046
rect 3154 39922 3250 39978
rect 3306 39922 3374 39978
rect 3430 39922 3498 39978
rect 3554 39922 3622 39978
rect 3678 39922 3774 39978
rect 3154 22350 3774 39922
rect 4172 42420 4228 42430
rect 4172 36932 4228 42364
rect 4172 36866 4228 36876
rect 4284 38612 4340 38622
rect 3154 22294 3250 22350
rect 3306 22294 3374 22350
rect 3430 22294 3498 22350
rect 3554 22294 3622 22350
rect 3678 22294 3774 22350
rect 3154 22226 3774 22294
rect 3154 22170 3250 22226
rect 3306 22170 3374 22226
rect 3430 22170 3498 22226
rect 3554 22170 3622 22226
rect 3678 22170 3774 22226
rect 3154 22102 3774 22170
rect 3154 22046 3250 22102
rect 3306 22046 3374 22102
rect 3430 22046 3498 22102
rect 3554 22046 3622 22102
rect 3678 22046 3774 22102
rect 3154 21978 3774 22046
rect 3154 21922 3250 21978
rect 3306 21922 3374 21978
rect 3430 21922 3498 21978
rect 3554 21922 3622 21978
rect 3678 21922 3774 21978
rect 3154 4350 3774 21922
rect 4172 34804 4228 34814
rect 4172 8820 4228 34748
rect 4284 22932 4340 38556
rect 4284 22866 4340 22876
rect 6874 28350 7494 45922
rect 6874 28294 6970 28350
rect 7026 28294 7094 28350
rect 7150 28294 7218 28350
rect 7274 28294 7342 28350
rect 7398 28294 7494 28350
rect 6874 28226 7494 28294
rect 6874 28170 6970 28226
rect 7026 28170 7094 28226
rect 7150 28170 7218 28226
rect 7274 28170 7342 28226
rect 7398 28170 7494 28226
rect 6874 28102 7494 28170
rect 6874 28046 6970 28102
rect 7026 28046 7094 28102
rect 7150 28046 7218 28102
rect 7274 28046 7342 28102
rect 7398 28046 7494 28102
rect 6874 27978 7494 28046
rect 6874 27922 6970 27978
rect 7026 27922 7094 27978
rect 7150 27922 7218 27978
rect 7274 27922 7342 27978
rect 7398 27922 7494 27978
rect 4172 8754 4228 8764
rect 6874 10350 7494 27922
rect 6874 10294 6970 10350
rect 7026 10294 7094 10350
rect 7150 10294 7218 10350
rect 7274 10294 7342 10350
rect 7398 10294 7494 10350
rect 6874 10226 7494 10294
rect 6874 10170 6970 10226
rect 7026 10170 7094 10226
rect 7150 10170 7218 10226
rect 7274 10170 7342 10226
rect 7398 10170 7494 10226
rect 6874 10102 7494 10170
rect 6874 10046 6970 10102
rect 7026 10046 7094 10102
rect 7150 10046 7218 10102
rect 7274 10046 7342 10102
rect 7398 10046 7494 10102
rect 6874 9978 7494 10046
rect 6874 9922 6970 9978
rect 7026 9922 7094 9978
rect 7150 9922 7218 9978
rect 7274 9922 7342 9978
rect 7398 9922 7494 9978
rect 3154 4294 3250 4350
rect 3306 4294 3374 4350
rect 3430 4294 3498 4350
rect 3554 4294 3622 4350
rect 3678 4294 3774 4350
rect 3154 4226 3774 4294
rect 3154 4170 3250 4226
rect 3306 4170 3374 4226
rect 3430 4170 3498 4226
rect 3554 4170 3622 4226
rect 3678 4170 3774 4226
rect 3154 4102 3774 4170
rect 3154 4046 3250 4102
rect 3306 4046 3374 4102
rect 3430 4046 3498 4102
rect 3554 4046 3622 4102
rect 3678 4046 3774 4102
rect 3154 3978 3774 4046
rect 3154 3922 3250 3978
rect 3306 3922 3374 3978
rect 3430 3922 3498 3978
rect 3554 3922 3622 3978
rect 3678 3922 3774 3978
rect 3154 -160 3774 3922
rect 3154 -216 3250 -160
rect 3306 -216 3374 -160
rect 3430 -216 3498 -160
rect 3554 -216 3622 -160
rect 3678 -216 3774 -160
rect 3154 -284 3774 -216
rect 3154 -340 3250 -284
rect 3306 -340 3374 -284
rect 3430 -340 3498 -284
rect 3554 -340 3622 -284
rect 3678 -340 3774 -284
rect 3154 -408 3774 -340
rect 3154 -464 3250 -408
rect 3306 -464 3374 -408
rect 3430 -464 3498 -408
rect 3554 -464 3622 -408
rect 3678 -464 3774 -408
rect 3154 -532 3774 -464
rect 3154 -588 3250 -532
rect 3306 -588 3374 -532
rect 3430 -588 3498 -532
rect 3554 -588 3622 -532
rect 3678 -588 3774 -532
rect -1916 -1176 -1820 -1120
rect -1764 -1176 -1696 -1120
rect -1640 -1176 -1572 -1120
rect -1516 -1176 -1448 -1120
rect -1392 -1176 -1296 -1120
rect -1916 -1244 -1296 -1176
rect -1916 -1300 -1820 -1244
rect -1764 -1300 -1696 -1244
rect -1640 -1300 -1572 -1244
rect -1516 -1300 -1448 -1244
rect -1392 -1300 -1296 -1244
rect -1916 -1368 -1296 -1300
rect -1916 -1424 -1820 -1368
rect -1764 -1424 -1696 -1368
rect -1640 -1424 -1572 -1368
rect -1516 -1424 -1448 -1368
rect -1392 -1424 -1296 -1368
rect -1916 -1492 -1296 -1424
rect -1916 -1548 -1820 -1492
rect -1764 -1548 -1696 -1492
rect -1640 -1548 -1572 -1492
rect -1516 -1548 -1448 -1492
rect -1392 -1548 -1296 -1492
rect -1916 -1644 -1296 -1548
rect 3154 -1644 3774 -588
rect 6874 -1120 7494 9922
rect 6874 -1176 6970 -1120
rect 7026 -1176 7094 -1120
rect 7150 -1176 7218 -1120
rect 7274 -1176 7342 -1120
rect 7398 -1176 7494 -1120
rect 6874 -1244 7494 -1176
rect 6874 -1300 6970 -1244
rect 7026 -1300 7094 -1244
rect 7150 -1300 7218 -1244
rect 7274 -1300 7342 -1244
rect 7398 -1300 7494 -1244
rect 6874 -1368 7494 -1300
rect 6874 -1424 6970 -1368
rect 7026 -1424 7094 -1368
rect 7150 -1424 7218 -1368
rect 7274 -1424 7342 -1368
rect 7398 -1424 7494 -1368
rect 6874 -1492 7494 -1424
rect 6874 -1548 6970 -1492
rect 7026 -1548 7094 -1492
rect 7150 -1548 7218 -1492
rect 7274 -1548 7342 -1492
rect 7398 -1548 7494 -1492
rect 6874 -1644 7494 -1548
rect 21154 58350 21774 75922
rect 21154 58294 21250 58350
rect 21306 58294 21374 58350
rect 21430 58294 21498 58350
rect 21554 58294 21622 58350
rect 21678 58294 21774 58350
rect 21154 58226 21774 58294
rect 21154 58170 21250 58226
rect 21306 58170 21374 58226
rect 21430 58170 21498 58226
rect 21554 58170 21622 58226
rect 21678 58170 21774 58226
rect 21154 58102 21774 58170
rect 21154 58046 21250 58102
rect 21306 58046 21374 58102
rect 21430 58046 21498 58102
rect 21554 58046 21622 58102
rect 21678 58046 21774 58102
rect 21154 57978 21774 58046
rect 21154 57922 21250 57978
rect 21306 57922 21374 57978
rect 21430 57922 21498 57978
rect 21554 57922 21622 57978
rect 21678 57922 21774 57978
rect 21154 40350 21774 57922
rect 21154 40294 21250 40350
rect 21306 40294 21374 40350
rect 21430 40294 21498 40350
rect 21554 40294 21622 40350
rect 21678 40294 21774 40350
rect 21154 40226 21774 40294
rect 21154 40170 21250 40226
rect 21306 40170 21374 40226
rect 21430 40170 21498 40226
rect 21554 40170 21622 40226
rect 21678 40170 21774 40226
rect 21154 40102 21774 40170
rect 21154 40046 21250 40102
rect 21306 40046 21374 40102
rect 21430 40046 21498 40102
rect 21554 40046 21622 40102
rect 21678 40046 21774 40102
rect 21154 39978 21774 40046
rect 21154 39922 21250 39978
rect 21306 39922 21374 39978
rect 21430 39922 21498 39978
rect 21554 39922 21622 39978
rect 21678 39922 21774 39978
rect 21154 22350 21774 39922
rect 21154 22294 21250 22350
rect 21306 22294 21374 22350
rect 21430 22294 21498 22350
rect 21554 22294 21622 22350
rect 21678 22294 21774 22350
rect 21154 22226 21774 22294
rect 21154 22170 21250 22226
rect 21306 22170 21374 22226
rect 21430 22170 21498 22226
rect 21554 22170 21622 22226
rect 21678 22170 21774 22226
rect 21154 22102 21774 22170
rect 21154 22046 21250 22102
rect 21306 22046 21374 22102
rect 21430 22046 21498 22102
rect 21554 22046 21622 22102
rect 21678 22046 21774 22102
rect 21154 21978 21774 22046
rect 21154 21922 21250 21978
rect 21306 21922 21374 21978
rect 21430 21922 21498 21978
rect 21554 21922 21622 21978
rect 21678 21922 21774 21978
rect 21154 4350 21774 21922
rect 21154 4294 21250 4350
rect 21306 4294 21374 4350
rect 21430 4294 21498 4350
rect 21554 4294 21622 4350
rect 21678 4294 21774 4350
rect 21154 4226 21774 4294
rect 21154 4170 21250 4226
rect 21306 4170 21374 4226
rect 21430 4170 21498 4226
rect 21554 4170 21622 4226
rect 21678 4170 21774 4226
rect 21154 4102 21774 4170
rect 21154 4046 21250 4102
rect 21306 4046 21374 4102
rect 21430 4046 21498 4102
rect 21554 4046 21622 4102
rect 21678 4046 21774 4102
rect 21154 3978 21774 4046
rect 21154 3922 21250 3978
rect 21306 3922 21374 3978
rect 21430 3922 21498 3978
rect 21554 3922 21622 3978
rect 21678 3922 21774 3978
rect 21154 -160 21774 3922
rect 21154 -216 21250 -160
rect 21306 -216 21374 -160
rect 21430 -216 21498 -160
rect 21554 -216 21622 -160
rect 21678 -216 21774 -160
rect 21154 -284 21774 -216
rect 21154 -340 21250 -284
rect 21306 -340 21374 -284
rect 21430 -340 21498 -284
rect 21554 -340 21622 -284
rect 21678 -340 21774 -284
rect 21154 -408 21774 -340
rect 21154 -464 21250 -408
rect 21306 -464 21374 -408
rect 21430 -464 21498 -408
rect 21554 -464 21622 -408
rect 21678 -464 21774 -408
rect 21154 -532 21774 -464
rect 21154 -588 21250 -532
rect 21306 -588 21374 -532
rect 21430 -588 21498 -532
rect 21554 -588 21622 -532
rect 21678 -588 21774 -532
rect 21154 -1644 21774 -588
rect 24874 100350 25494 117922
rect 27804 101668 27860 248444
rect 29372 126196 29428 347228
rect 29372 126130 29428 126140
rect 29484 206164 29540 206174
rect 27804 101602 27860 101612
rect 24874 100294 24970 100350
rect 25026 100294 25094 100350
rect 25150 100294 25218 100350
rect 25274 100294 25342 100350
rect 25398 100294 25494 100350
rect 24874 100226 25494 100294
rect 24874 100170 24970 100226
rect 25026 100170 25094 100226
rect 25150 100170 25218 100226
rect 25274 100170 25342 100226
rect 25398 100170 25494 100226
rect 24874 100102 25494 100170
rect 24874 100046 24970 100102
rect 25026 100046 25094 100102
rect 25150 100046 25218 100102
rect 25274 100046 25342 100102
rect 25398 100046 25494 100102
rect 24874 99978 25494 100046
rect 24874 99922 24970 99978
rect 25026 99922 25094 99978
rect 25150 99922 25218 99978
rect 25274 99922 25342 99978
rect 25398 99922 25494 99978
rect 24874 82350 25494 99922
rect 29484 88116 29540 206108
rect 31052 150388 31108 431900
rect 31052 150322 31108 150332
rect 32732 304948 32788 304958
rect 32732 114772 32788 304892
rect 34412 171892 34468 516572
rect 34412 171826 34468 171836
rect 34524 276724 34580 276734
rect 32732 114706 32788 114716
rect 34524 107156 34580 276668
rect 36092 183316 36148 558908
rect 36092 183250 36148 183260
rect 36204 319060 36260 319070
rect 36204 120148 36260 319004
rect 37772 190932 37828 587132
rect 39154 580350 39774 596784
rect 39154 580294 39250 580350
rect 39306 580294 39374 580350
rect 39430 580294 39498 580350
rect 39554 580294 39622 580350
rect 39678 580294 39774 580350
rect 39154 580226 39774 580294
rect 39154 580170 39250 580226
rect 39306 580170 39374 580226
rect 39430 580170 39498 580226
rect 39554 580170 39622 580226
rect 39678 580170 39774 580226
rect 39154 580102 39774 580170
rect 39154 580046 39250 580102
rect 39306 580046 39374 580102
rect 39430 580046 39498 580102
rect 39554 580046 39622 580102
rect 39678 580046 39774 580102
rect 39154 579978 39774 580046
rect 39154 579922 39250 579978
rect 39306 579922 39374 579978
rect 39430 579922 39498 579978
rect 39554 579922 39622 579978
rect 39678 579922 39774 579978
rect 39154 562350 39774 579922
rect 39154 562294 39250 562350
rect 39306 562294 39374 562350
rect 39430 562294 39498 562350
rect 39554 562294 39622 562350
rect 39678 562294 39774 562350
rect 39154 562226 39774 562294
rect 39154 562170 39250 562226
rect 39306 562170 39374 562226
rect 39430 562170 39498 562226
rect 39554 562170 39622 562226
rect 39678 562170 39774 562226
rect 39154 562102 39774 562170
rect 39154 562046 39250 562102
rect 39306 562046 39374 562102
rect 39430 562046 39498 562102
rect 39554 562046 39622 562102
rect 39678 562046 39774 562102
rect 39154 561978 39774 562046
rect 39154 561922 39250 561978
rect 39306 561922 39374 561978
rect 39430 561922 39498 561978
rect 39554 561922 39622 561978
rect 39678 561922 39774 561978
rect 39154 544350 39774 561922
rect 39154 544294 39250 544350
rect 39306 544294 39374 544350
rect 39430 544294 39498 544350
rect 39554 544294 39622 544350
rect 39678 544294 39774 544350
rect 39154 544226 39774 544294
rect 39154 544170 39250 544226
rect 39306 544170 39374 544226
rect 39430 544170 39498 544226
rect 39554 544170 39622 544226
rect 39678 544170 39774 544226
rect 39154 544102 39774 544170
rect 39154 544046 39250 544102
rect 39306 544046 39374 544102
rect 39430 544046 39498 544102
rect 39554 544046 39622 544102
rect 39678 544046 39774 544102
rect 39154 543978 39774 544046
rect 39154 543922 39250 543978
rect 39306 543922 39374 543978
rect 39430 543922 39498 543978
rect 39554 543922 39622 543978
rect 39678 543922 39774 543978
rect 39154 526350 39774 543922
rect 39154 526294 39250 526350
rect 39306 526294 39374 526350
rect 39430 526294 39498 526350
rect 39554 526294 39622 526350
rect 39678 526294 39774 526350
rect 39154 526226 39774 526294
rect 39154 526170 39250 526226
rect 39306 526170 39374 526226
rect 39430 526170 39498 526226
rect 39554 526170 39622 526226
rect 39678 526170 39774 526226
rect 39154 526102 39774 526170
rect 39154 526046 39250 526102
rect 39306 526046 39374 526102
rect 39430 526046 39498 526102
rect 39554 526046 39622 526102
rect 39678 526046 39774 526102
rect 39154 525978 39774 526046
rect 39154 525922 39250 525978
rect 39306 525922 39374 525978
rect 39430 525922 39498 525978
rect 39554 525922 39622 525978
rect 39678 525922 39774 525978
rect 39154 508350 39774 525922
rect 39154 508294 39250 508350
rect 39306 508294 39374 508350
rect 39430 508294 39498 508350
rect 39554 508294 39622 508350
rect 39678 508294 39774 508350
rect 39154 508226 39774 508294
rect 39154 508170 39250 508226
rect 39306 508170 39374 508226
rect 39430 508170 39498 508226
rect 39554 508170 39622 508226
rect 39678 508170 39774 508226
rect 39154 508102 39774 508170
rect 39154 508046 39250 508102
rect 39306 508046 39374 508102
rect 39430 508046 39498 508102
rect 39554 508046 39622 508102
rect 39678 508046 39774 508102
rect 39154 507978 39774 508046
rect 39154 507922 39250 507978
rect 39306 507922 39374 507978
rect 39430 507922 39498 507978
rect 39554 507922 39622 507978
rect 39678 507922 39774 507978
rect 39154 490350 39774 507922
rect 39154 490294 39250 490350
rect 39306 490294 39374 490350
rect 39430 490294 39498 490350
rect 39554 490294 39622 490350
rect 39678 490294 39774 490350
rect 39154 490226 39774 490294
rect 39154 490170 39250 490226
rect 39306 490170 39374 490226
rect 39430 490170 39498 490226
rect 39554 490170 39622 490226
rect 39678 490170 39774 490226
rect 39154 490102 39774 490170
rect 39154 490046 39250 490102
rect 39306 490046 39374 490102
rect 39430 490046 39498 490102
rect 39554 490046 39622 490102
rect 39678 490046 39774 490102
rect 39154 489978 39774 490046
rect 39154 489922 39250 489978
rect 39306 489922 39374 489978
rect 39430 489922 39498 489978
rect 39554 489922 39622 489978
rect 39678 489922 39774 489978
rect 39154 472350 39774 489922
rect 39154 472294 39250 472350
rect 39306 472294 39374 472350
rect 39430 472294 39498 472350
rect 39554 472294 39622 472350
rect 39678 472294 39774 472350
rect 39154 472226 39774 472294
rect 39154 472170 39250 472226
rect 39306 472170 39374 472226
rect 39430 472170 39498 472226
rect 39554 472170 39622 472226
rect 39678 472170 39774 472226
rect 39154 472102 39774 472170
rect 39154 472046 39250 472102
rect 39306 472046 39374 472102
rect 39430 472046 39498 472102
rect 39554 472046 39622 472102
rect 39678 472046 39774 472102
rect 39154 471978 39774 472046
rect 39154 471922 39250 471978
rect 39306 471922 39374 471978
rect 39430 471922 39498 471978
rect 39554 471922 39622 471978
rect 39678 471922 39774 471978
rect 39154 454350 39774 471922
rect 39154 454294 39250 454350
rect 39306 454294 39374 454350
rect 39430 454294 39498 454350
rect 39554 454294 39622 454350
rect 39678 454294 39774 454350
rect 39154 454226 39774 454294
rect 39154 454170 39250 454226
rect 39306 454170 39374 454226
rect 39430 454170 39498 454226
rect 39554 454170 39622 454226
rect 39678 454170 39774 454226
rect 39154 454102 39774 454170
rect 39154 454046 39250 454102
rect 39306 454046 39374 454102
rect 39430 454046 39498 454102
rect 39554 454046 39622 454102
rect 39678 454046 39774 454102
rect 39154 453978 39774 454046
rect 39154 453922 39250 453978
rect 39306 453922 39374 453978
rect 39430 453922 39498 453978
rect 39554 453922 39622 453978
rect 39678 453922 39774 453978
rect 39154 436350 39774 453922
rect 39154 436294 39250 436350
rect 39306 436294 39374 436350
rect 39430 436294 39498 436350
rect 39554 436294 39622 436350
rect 39678 436294 39774 436350
rect 39154 436226 39774 436294
rect 39154 436170 39250 436226
rect 39306 436170 39374 436226
rect 39430 436170 39498 436226
rect 39554 436170 39622 436226
rect 39678 436170 39774 436226
rect 39154 436102 39774 436170
rect 39154 436046 39250 436102
rect 39306 436046 39374 436102
rect 39430 436046 39498 436102
rect 39554 436046 39622 436102
rect 39678 436046 39774 436102
rect 39154 435978 39774 436046
rect 39154 435922 39250 435978
rect 39306 435922 39374 435978
rect 39430 435922 39498 435978
rect 39554 435922 39622 435978
rect 39678 435922 39774 435978
rect 39154 418350 39774 435922
rect 39154 418294 39250 418350
rect 39306 418294 39374 418350
rect 39430 418294 39498 418350
rect 39554 418294 39622 418350
rect 39678 418294 39774 418350
rect 39154 418226 39774 418294
rect 39154 418170 39250 418226
rect 39306 418170 39374 418226
rect 39430 418170 39498 418226
rect 39554 418170 39622 418226
rect 39678 418170 39774 418226
rect 39154 418102 39774 418170
rect 39154 418046 39250 418102
rect 39306 418046 39374 418102
rect 39430 418046 39498 418102
rect 39554 418046 39622 418102
rect 39678 418046 39774 418102
rect 39154 417978 39774 418046
rect 39154 417922 39250 417978
rect 39306 417922 39374 417978
rect 39430 417922 39498 417978
rect 39554 417922 39622 417978
rect 39678 417922 39774 417978
rect 39154 400350 39774 417922
rect 39154 400294 39250 400350
rect 39306 400294 39374 400350
rect 39430 400294 39498 400350
rect 39554 400294 39622 400350
rect 39678 400294 39774 400350
rect 39154 400226 39774 400294
rect 39154 400170 39250 400226
rect 39306 400170 39374 400226
rect 39430 400170 39498 400226
rect 39554 400170 39622 400226
rect 39678 400170 39774 400226
rect 39154 400102 39774 400170
rect 39154 400046 39250 400102
rect 39306 400046 39374 400102
rect 39430 400046 39498 400102
rect 39554 400046 39622 400102
rect 39678 400046 39774 400102
rect 39154 399978 39774 400046
rect 39154 399922 39250 399978
rect 39306 399922 39374 399978
rect 39430 399922 39498 399978
rect 39554 399922 39622 399978
rect 39678 399922 39774 399978
rect 39154 382350 39774 399922
rect 39154 382294 39250 382350
rect 39306 382294 39374 382350
rect 39430 382294 39498 382350
rect 39554 382294 39622 382350
rect 39678 382294 39774 382350
rect 39154 382226 39774 382294
rect 39154 382170 39250 382226
rect 39306 382170 39374 382226
rect 39430 382170 39498 382226
rect 39554 382170 39622 382226
rect 39678 382170 39774 382226
rect 39154 382102 39774 382170
rect 39154 382046 39250 382102
rect 39306 382046 39374 382102
rect 39430 382046 39498 382102
rect 39554 382046 39622 382102
rect 39678 382046 39774 382102
rect 39154 381978 39774 382046
rect 39154 381922 39250 381978
rect 39306 381922 39374 381978
rect 39430 381922 39498 381978
rect 39554 381922 39622 381978
rect 39678 381922 39774 381978
rect 39154 364350 39774 381922
rect 39154 364294 39250 364350
rect 39306 364294 39374 364350
rect 39430 364294 39498 364350
rect 39554 364294 39622 364350
rect 39678 364294 39774 364350
rect 39154 364226 39774 364294
rect 39154 364170 39250 364226
rect 39306 364170 39374 364226
rect 39430 364170 39498 364226
rect 39554 364170 39622 364226
rect 39678 364170 39774 364226
rect 39154 364102 39774 364170
rect 39154 364046 39250 364102
rect 39306 364046 39374 364102
rect 39430 364046 39498 364102
rect 39554 364046 39622 364102
rect 39678 364046 39774 364102
rect 39154 363978 39774 364046
rect 39154 363922 39250 363978
rect 39306 363922 39374 363978
rect 39430 363922 39498 363978
rect 39554 363922 39622 363978
rect 39678 363922 39774 363978
rect 37772 190866 37828 190876
rect 37884 361396 37940 361406
rect 37884 131908 37940 361340
rect 37884 131842 37940 131852
rect 39154 346350 39774 363922
rect 39154 346294 39250 346350
rect 39306 346294 39374 346350
rect 39430 346294 39498 346350
rect 39554 346294 39622 346350
rect 39678 346294 39774 346350
rect 39154 346226 39774 346294
rect 39154 346170 39250 346226
rect 39306 346170 39374 346226
rect 39430 346170 39498 346226
rect 39554 346170 39622 346226
rect 39678 346170 39774 346226
rect 39154 346102 39774 346170
rect 39154 346046 39250 346102
rect 39306 346046 39374 346102
rect 39430 346046 39498 346102
rect 39554 346046 39622 346102
rect 39678 346046 39774 346102
rect 39154 345978 39774 346046
rect 39154 345922 39250 345978
rect 39306 345922 39374 345978
rect 39430 345922 39498 345978
rect 39554 345922 39622 345978
rect 39678 345922 39774 345978
rect 39154 328350 39774 345922
rect 39154 328294 39250 328350
rect 39306 328294 39374 328350
rect 39430 328294 39498 328350
rect 39554 328294 39622 328350
rect 39678 328294 39774 328350
rect 39154 328226 39774 328294
rect 39154 328170 39250 328226
rect 39306 328170 39374 328226
rect 39430 328170 39498 328226
rect 39554 328170 39622 328226
rect 39678 328170 39774 328226
rect 39154 328102 39774 328170
rect 39154 328046 39250 328102
rect 39306 328046 39374 328102
rect 39430 328046 39498 328102
rect 39554 328046 39622 328102
rect 39678 328046 39774 328102
rect 39154 327978 39774 328046
rect 39154 327922 39250 327978
rect 39306 327922 39374 327978
rect 39430 327922 39498 327978
rect 39554 327922 39622 327978
rect 39678 327922 39774 327978
rect 39154 310350 39774 327922
rect 39154 310294 39250 310350
rect 39306 310294 39374 310350
rect 39430 310294 39498 310350
rect 39554 310294 39622 310350
rect 39678 310294 39774 310350
rect 39154 310226 39774 310294
rect 39154 310170 39250 310226
rect 39306 310170 39374 310226
rect 39430 310170 39498 310226
rect 39554 310170 39622 310226
rect 39678 310170 39774 310226
rect 39154 310102 39774 310170
rect 39154 310046 39250 310102
rect 39306 310046 39374 310102
rect 39430 310046 39498 310102
rect 39554 310046 39622 310102
rect 39678 310046 39774 310102
rect 39154 309978 39774 310046
rect 39154 309922 39250 309978
rect 39306 309922 39374 309978
rect 39430 309922 39498 309978
rect 39554 309922 39622 309978
rect 39678 309922 39774 309978
rect 39154 292350 39774 309922
rect 39154 292294 39250 292350
rect 39306 292294 39374 292350
rect 39430 292294 39498 292350
rect 39554 292294 39622 292350
rect 39678 292294 39774 292350
rect 39154 292226 39774 292294
rect 39154 292170 39250 292226
rect 39306 292170 39374 292226
rect 39430 292170 39498 292226
rect 39554 292170 39622 292226
rect 39678 292170 39774 292226
rect 39154 292102 39774 292170
rect 39154 292046 39250 292102
rect 39306 292046 39374 292102
rect 39430 292046 39498 292102
rect 39554 292046 39622 292102
rect 39678 292046 39774 292102
rect 39154 291978 39774 292046
rect 39154 291922 39250 291978
rect 39306 291922 39374 291978
rect 39430 291922 39498 291978
rect 39554 291922 39622 291978
rect 39678 291922 39774 291978
rect 39154 274350 39774 291922
rect 39154 274294 39250 274350
rect 39306 274294 39374 274350
rect 39430 274294 39498 274350
rect 39554 274294 39622 274350
rect 39678 274294 39774 274350
rect 39154 274226 39774 274294
rect 39154 274170 39250 274226
rect 39306 274170 39374 274226
rect 39430 274170 39498 274226
rect 39554 274170 39622 274226
rect 39678 274170 39774 274226
rect 39154 274102 39774 274170
rect 39154 274046 39250 274102
rect 39306 274046 39374 274102
rect 39430 274046 39498 274102
rect 39554 274046 39622 274102
rect 39678 274046 39774 274102
rect 39154 273978 39774 274046
rect 39154 273922 39250 273978
rect 39306 273922 39374 273978
rect 39430 273922 39498 273978
rect 39554 273922 39622 273978
rect 39678 273922 39774 273978
rect 39154 256350 39774 273922
rect 39154 256294 39250 256350
rect 39306 256294 39374 256350
rect 39430 256294 39498 256350
rect 39554 256294 39622 256350
rect 39678 256294 39774 256350
rect 39154 256226 39774 256294
rect 39154 256170 39250 256226
rect 39306 256170 39374 256226
rect 39430 256170 39498 256226
rect 39554 256170 39622 256226
rect 39678 256170 39774 256226
rect 39154 256102 39774 256170
rect 39154 256046 39250 256102
rect 39306 256046 39374 256102
rect 39430 256046 39498 256102
rect 39554 256046 39622 256102
rect 39678 256046 39774 256102
rect 39154 255978 39774 256046
rect 39154 255922 39250 255978
rect 39306 255922 39374 255978
rect 39430 255922 39498 255978
rect 39554 255922 39622 255978
rect 39678 255922 39774 255978
rect 39154 238350 39774 255922
rect 39154 238294 39250 238350
rect 39306 238294 39374 238350
rect 39430 238294 39498 238350
rect 39554 238294 39622 238350
rect 39678 238294 39774 238350
rect 39154 238226 39774 238294
rect 39154 238170 39250 238226
rect 39306 238170 39374 238226
rect 39430 238170 39498 238226
rect 39554 238170 39622 238226
rect 39678 238170 39774 238226
rect 39154 238102 39774 238170
rect 39154 238046 39250 238102
rect 39306 238046 39374 238102
rect 39430 238046 39498 238102
rect 39554 238046 39622 238102
rect 39678 238046 39774 238102
rect 39154 237978 39774 238046
rect 39154 237922 39250 237978
rect 39306 237922 39374 237978
rect 39430 237922 39498 237978
rect 39554 237922 39622 237978
rect 39678 237922 39774 237978
rect 39154 220350 39774 237922
rect 39154 220294 39250 220350
rect 39306 220294 39374 220350
rect 39430 220294 39498 220350
rect 39554 220294 39622 220350
rect 39678 220294 39774 220350
rect 39154 220226 39774 220294
rect 39154 220170 39250 220226
rect 39306 220170 39374 220226
rect 39430 220170 39498 220226
rect 39554 220170 39622 220226
rect 39678 220170 39774 220226
rect 39154 220102 39774 220170
rect 39154 220046 39250 220102
rect 39306 220046 39374 220102
rect 39430 220046 39498 220102
rect 39554 220046 39622 220102
rect 39678 220046 39774 220102
rect 39154 219978 39774 220046
rect 39154 219922 39250 219978
rect 39306 219922 39374 219978
rect 39430 219922 39498 219978
rect 39554 219922 39622 219978
rect 39678 219922 39774 219978
rect 39154 202350 39774 219922
rect 39154 202294 39250 202350
rect 39306 202294 39374 202350
rect 39430 202294 39498 202350
rect 39554 202294 39622 202350
rect 39678 202294 39774 202350
rect 39154 202226 39774 202294
rect 39154 202170 39250 202226
rect 39306 202170 39374 202226
rect 39430 202170 39498 202226
rect 39554 202170 39622 202226
rect 39678 202170 39774 202226
rect 39154 202102 39774 202170
rect 39154 202046 39250 202102
rect 39306 202046 39374 202102
rect 39430 202046 39498 202102
rect 39554 202046 39622 202102
rect 39678 202046 39774 202102
rect 39154 201978 39774 202046
rect 39154 201922 39250 201978
rect 39306 201922 39374 201978
rect 39430 201922 39498 201978
rect 39554 201922 39622 201978
rect 39678 201922 39774 201978
rect 39154 184350 39774 201922
rect 42874 598172 43494 598268
rect 42874 598116 42970 598172
rect 43026 598116 43094 598172
rect 43150 598116 43218 598172
rect 43274 598116 43342 598172
rect 43398 598116 43494 598172
rect 42874 598048 43494 598116
rect 42874 597992 42970 598048
rect 43026 597992 43094 598048
rect 43150 597992 43218 598048
rect 43274 597992 43342 598048
rect 43398 597992 43494 598048
rect 42874 597924 43494 597992
rect 42874 597868 42970 597924
rect 43026 597868 43094 597924
rect 43150 597868 43218 597924
rect 43274 597868 43342 597924
rect 43398 597868 43494 597924
rect 42874 597800 43494 597868
rect 42874 597744 42970 597800
rect 43026 597744 43094 597800
rect 43150 597744 43218 597800
rect 43274 597744 43342 597800
rect 43398 597744 43494 597800
rect 42874 586350 43494 597744
rect 42874 586294 42970 586350
rect 43026 586294 43094 586350
rect 43150 586294 43218 586350
rect 43274 586294 43342 586350
rect 43398 586294 43494 586350
rect 42874 586226 43494 586294
rect 42874 586170 42970 586226
rect 43026 586170 43094 586226
rect 43150 586170 43218 586226
rect 43274 586170 43342 586226
rect 43398 586170 43494 586226
rect 42874 586102 43494 586170
rect 42874 586046 42970 586102
rect 43026 586046 43094 586102
rect 43150 586046 43218 586102
rect 43274 586046 43342 586102
rect 43398 586046 43494 586102
rect 42874 585978 43494 586046
rect 42874 585922 42970 585978
rect 43026 585922 43094 585978
rect 43150 585922 43218 585978
rect 43274 585922 43342 585978
rect 43398 585922 43494 585978
rect 42874 568350 43494 585922
rect 42874 568294 42970 568350
rect 43026 568294 43094 568350
rect 43150 568294 43218 568350
rect 43274 568294 43342 568350
rect 43398 568294 43494 568350
rect 42874 568226 43494 568294
rect 42874 568170 42970 568226
rect 43026 568170 43094 568226
rect 43150 568170 43218 568226
rect 43274 568170 43342 568226
rect 43398 568170 43494 568226
rect 42874 568102 43494 568170
rect 42874 568046 42970 568102
rect 43026 568046 43094 568102
rect 43150 568046 43218 568102
rect 43274 568046 43342 568102
rect 43398 568046 43494 568102
rect 42874 567978 43494 568046
rect 42874 567922 42970 567978
rect 43026 567922 43094 567978
rect 43150 567922 43218 567978
rect 43274 567922 43342 567978
rect 43398 567922 43494 567978
rect 42874 550350 43494 567922
rect 42874 550294 42970 550350
rect 43026 550294 43094 550350
rect 43150 550294 43218 550350
rect 43274 550294 43342 550350
rect 43398 550294 43494 550350
rect 42874 550226 43494 550294
rect 42874 550170 42970 550226
rect 43026 550170 43094 550226
rect 43150 550170 43218 550226
rect 43274 550170 43342 550226
rect 43398 550170 43494 550226
rect 42874 550102 43494 550170
rect 42874 550046 42970 550102
rect 43026 550046 43094 550102
rect 43150 550046 43218 550102
rect 43274 550046 43342 550102
rect 43398 550046 43494 550102
rect 42874 549978 43494 550046
rect 42874 549922 42970 549978
rect 43026 549922 43094 549978
rect 43150 549922 43218 549978
rect 43274 549922 43342 549978
rect 43398 549922 43494 549978
rect 42874 532350 43494 549922
rect 42874 532294 42970 532350
rect 43026 532294 43094 532350
rect 43150 532294 43218 532350
rect 43274 532294 43342 532350
rect 43398 532294 43494 532350
rect 42874 532226 43494 532294
rect 42874 532170 42970 532226
rect 43026 532170 43094 532226
rect 43150 532170 43218 532226
rect 43274 532170 43342 532226
rect 43398 532170 43494 532226
rect 42874 532102 43494 532170
rect 42874 532046 42970 532102
rect 43026 532046 43094 532102
rect 43150 532046 43218 532102
rect 43274 532046 43342 532102
rect 43398 532046 43494 532102
rect 42874 531978 43494 532046
rect 42874 531922 42970 531978
rect 43026 531922 43094 531978
rect 43150 531922 43218 531978
rect 43274 531922 43342 531978
rect 43398 531922 43494 531978
rect 42874 514350 43494 531922
rect 42874 514294 42970 514350
rect 43026 514294 43094 514350
rect 43150 514294 43218 514350
rect 43274 514294 43342 514350
rect 43398 514294 43494 514350
rect 42874 514226 43494 514294
rect 42874 514170 42970 514226
rect 43026 514170 43094 514226
rect 43150 514170 43218 514226
rect 43274 514170 43342 514226
rect 43398 514170 43494 514226
rect 42874 514102 43494 514170
rect 42874 514046 42970 514102
rect 43026 514046 43094 514102
rect 43150 514046 43218 514102
rect 43274 514046 43342 514102
rect 43398 514046 43494 514102
rect 42874 513978 43494 514046
rect 42874 513922 42970 513978
rect 43026 513922 43094 513978
rect 43150 513922 43218 513978
rect 43274 513922 43342 513978
rect 43398 513922 43494 513978
rect 42874 496350 43494 513922
rect 42874 496294 42970 496350
rect 43026 496294 43094 496350
rect 43150 496294 43218 496350
rect 43274 496294 43342 496350
rect 43398 496294 43494 496350
rect 42874 496226 43494 496294
rect 42874 496170 42970 496226
rect 43026 496170 43094 496226
rect 43150 496170 43218 496226
rect 43274 496170 43342 496226
rect 43398 496170 43494 496226
rect 42874 496102 43494 496170
rect 42874 496046 42970 496102
rect 43026 496046 43094 496102
rect 43150 496046 43218 496102
rect 43274 496046 43342 496102
rect 43398 496046 43494 496102
rect 42874 495978 43494 496046
rect 42874 495922 42970 495978
rect 43026 495922 43094 495978
rect 43150 495922 43218 495978
rect 43274 495922 43342 495978
rect 43398 495922 43494 495978
rect 42874 478350 43494 495922
rect 42874 478294 42970 478350
rect 43026 478294 43094 478350
rect 43150 478294 43218 478350
rect 43274 478294 43342 478350
rect 43398 478294 43494 478350
rect 42874 478226 43494 478294
rect 42874 478170 42970 478226
rect 43026 478170 43094 478226
rect 43150 478170 43218 478226
rect 43274 478170 43342 478226
rect 43398 478170 43494 478226
rect 42874 478102 43494 478170
rect 42874 478046 42970 478102
rect 43026 478046 43094 478102
rect 43150 478046 43218 478102
rect 43274 478046 43342 478102
rect 43398 478046 43494 478102
rect 42874 477978 43494 478046
rect 42874 477922 42970 477978
rect 43026 477922 43094 477978
rect 43150 477922 43218 477978
rect 43274 477922 43342 477978
rect 43398 477922 43494 477978
rect 42874 460350 43494 477922
rect 42874 460294 42970 460350
rect 43026 460294 43094 460350
rect 43150 460294 43218 460350
rect 43274 460294 43342 460350
rect 43398 460294 43494 460350
rect 42874 460226 43494 460294
rect 42874 460170 42970 460226
rect 43026 460170 43094 460226
rect 43150 460170 43218 460226
rect 43274 460170 43342 460226
rect 43398 460170 43494 460226
rect 42874 460102 43494 460170
rect 42874 460046 42970 460102
rect 43026 460046 43094 460102
rect 43150 460046 43218 460102
rect 43274 460046 43342 460102
rect 43398 460046 43494 460102
rect 42874 459978 43494 460046
rect 42874 459922 42970 459978
rect 43026 459922 43094 459978
rect 43150 459922 43218 459978
rect 43274 459922 43342 459978
rect 43398 459922 43494 459978
rect 42874 442350 43494 459922
rect 42874 442294 42970 442350
rect 43026 442294 43094 442350
rect 43150 442294 43218 442350
rect 43274 442294 43342 442350
rect 43398 442294 43494 442350
rect 42874 442226 43494 442294
rect 42874 442170 42970 442226
rect 43026 442170 43094 442226
rect 43150 442170 43218 442226
rect 43274 442170 43342 442226
rect 43398 442170 43494 442226
rect 42874 442102 43494 442170
rect 42874 442046 42970 442102
rect 43026 442046 43094 442102
rect 43150 442046 43218 442102
rect 43274 442046 43342 442102
rect 43398 442046 43494 442102
rect 42874 441978 43494 442046
rect 42874 441922 42970 441978
rect 43026 441922 43094 441978
rect 43150 441922 43218 441978
rect 43274 441922 43342 441978
rect 43398 441922 43494 441978
rect 42874 424350 43494 441922
rect 42874 424294 42970 424350
rect 43026 424294 43094 424350
rect 43150 424294 43218 424350
rect 43274 424294 43342 424350
rect 43398 424294 43494 424350
rect 42874 424226 43494 424294
rect 42874 424170 42970 424226
rect 43026 424170 43094 424226
rect 43150 424170 43218 424226
rect 43274 424170 43342 424226
rect 43398 424170 43494 424226
rect 42874 424102 43494 424170
rect 42874 424046 42970 424102
rect 43026 424046 43094 424102
rect 43150 424046 43218 424102
rect 43274 424046 43342 424102
rect 43398 424046 43494 424102
rect 42874 423978 43494 424046
rect 42874 423922 42970 423978
rect 43026 423922 43094 423978
rect 43150 423922 43218 423978
rect 43274 423922 43342 423978
rect 43398 423922 43494 423978
rect 42874 406350 43494 423922
rect 42874 406294 42970 406350
rect 43026 406294 43094 406350
rect 43150 406294 43218 406350
rect 43274 406294 43342 406350
rect 43398 406294 43494 406350
rect 42874 406226 43494 406294
rect 42874 406170 42970 406226
rect 43026 406170 43094 406226
rect 43150 406170 43218 406226
rect 43274 406170 43342 406226
rect 43398 406170 43494 406226
rect 42874 406102 43494 406170
rect 42874 406046 42970 406102
rect 43026 406046 43094 406102
rect 43150 406046 43218 406102
rect 43274 406046 43342 406102
rect 43398 406046 43494 406102
rect 42874 405978 43494 406046
rect 42874 405922 42970 405978
rect 43026 405922 43094 405978
rect 43150 405922 43218 405978
rect 43274 405922 43342 405978
rect 43398 405922 43494 405978
rect 42874 388350 43494 405922
rect 42874 388294 42970 388350
rect 43026 388294 43094 388350
rect 43150 388294 43218 388350
rect 43274 388294 43342 388350
rect 43398 388294 43494 388350
rect 42874 388226 43494 388294
rect 42874 388170 42970 388226
rect 43026 388170 43094 388226
rect 43150 388170 43218 388226
rect 43274 388170 43342 388226
rect 43398 388170 43494 388226
rect 42874 388102 43494 388170
rect 42874 388046 42970 388102
rect 43026 388046 43094 388102
rect 43150 388046 43218 388102
rect 43274 388046 43342 388102
rect 43398 388046 43494 388102
rect 42874 387978 43494 388046
rect 42874 387922 42970 387978
rect 43026 387922 43094 387978
rect 43150 387922 43218 387978
rect 43274 387922 43342 387978
rect 43398 387922 43494 387978
rect 42874 370350 43494 387922
rect 42874 370294 42970 370350
rect 43026 370294 43094 370350
rect 43150 370294 43218 370350
rect 43274 370294 43342 370350
rect 43398 370294 43494 370350
rect 42874 370226 43494 370294
rect 42874 370170 42970 370226
rect 43026 370170 43094 370226
rect 43150 370170 43218 370226
rect 43274 370170 43342 370226
rect 43398 370170 43494 370226
rect 42874 370102 43494 370170
rect 42874 370046 42970 370102
rect 43026 370046 43094 370102
rect 43150 370046 43218 370102
rect 43274 370046 43342 370102
rect 43398 370046 43494 370102
rect 42874 369978 43494 370046
rect 42874 369922 42970 369978
rect 43026 369922 43094 369978
rect 43150 369922 43218 369978
rect 43274 369922 43342 369978
rect 43398 369922 43494 369978
rect 42874 352350 43494 369922
rect 42874 352294 42970 352350
rect 43026 352294 43094 352350
rect 43150 352294 43218 352350
rect 43274 352294 43342 352350
rect 43398 352294 43494 352350
rect 42874 352226 43494 352294
rect 42874 352170 42970 352226
rect 43026 352170 43094 352226
rect 43150 352170 43218 352226
rect 43274 352170 43342 352226
rect 43398 352170 43494 352226
rect 42874 352102 43494 352170
rect 42874 352046 42970 352102
rect 43026 352046 43094 352102
rect 43150 352046 43218 352102
rect 43274 352046 43342 352102
rect 43398 352046 43494 352102
rect 42874 351978 43494 352046
rect 42874 351922 42970 351978
rect 43026 351922 43094 351978
rect 43150 351922 43218 351978
rect 43274 351922 43342 351978
rect 43398 351922 43494 351978
rect 42874 334350 43494 351922
rect 42874 334294 42970 334350
rect 43026 334294 43094 334350
rect 43150 334294 43218 334350
rect 43274 334294 43342 334350
rect 43398 334294 43494 334350
rect 42874 334226 43494 334294
rect 42874 334170 42970 334226
rect 43026 334170 43094 334226
rect 43150 334170 43218 334226
rect 43274 334170 43342 334226
rect 43398 334170 43494 334226
rect 42874 334102 43494 334170
rect 42874 334046 42970 334102
rect 43026 334046 43094 334102
rect 43150 334046 43218 334102
rect 43274 334046 43342 334102
rect 43398 334046 43494 334102
rect 42874 333978 43494 334046
rect 42874 333922 42970 333978
rect 43026 333922 43094 333978
rect 43150 333922 43218 333978
rect 43274 333922 43342 333978
rect 43398 333922 43494 333978
rect 42874 316350 43494 333922
rect 42874 316294 42970 316350
rect 43026 316294 43094 316350
rect 43150 316294 43218 316350
rect 43274 316294 43342 316350
rect 43398 316294 43494 316350
rect 42874 316226 43494 316294
rect 42874 316170 42970 316226
rect 43026 316170 43094 316226
rect 43150 316170 43218 316226
rect 43274 316170 43342 316226
rect 43398 316170 43494 316226
rect 42874 316102 43494 316170
rect 42874 316046 42970 316102
rect 43026 316046 43094 316102
rect 43150 316046 43218 316102
rect 43274 316046 43342 316102
rect 43398 316046 43494 316102
rect 42874 315978 43494 316046
rect 42874 315922 42970 315978
rect 43026 315922 43094 315978
rect 43150 315922 43218 315978
rect 43274 315922 43342 315978
rect 43398 315922 43494 315978
rect 42874 298350 43494 315922
rect 42874 298294 42970 298350
rect 43026 298294 43094 298350
rect 43150 298294 43218 298350
rect 43274 298294 43342 298350
rect 43398 298294 43494 298350
rect 42874 298226 43494 298294
rect 42874 298170 42970 298226
rect 43026 298170 43094 298226
rect 43150 298170 43218 298226
rect 43274 298170 43342 298226
rect 43398 298170 43494 298226
rect 42874 298102 43494 298170
rect 42874 298046 42970 298102
rect 43026 298046 43094 298102
rect 43150 298046 43218 298102
rect 43274 298046 43342 298102
rect 43398 298046 43494 298102
rect 42874 297978 43494 298046
rect 42874 297922 42970 297978
rect 43026 297922 43094 297978
rect 43150 297922 43218 297978
rect 43274 297922 43342 297978
rect 43398 297922 43494 297978
rect 42874 280350 43494 297922
rect 42874 280294 42970 280350
rect 43026 280294 43094 280350
rect 43150 280294 43218 280350
rect 43274 280294 43342 280350
rect 43398 280294 43494 280350
rect 42874 280226 43494 280294
rect 42874 280170 42970 280226
rect 43026 280170 43094 280226
rect 43150 280170 43218 280226
rect 43274 280170 43342 280226
rect 43398 280170 43494 280226
rect 42874 280102 43494 280170
rect 42874 280046 42970 280102
rect 43026 280046 43094 280102
rect 43150 280046 43218 280102
rect 43274 280046 43342 280102
rect 43398 280046 43494 280102
rect 42874 279978 43494 280046
rect 42874 279922 42970 279978
rect 43026 279922 43094 279978
rect 43150 279922 43218 279978
rect 43274 279922 43342 279978
rect 43398 279922 43494 279978
rect 42874 262350 43494 279922
rect 42874 262294 42970 262350
rect 43026 262294 43094 262350
rect 43150 262294 43218 262350
rect 43274 262294 43342 262350
rect 43398 262294 43494 262350
rect 42874 262226 43494 262294
rect 42874 262170 42970 262226
rect 43026 262170 43094 262226
rect 43150 262170 43218 262226
rect 43274 262170 43342 262226
rect 43398 262170 43494 262226
rect 42874 262102 43494 262170
rect 42874 262046 42970 262102
rect 43026 262046 43094 262102
rect 43150 262046 43218 262102
rect 43274 262046 43342 262102
rect 43398 262046 43494 262102
rect 42874 261978 43494 262046
rect 42874 261922 42970 261978
rect 43026 261922 43094 261978
rect 43150 261922 43218 261978
rect 43274 261922 43342 261978
rect 43398 261922 43494 261978
rect 42874 244350 43494 261922
rect 42874 244294 42970 244350
rect 43026 244294 43094 244350
rect 43150 244294 43218 244350
rect 43274 244294 43342 244350
rect 43398 244294 43494 244350
rect 42874 244226 43494 244294
rect 42874 244170 42970 244226
rect 43026 244170 43094 244226
rect 43150 244170 43218 244226
rect 43274 244170 43342 244226
rect 43398 244170 43494 244226
rect 42874 244102 43494 244170
rect 42874 244046 42970 244102
rect 43026 244046 43094 244102
rect 43150 244046 43218 244102
rect 43274 244046 43342 244102
rect 43398 244046 43494 244102
rect 42874 243978 43494 244046
rect 42874 243922 42970 243978
rect 43026 243922 43094 243978
rect 43150 243922 43218 243978
rect 43274 243922 43342 243978
rect 43398 243922 43494 243978
rect 42874 226350 43494 243922
rect 57154 597212 57774 598268
rect 57154 597156 57250 597212
rect 57306 597156 57374 597212
rect 57430 597156 57498 597212
rect 57554 597156 57622 597212
rect 57678 597156 57774 597212
rect 57154 597088 57774 597156
rect 57154 597032 57250 597088
rect 57306 597032 57374 597088
rect 57430 597032 57498 597088
rect 57554 597032 57622 597088
rect 57678 597032 57774 597088
rect 57154 596964 57774 597032
rect 57154 596908 57250 596964
rect 57306 596908 57374 596964
rect 57430 596908 57498 596964
rect 57554 596908 57622 596964
rect 57678 596908 57774 596964
rect 57154 596840 57774 596908
rect 57154 596784 57250 596840
rect 57306 596784 57374 596840
rect 57430 596784 57498 596840
rect 57554 596784 57622 596840
rect 57678 596784 57774 596840
rect 57154 580350 57774 596784
rect 57154 580294 57250 580350
rect 57306 580294 57374 580350
rect 57430 580294 57498 580350
rect 57554 580294 57622 580350
rect 57678 580294 57774 580350
rect 57154 580226 57774 580294
rect 57154 580170 57250 580226
rect 57306 580170 57374 580226
rect 57430 580170 57498 580226
rect 57554 580170 57622 580226
rect 57678 580170 57774 580226
rect 57154 580102 57774 580170
rect 57154 580046 57250 580102
rect 57306 580046 57374 580102
rect 57430 580046 57498 580102
rect 57554 580046 57622 580102
rect 57678 580046 57774 580102
rect 57154 579978 57774 580046
rect 57154 579922 57250 579978
rect 57306 579922 57374 579978
rect 57430 579922 57498 579978
rect 57554 579922 57622 579978
rect 57678 579922 57774 579978
rect 57154 562350 57774 579922
rect 57154 562294 57250 562350
rect 57306 562294 57374 562350
rect 57430 562294 57498 562350
rect 57554 562294 57622 562350
rect 57678 562294 57774 562350
rect 57154 562226 57774 562294
rect 57154 562170 57250 562226
rect 57306 562170 57374 562226
rect 57430 562170 57498 562226
rect 57554 562170 57622 562226
rect 57678 562170 57774 562226
rect 57154 562102 57774 562170
rect 57154 562046 57250 562102
rect 57306 562046 57374 562102
rect 57430 562046 57498 562102
rect 57554 562046 57622 562102
rect 57678 562046 57774 562102
rect 57154 561978 57774 562046
rect 57154 561922 57250 561978
rect 57306 561922 57374 561978
rect 57430 561922 57498 561978
rect 57554 561922 57622 561978
rect 57678 561922 57774 561978
rect 57154 544350 57774 561922
rect 57154 544294 57250 544350
rect 57306 544294 57374 544350
rect 57430 544294 57498 544350
rect 57554 544294 57622 544350
rect 57678 544294 57774 544350
rect 57154 544226 57774 544294
rect 57154 544170 57250 544226
rect 57306 544170 57374 544226
rect 57430 544170 57498 544226
rect 57554 544170 57622 544226
rect 57678 544170 57774 544226
rect 57154 544102 57774 544170
rect 57154 544046 57250 544102
rect 57306 544046 57374 544102
rect 57430 544046 57498 544102
rect 57554 544046 57622 544102
rect 57678 544046 57774 544102
rect 57154 543978 57774 544046
rect 57154 543922 57250 543978
rect 57306 543922 57374 543978
rect 57430 543922 57498 543978
rect 57554 543922 57622 543978
rect 57678 543922 57774 543978
rect 57154 526350 57774 543922
rect 57154 526294 57250 526350
rect 57306 526294 57374 526350
rect 57430 526294 57498 526350
rect 57554 526294 57622 526350
rect 57678 526294 57774 526350
rect 57154 526226 57774 526294
rect 57154 526170 57250 526226
rect 57306 526170 57374 526226
rect 57430 526170 57498 526226
rect 57554 526170 57622 526226
rect 57678 526170 57774 526226
rect 57154 526102 57774 526170
rect 57154 526046 57250 526102
rect 57306 526046 57374 526102
rect 57430 526046 57498 526102
rect 57554 526046 57622 526102
rect 57678 526046 57774 526102
rect 57154 525978 57774 526046
rect 57154 525922 57250 525978
rect 57306 525922 57374 525978
rect 57430 525922 57498 525978
rect 57554 525922 57622 525978
rect 57678 525922 57774 525978
rect 57154 508350 57774 525922
rect 57154 508294 57250 508350
rect 57306 508294 57374 508350
rect 57430 508294 57498 508350
rect 57554 508294 57622 508350
rect 57678 508294 57774 508350
rect 57154 508226 57774 508294
rect 57154 508170 57250 508226
rect 57306 508170 57374 508226
rect 57430 508170 57498 508226
rect 57554 508170 57622 508226
rect 57678 508170 57774 508226
rect 57154 508102 57774 508170
rect 57154 508046 57250 508102
rect 57306 508046 57374 508102
rect 57430 508046 57498 508102
rect 57554 508046 57622 508102
rect 57678 508046 57774 508102
rect 57154 507978 57774 508046
rect 57154 507922 57250 507978
rect 57306 507922 57374 507978
rect 57430 507922 57498 507978
rect 57554 507922 57622 507978
rect 57678 507922 57774 507978
rect 57154 490350 57774 507922
rect 57154 490294 57250 490350
rect 57306 490294 57374 490350
rect 57430 490294 57498 490350
rect 57554 490294 57622 490350
rect 57678 490294 57774 490350
rect 57154 490226 57774 490294
rect 57154 490170 57250 490226
rect 57306 490170 57374 490226
rect 57430 490170 57498 490226
rect 57554 490170 57622 490226
rect 57678 490170 57774 490226
rect 57154 490102 57774 490170
rect 57154 490046 57250 490102
rect 57306 490046 57374 490102
rect 57430 490046 57498 490102
rect 57554 490046 57622 490102
rect 57678 490046 57774 490102
rect 57154 489978 57774 490046
rect 57154 489922 57250 489978
rect 57306 489922 57374 489978
rect 57430 489922 57498 489978
rect 57554 489922 57622 489978
rect 57678 489922 57774 489978
rect 57154 472350 57774 489922
rect 57154 472294 57250 472350
rect 57306 472294 57374 472350
rect 57430 472294 57498 472350
rect 57554 472294 57622 472350
rect 57678 472294 57774 472350
rect 57154 472226 57774 472294
rect 57154 472170 57250 472226
rect 57306 472170 57374 472226
rect 57430 472170 57498 472226
rect 57554 472170 57622 472226
rect 57678 472170 57774 472226
rect 57154 472102 57774 472170
rect 57154 472046 57250 472102
rect 57306 472046 57374 472102
rect 57430 472046 57498 472102
rect 57554 472046 57622 472102
rect 57678 472046 57774 472102
rect 57154 471978 57774 472046
rect 57154 471922 57250 471978
rect 57306 471922 57374 471978
rect 57430 471922 57498 471978
rect 57554 471922 57622 471978
rect 57678 471922 57774 471978
rect 57154 454350 57774 471922
rect 57154 454294 57250 454350
rect 57306 454294 57374 454350
rect 57430 454294 57498 454350
rect 57554 454294 57622 454350
rect 57678 454294 57774 454350
rect 57154 454226 57774 454294
rect 57154 454170 57250 454226
rect 57306 454170 57374 454226
rect 57430 454170 57498 454226
rect 57554 454170 57622 454226
rect 57678 454170 57774 454226
rect 57154 454102 57774 454170
rect 57154 454046 57250 454102
rect 57306 454046 57374 454102
rect 57430 454046 57498 454102
rect 57554 454046 57622 454102
rect 57678 454046 57774 454102
rect 57154 453978 57774 454046
rect 57154 453922 57250 453978
rect 57306 453922 57374 453978
rect 57430 453922 57498 453978
rect 57554 453922 57622 453978
rect 57678 453922 57774 453978
rect 57154 436350 57774 453922
rect 57154 436294 57250 436350
rect 57306 436294 57374 436350
rect 57430 436294 57498 436350
rect 57554 436294 57622 436350
rect 57678 436294 57774 436350
rect 57154 436226 57774 436294
rect 57154 436170 57250 436226
rect 57306 436170 57374 436226
rect 57430 436170 57498 436226
rect 57554 436170 57622 436226
rect 57678 436170 57774 436226
rect 57154 436102 57774 436170
rect 57154 436046 57250 436102
rect 57306 436046 57374 436102
rect 57430 436046 57498 436102
rect 57554 436046 57622 436102
rect 57678 436046 57774 436102
rect 57154 435978 57774 436046
rect 57154 435922 57250 435978
rect 57306 435922 57374 435978
rect 57430 435922 57498 435978
rect 57554 435922 57622 435978
rect 57678 435922 57774 435978
rect 57154 418350 57774 435922
rect 57154 418294 57250 418350
rect 57306 418294 57374 418350
rect 57430 418294 57498 418350
rect 57554 418294 57622 418350
rect 57678 418294 57774 418350
rect 57154 418226 57774 418294
rect 57154 418170 57250 418226
rect 57306 418170 57374 418226
rect 57430 418170 57498 418226
rect 57554 418170 57622 418226
rect 57678 418170 57774 418226
rect 57154 418102 57774 418170
rect 57154 418046 57250 418102
rect 57306 418046 57374 418102
rect 57430 418046 57498 418102
rect 57554 418046 57622 418102
rect 57678 418046 57774 418102
rect 57154 417978 57774 418046
rect 57154 417922 57250 417978
rect 57306 417922 57374 417978
rect 57430 417922 57498 417978
rect 57554 417922 57622 417978
rect 57678 417922 57774 417978
rect 57154 400350 57774 417922
rect 57154 400294 57250 400350
rect 57306 400294 57374 400350
rect 57430 400294 57498 400350
rect 57554 400294 57622 400350
rect 57678 400294 57774 400350
rect 57154 400226 57774 400294
rect 57154 400170 57250 400226
rect 57306 400170 57374 400226
rect 57430 400170 57498 400226
rect 57554 400170 57622 400226
rect 57678 400170 57774 400226
rect 57154 400102 57774 400170
rect 57154 400046 57250 400102
rect 57306 400046 57374 400102
rect 57430 400046 57498 400102
rect 57554 400046 57622 400102
rect 57678 400046 57774 400102
rect 57154 399978 57774 400046
rect 57154 399922 57250 399978
rect 57306 399922 57374 399978
rect 57430 399922 57498 399978
rect 57554 399922 57622 399978
rect 57678 399922 57774 399978
rect 57154 382350 57774 399922
rect 57154 382294 57250 382350
rect 57306 382294 57374 382350
rect 57430 382294 57498 382350
rect 57554 382294 57622 382350
rect 57678 382294 57774 382350
rect 57154 382226 57774 382294
rect 57154 382170 57250 382226
rect 57306 382170 57374 382226
rect 57430 382170 57498 382226
rect 57554 382170 57622 382226
rect 57678 382170 57774 382226
rect 57154 382102 57774 382170
rect 57154 382046 57250 382102
rect 57306 382046 57374 382102
rect 57430 382046 57498 382102
rect 57554 382046 57622 382102
rect 57678 382046 57774 382102
rect 57154 381978 57774 382046
rect 57154 381922 57250 381978
rect 57306 381922 57374 381978
rect 57430 381922 57498 381978
rect 57554 381922 57622 381978
rect 57678 381922 57774 381978
rect 57154 364350 57774 381922
rect 57154 364294 57250 364350
rect 57306 364294 57374 364350
rect 57430 364294 57498 364350
rect 57554 364294 57622 364350
rect 57678 364294 57774 364350
rect 57154 364226 57774 364294
rect 57154 364170 57250 364226
rect 57306 364170 57374 364226
rect 57430 364170 57498 364226
rect 57554 364170 57622 364226
rect 57678 364170 57774 364226
rect 57154 364102 57774 364170
rect 57154 364046 57250 364102
rect 57306 364046 57374 364102
rect 57430 364046 57498 364102
rect 57554 364046 57622 364102
rect 57678 364046 57774 364102
rect 57154 363978 57774 364046
rect 57154 363922 57250 363978
rect 57306 363922 57374 363978
rect 57430 363922 57498 363978
rect 57554 363922 57622 363978
rect 57678 363922 57774 363978
rect 57154 346350 57774 363922
rect 57154 346294 57250 346350
rect 57306 346294 57374 346350
rect 57430 346294 57498 346350
rect 57554 346294 57622 346350
rect 57678 346294 57774 346350
rect 57154 346226 57774 346294
rect 57154 346170 57250 346226
rect 57306 346170 57374 346226
rect 57430 346170 57498 346226
rect 57554 346170 57622 346226
rect 57678 346170 57774 346226
rect 57154 346102 57774 346170
rect 57154 346046 57250 346102
rect 57306 346046 57374 346102
rect 57430 346046 57498 346102
rect 57554 346046 57622 346102
rect 57678 346046 57774 346102
rect 57154 345978 57774 346046
rect 57154 345922 57250 345978
rect 57306 345922 57374 345978
rect 57430 345922 57498 345978
rect 57554 345922 57622 345978
rect 57678 345922 57774 345978
rect 57154 328350 57774 345922
rect 57154 328294 57250 328350
rect 57306 328294 57374 328350
rect 57430 328294 57498 328350
rect 57554 328294 57622 328350
rect 57678 328294 57774 328350
rect 57154 328226 57774 328294
rect 57154 328170 57250 328226
rect 57306 328170 57374 328226
rect 57430 328170 57498 328226
rect 57554 328170 57622 328226
rect 57678 328170 57774 328226
rect 57154 328102 57774 328170
rect 57154 328046 57250 328102
rect 57306 328046 57374 328102
rect 57430 328046 57498 328102
rect 57554 328046 57622 328102
rect 57678 328046 57774 328102
rect 57154 327978 57774 328046
rect 57154 327922 57250 327978
rect 57306 327922 57374 327978
rect 57430 327922 57498 327978
rect 57554 327922 57622 327978
rect 57678 327922 57774 327978
rect 57154 310350 57774 327922
rect 57154 310294 57250 310350
rect 57306 310294 57374 310350
rect 57430 310294 57498 310350
rect 57554 310294 57622 310350
rect 57678 310294 57774 310350
rect 57154 310226 57774 310294
rect 57154 310170 57250 310226
rect 57306 310170 57374 310226
rect 57430 310170 57498 310226
rect 57554 310170 57622 310226
rect 57678 310170 57774 310226
rect 57154 310102 57774 310170
rect 57154 310046 57250 310102
rect 57306 310046 57374 310102
rect 57430 310046 57498 310102
rect 57554 310046 57622 310102
rect 57678 310046 57774 310102
rect 57154 309978 57774 310046
rect 57154 309922 57250 309978
rect 57306 309922 57374 309978
rect 57430 309922 57498 309978
rect 57554 309922 57622 309978
rect 57678 309922 57774 309978
rect 57154 292350 57774 309922
rect 57154 292294 57250 292350
rect 57306 292294 57374 292350
rect 57430 292294 57498 292350
rect 57554 292294 57622 292350
rect 57678 292294 57774 292350
rect 57154 292226 57774 292294
rect 57154 292170 57250 292226
rect 57306 292170 57374 292226
rect 57430 292170 57498 292226
rect 57554 292170 57622 292226
rect 57678 292170 57774 292226
rect 57154 292102 57774 292170
rect 57154 292046 57250 292102
rect 57306 292046 57374 292102
rect 57430 292046 57498 292102
rect 57554 292046 57622 292102
rect 57678 292046 57774 292102
rect 57154 291978 57774 292046
rect 57154 291922 57250 291978
rect 57306 291922 57374 291978
rect 57430 291922 57498 291978
rect 57554 291922 57622 291978
rect 57678 291922 57774 291978
rect 57154 274350 57774 291922
rect 57154 274294 57250 274350
rect 57306 274294 57374 274350
rect 57430 274294 57498 274350
rect 57554 274294 57622 274350
rect 57678 274294 57774 274350
rect 57154 274226 57774 274294
rect 57154 274170 57250 274226
rect 57306 274170 57374 274226
rect 57430 274170 57498 274226
rect 57554 274170 57622 274226
rect 57678 274170 57774 274226
rect 57154 274102 57774 274170
rect 57154 274046 57250 274102
rect 57306 274046 57374 274102
rect 57430 274046 57498 274102
rect 57554 274046 57622 274102
rect 57678 274046 57774 274102
rect 57154 273978 57774 274046
rect 57154 273922 57250 273978
rect 57306 273922 57374 273978
rect 57430 273922 57498 273978
rect 57554 273922 57622 273978
rect 57678 273922 57774 273978
rect 57154 256350 57774 273922
rect 57154 256294 57250 256350
rect 57306 256294 57374 256350
rect 57430 256294 57498 256350
rect 57554 256294 57622 256350
rect 57678 256294 57774 256350
rect 57154 256226 57774 256294
rect 57154 256170 57250 256226
rect 57306 256170 57374 256226
rect 57430 256170 57498 256226
rect 57554 256170 57622 256226
rect 57678 256170 57774 256226
rect 57154 256102 57774 256170
rect 57154 256046 57250 256102
rect 57306 256046 57374 256102
rect 57430 256046 57498 256102
rect 57554 256046 57622 256102
rect 57678 256046 57774 256102
rect 57154 255978 57774 256046
rect 57154 255922 57250 255978
rect 57306 255922 57374 255978
rect 57430 255922 57498 255978
rect 57554 255922 57622 255978
rect 57678 255922 57774 255978
rect 57154 238350 57774 255922
rect 57154 238294 57250 238350
rect 57306 238294 57374 238350
rect 57430 238294 57498 238350
rect 57554 238294 57622 238350
rect 57678 238294 57774 238350
rect 57154 238226 57774 238294
rect 57154 238170 57250 238226
rect 57306 238170 57374 238226
rect 57430 238170 57498 238226
rect 57554 238170 57622 238226
rect 57678 238170 57774 238226
rect 57154 238102 57774 238170
rect 57154 238046 57250 238102
rect 57306 238046 57374 238102
rect 57430 238046 57498 238102
rect 57554 238046 57622 238102
rect 57678 238046 57774 238102
rect 57154 237978 57774 238046
rect 57154 237922 57250 237978
rect 57306 237922 57374 237978
rect 57430 237922 57498 237978
rect 57554 237922 57622 237978
rect 57678 237922 57774 237978
rect 42874 226294 42970 226350
rect 43026 226294 43094 226350
rect 43150 226294 43218 226350
rect 43274 226294 43342 226350
rect 43398 226294 43494 226350
rect 42874 226226 43494 226294
rect 42874 226170 42970 226226
rect 43026 226170 43094 226226
rect 43150 226170 43218 226226
rect 43274 226170 43342 226226
rect 43398 226170 43494 226226
rect 42874 226102 43494 226170
rect 42874 226046 42970 226102
rect 43026 226046 43094 226102
rect 43150 226046 43218 226102
rect 43274 226046 43342 226102
rect 43398 226046 43494 226102
rect 42874 225978 43494 226046
rect 42874 225922 42970 225978
rect 43026 225922 43094 225978
rect 43150 225922 43218 225978
rect 43274 225922 43342 225978
rect 43398 225922 43494 225978
rect 42874 208350 43494 225922
rect 42874 208294 42970 208350
rect 43026 208294 43094 208350
rect 43150 208294 43218 208350
rect 43274 208294 43342 208350
rect 43398 208294 43494 208350
rect 42874 208226 43494 208294
rect 42874 208170 42970 208226
rect 43026 208170 43094 208226
rect 43150 208170 43218 208226
rect 43274 208170 43342 208226
rect 43398 208170 43494 208226
rect 42874 208102 43494 208170
rect 42874 208046 42970 208102
rect 43026 208046 43094 208102
rect 43150 208046 43218 208102
rect 43274 208046 43342 208102
rect 43398 208046 43494 208102
rect 42874 207978 43494 208046
rect 42874 207922 42970 207978
rect 43026 207922 43094 207978
rect 43150 207922 43218 207978
rect 43274 207922 43342 207978
rect 43398 207922 43494 207978
rect 39154 184294 39250 184350
rect 39306 184294 39374 184350
rect 39430 184294 39498 184350
rect 39554 184294 39622 184350
rect 39678 184294 39774 184350
rect 39154 184226 39774 184294
rect 39154 184170 39250 184226
rect 39306 184170 39374 184226
rect 39430 184170 39498 184226
rect 39554 184170 39622 184226
rect 39678 184170 39774 184226
rect 39154 184102 39774 184170
rect 39154 184046 39250 184102
rect 39306 184046 39374 184102
rect 39430 184046 39498 184102
rect 39554 184046 39622 184102
rect 39678 184046 39774 184102
rect 39154 183978 39774 184046
rect 39154 183922 39250 183978
rect 39306 183922 39374 183978
rect 39430 183922 39498 183978
rect 39554 183922 39622 183978
rect 39678 183922 39774 183978
rect 39154 166350 39774 183922
rect 39154 166294 39250 166350
rect 39306 166294 39374 166350
rect 39430 166294 39498 166350
rect 39554 166294 39622 166350
rect 39678 166294 39774 166350
rect 39154 166226 39774 166294
rect 39154 166170 39250 166226
rect 39306 166170 39374 166226
rect 39430 166170 39498 166226
rect 39554 166170 39622 166226
rect 39678 166170 39774 166226
rect 39154 166102 39774 166170
rect 39154 166046 39250 166102
rect 39306 166046 39374 166102
rect 39430 166046 39498 166102
rect 39554 166046 39622 166102
rect 39678 166046 39774 166102
rect 39154 165978 39774 166046
rect 39154 165922 39250 165978
rect 39306 165922 39374 165978
rect 39430 165922 39498 165978
rect 39554 165922 39622 165978
rect 39678 165922 39774 165978
rect 39154 148350 39774 165922
rect 39154 148294 39250 148350
rect 39306 148294 39374 148350
rect 39430 148294 39498 148350
rect 39554 148294 39622 148350
rect 39678 148294 39774 148350
rect 39154 148226 39774 148294
rect 39154 148170 39250 148226
rect 39306 148170 39374 148226
rect 39430 148170 39498 148226
rect 39554 148170 39622 148226
rect 39678 148170 39774 148226
rect 39154 148102 39774 148170
rect 39154 148046 39250 148102
rect 39306 148046 39374 148102
rect 39430 148046 39498 148102
rect 39554 148046 39622 148102
rect 39678 148046 39774 148102
rect 39154 147978 39774 148046
rect 39154 147922 39250 147978
rect 39306 147922 39374 147978
rect 39430 147922 39498 147978
rect 39554 147922 39622 147978
rect 39678 147922 39774 147978
rect 36204 120082 36260 120092
rect 39154 130350 39774 147922
rect 39154 130294 39250 130350
rect 39306 130294 39374 130350
rect 39430 130294 39498 130350
rect 39554 130294 39622 130350
rect 39678 130294 39774 130350
rect 39154 130226 39774 130294
rect 39154 130170 39250 130226
rect 39306 130170 39374 130226
rect 39430 130170 39498 130226
rect 39554 130170 39622 130226
rect 39678 130170 39774 130226
rect 39154 130102 39774 130170
rect 39154 130046 39250 130102
rect 39306 130046 39374 130102
rect 39430 130046 39498 130102
rect 39554 130046 39622 130102
rect 39678 130046 39774 130102
rect 39154 129978 39774 130046
rect 39154 129922 39250 129978
rect 39306 129922 39374 129978
rect 39430 129922 39498 129978
rect 39554 129922 39622 129978
rect 39678 129922 39774 129978
rect 34524 107090 34580 107100
rect 39154 112350 39774 129922
rect 39154 112294 39250 112350
rect 39306 112294 39374 112350
rect 39430 112294 39498 112350
rect 39554 112294 39622 112350
rect 39678 112294 39774 112350
rect 39154 112226 39774 112294
rect 39154 112170 39250 112226
rect 39306 112170 39374 112226
rect 39430 112170 39498 112226
rect 39554 112170 39622 112226
rect 39678 112170 39774 112226
rect 39154 112102 39774 112170
rect 39154 112046 39250 112102
rect 39306 112046 39374 112102
rect 39430 112046 39498 112102
rect 39554 112046 39622 112102
rect 39678 112046 39774 112102
rect 39154 111978 39774 112046
rect 39154 111922 39250 111978
rect 39306 111922 39374 111978
rect 39430 111922 39498 111978
rect 39554 111922 39622 111978
rect 39678 111922 39774 111978
rect 29484 88050 29540 88060
rect 39154 94350 39774 111922
rect 39154 94294 39250 94350
rect 39306 94294 39374 94350
rect 39430 94294 39498 94350
rect 39554 94294 39622 94350
rect 39678 94294 39774 94350
rect 39154 94226 39774 94294
rect 39154 94170 39250 94226
rect 39306 94170 39374 94226
rect 39430 94170 39498 94226
rect 39554 94170 39622 94226
rect 39678 94170 39774 94226
rect 39154 94102 39774 94170
rect 39154 94046 39250 94102
rect 39306 94046 39374 94102
rect 39430 94046 39498 94102
rect 39554 94046 39622 94102
rect 39678 94046 39774 94102
rect 39154 93978 39774 94046
rect 39154 93922 39250 93978
rect 39306 93922 39374 93978
rect 39430 93922 39498 93978
rect 39554 93922 39622 93978
rect 39678 93922 39774 93978
rect 24874 82294 24970 82350
rect 25026 82294 25094 82350
rect 25150 82294 25218 82350
rect 25274 82294 25342 82350
rect 25398 82294 25494 82350
rect 24874 82226 25494 82294
rect 24874 82170 24970 82226
rect 25026 82170 25094 82226
rect 25150 82170 25218 82226
rect 25274 82170 25342 82226
rect 25398 82170 25494 82226
rect 24874 82102 25494 82170
rect 24874 82046 24970 82102
rect 25026 82046 25094 82102
rect 25150 82046 25218 82102
rect 25274 82046 25342 82102
rect 25398 82046 25494 82102
rect 24874 81978 25494 82046
rect 24874 81922 24970 81978
rect 25026 81922 25094 81978
rect 25150 81922 25218 81978
rect 25274 81922 25342 81978
rect 25398 81922 25494 81978
rect 24874 64350 25494 81922
rect 24874 64294 24970 64350
rect 25026 64294 25094 64350
rect 25150 64294 25218 64350
rect 25274 64294 25342 64350
rect 25398 64294 25494 64350
rect 24874 64226 25494 64294
rect 24874 64170 24970 64226
rect 25026 64170 25094 64226
rect 25150 64170 25218 64226
rect 25274 64170 25342 64226
rect 25398 64170 25494 64226
rect 24874 64102 25494 64170
rect 24874 64046 24970 64102
rect 25026 64046 25094 64102
rect 25150 64046 25218 64102
rect 25274 64046 25342 64102
rect 25398 64046 25494 64102
rect 24874 63978 25494 64046
rect 24874 63922 24970 63978
rect 25026 63922 25094 63978
rect 25150 63922 25218 63978
rect 25274 63922 25342 63978
rect 25398 63922 25494 63978
rect 24874 46350 25494 63922
rect 24874 46294 24970 46350
rect 25026 46294 25094 46350
rect 25150 46294 25218 46350
rect 25274 46294 25342 46350
rect 25398 46294 25494 46350
rect 24874 46226 25494 46294
rect 24874 46170 24970 46226
rect 25026 46170 25094 46226
rect 25150 46170 25218 46226
rect 25274 46170 25342 46226
rect 25398 46170 25494 46226
rect 24874 46102 25494 46170
rect 24874 46046 24970 46102
rect 25026 46046 25094 46102
rect 25150 46046 25218 46102
rect 25274 46046 25342 46102
rect 25398 46046 25494 46102
rect 24874 45978 25494 46046
rect 24874 45922 24970 45978
rect 25026 45922 25094 45978
rect 25150 45922 25218 45978
rect 25274 45922 25342 45978
rect 25398 45922 25494 45978
rect 24874 28350 25494 45922
rect 24874 28294 24970 28350
rect 25026 28294 25094 28350
rect 25150 28294 25218 28350
rect 25274 28294 25342 28350
rect 25398 28294 25494 28350
rect 24874 28226 25494 28294
rect 24874 28170 24970 28226
rect 25026 28170 25094 28226
rect 25150 28170 25218 28226
rect 25274 28170 25342 28226
rect 25398 28170 25494 28226
rect 24874 28102 25494 28170
rect 24874 28046 24970 28102
rect 25026 28046 25094 28102
rect 25150 28046 25218 28102
rect 25274 28046 25342 28102
rect 25398 28046 25494 28102
rect 24874 27978 25494 28046
rect 24874 27922 24970 27978
rect 25026 27922 25094 27978
rect 25150 27922 25218 27978
rect 25274 27922 25342 27978
rect 25398 27922 25494 27978
rect 24874 10350 25494 27922
rect 24874 10294 24970 10350
rect 25026 10294 25094 10350
rect 25150 10294 25218 10350
rect 25274 10294 25342 10350
rect 25398 10294 25494 10350
rect 24874 10226 25494 10294
rect 24874 10170 24970 10226
rect 25026 10170 25094 10226
rect 25150 10170 25218 10226
rect 25274 10170 25342 10226
rect 25398 10170 25494 10226
rect 24874 10102 25494 10170
rect 24874 10046 24970 10102
rect 25026 10046 25094 10102
rect 25150 10046 25218 10102
rect 25274 10046 25342 10102
rect 25398 10046 25494 10102
rect 24874 9978 25494 10046
rect 24874 9922 24970 9978
rect 25026 9922 25094 9978
rect 25150 9922 25218 9978
rect 25274 9922 25342 9978
rect 25398 9922 25494 9978
rect 24874 -1120 25494 9922
rect 24874 -1176 24970 -1120
rect 25026 -1176 25094 -1120
rect 25150 -1176 25218 -1120
rect 25274 -1176 25342 -1120
rect 25398 -1176 25494 -1120
rect 24874 -1244 25494 -1176
rect 24874 -1300 24970 -1244
rect 25026 -1300 25094 -1244
rect 25150 -1300 25218 -1244
rect 25274 -1300 25342 -1244
rect 25398 -1300 25494 -1244
rect 24874 -1368 25494 -1300
rect 24874 -1424 24970 -1368
rect 25026 -1424 25094 -1368
rect 25150 -1424 25218 -1368
rect 25274 -1424 25342 -1368
rect 25398 -1424 25494 -1368
rect 24874 -1492 25494 -1424
rect 24874 -1548 24970 -1492
rect 25026 -1548 25094 -1492
rect 25150 -1548 25218 -1492
rect 25274 -1548 25342 -1492
rect 25398 -1548 25494 -1492
rect 24874 -1644 25494 -1548
rect 39154 76350 39774 93922
rect 41132 192052 41188 192062
rect 41132 89908 41188 191996
rect 41132 89842 41188 89852
rect 42874 190350 43494 207922
rect 42874 190294 42970 190350
rect 43026 190294 43094 190350
rect 43150 190294 43218 190350
rect 43274 190294 43342 190350
rect 43398 190294 43494 190350
rect 42874 190226 43494 190294
rect 42874 190170 42970 190226
rect 43026 190170 43094 190226
rect 43150 190170 43218 190226
rect 43274 190170 43342 190226
rect 43398 190170 43494 190226
rect 42874 190102 43494 190170
rect 42874 190046 42970 190102
rect 43026 190046 43094 190102
rect 43150 190046 43218 190102
rect 43274 190046 43342 190102
rect 43398 190046 43494 190102
rect 42874 189978 43494 190046
rect 42874 189922 42970 189978
rect 43026 189922 43094 189978
rect 43150 189922 43218 189978
rect 43274 189922 43342 189978
rect 43398 189922 43494 189978
rect 42874 172350 43494 189922
rect 42874 172294 42970 172350
rect 43026 172294 43094 172350
rect 43150 172294 43218 172350
rect 43274 172294 43342 172350
rect 43398 172294 43494 172350
rect 42874 172226 43494 172294
rect 42874 172170 42970 172226
rect 43026 172170 43094 172226
rect 43150 172170 43218 172226
rect 43274 172170 43342 172226
rect 43398 172170 43494 172226
rect 42874 172102 43494 172170
rect 42874 172046 42970 172102
rect 43026 172046 43094 172102
rect 43150 172046 43218 172102
rect 43274 172046 43342 172102
rect 43398 172046 43494 172102
rect 42874 171978 43494 172046
rect 42874 171922 42970 171978
rect 43026 171922 43094 171978
rect 43150 171922 43218 171978
rect 43274 171922 43342 171978
rect 43398 171922 43494 171978
rect 42874 154350 43494 171922
rect 42874 154294 42970 154350
rect 43026 154294 43094 154350
rect 43150 154294 43218 154350
rect 43274 154294 43342 154350
rect 43398 154294 43494 154350
rect 42874 154226 43494 154294
rect 42874 154170 42970 154226
rect 43026 154170 43094 154226
rect 43150 154170 43218 154226
rect 43274 154170 43342 154226
rect 43398 154170 43494 154226
rect 42874 154102 43494 154170
rect 42874 154046 42970 154102
rect 43026 154046 43094 154102
rect 43150 154046 43218 154102
rect 43274 154046 43342 154102
rect 43398 154046 43494 154102
rect 42874 153978 43494 154046
rect 42874 153922 42970 153978
rect 43026 153922 43094 153978
rect 43150 153922 43218 153978
rect 43274 153922 43342 153978
rect 43398 153922 43494 153978
rect 42874 136350 43494 153922
rect 42874 136294 42970 136350
rect 43026 136294 43094 136350
rect 43150 136294 43218 136350
rect 43274 136294 43342 136350
rect 43398 136294 43494 136350
rect 42874 136226 43494 136294
rect 42874 136170 42970 136226
rect 43026 136170 43094 136226
rect 43150 136170 43218 136226
rect 43274 136170 43342 136226
rect 43398 136170 43494 136226
rect 42874 136102 43494 136170
rect 42874 136046 42970 136102
rect 43026 136046 43094 136102
rect 43150 136046 43218 136102
rect 43274 136046 43342 136102
rect 43398 136046 43494 136102
rect 42874 135978 43494 136046
rect 42874 135922 42970 135978
rect 43026 135922 43094 135978
rect 43150 135922 43218 135978
rect 43274 135922 43342 135978
rect 43398 135922 43494 135978
rect 42874 118350 43494 135922
rect 42874 118294 42970 118350
rect 43026 118294 43094 118350
rect 43150 118294 43218 118350
rect 43274 118294 43342 118350
rect 43398 118294 43494 118350
rect 42874 118226 43494 118294
rect 42874 118170 42970 118226
rect 43026 118170 43094 118226
rect 43150 118170 43218 118226
rect 43274 118170 43342 118226
rect 43398 118170 43494 118226
rect 42874 118102 43494 118170
rect 42874 118046 42970 118102
rect 43026 118046 43094 118102
rect 43150 118046 43218 118102
rect 43274 118046 43342 118102
rect 43398 118046 43494 118102
rect 42874 117978 43494 118046
rect 42874 117922 42970 117978
rect 43026 117922 43094 117978
rect 43150 117922 43218 117978
rect 43274 117922 43342 117978
rect 43398 117922 43494 117978
rect 42874 100350 43494 117922
rect 42874 100294 42970 100350
rect 43026 100294 43094 100350
rect 43150 100294 43218 100350
rect 43274 100294 43342 100350
rect 43398 100294 43494 100350
rect 42874 100226 43494 100294
rect 42874 100170 42970 100226
rect 43026 100170 43094 100226
rect 43150 100170 43218 100226
rect 43274 100170 43342 100226
rect 43398 100170 43494 100226
rect 42874 100102 43494 100170
rect 42874 100046 42970 100102
rect 43026 100046 43094 100102
rect 43150 100046 43218 100102
rect 43274 100046 43342 100102
rect 43398 100046 43494 100102
rect 42874 99978 43494 100046
rect 42874 99922 42970 99978
rect 43026 99922 43094 99978
rect 43150 99922 43218 99978
rect 43274 99922 43342 99978
rect 43398 99922 43494 99978
rect 39154 76294 39250 76350
rect 39306 76294 39374 76350
rect 39430 76294 39498 76350
rect 39554 76294 39622 76350
rect 39678 76294 39774 76350
rect 39154 76226 39774 76294
rect 39154 76170 39250 76226
rect 39306 76170 39374 76226
rect 39430 76170 39498 76226
rect 39554 76170 39622 76226
rect 39678 76170 39774 76226
rect 39154 76102 39774 76170
rect 39154 76046 39250 76102
rect 39306 76046 39374 76102
rect 39430 76046 39498 76102
rect 39554 76046 39622 76102
rect 39678 76046 39774 76102
rect 39154 75978 39774 76046
rect 39154 75922 39250 75978
rect 39306 75922 39374 75978
rect 39430 75922 39498 75978
rect 39554 75922 39622 75978
rect 39678 75922 39774 75978
rect 39154 58350 39774 75922
rect 39154 58294 39250 58350
rect 39306 58294 39374 58350
rect 39430 58294 39498 58350
rect 39554 58294 39622 58350
rect 39678 58294 39774 58350
rect 39154 58226 39774 58294
rect 39154 58170 39250 58226
rect 39306 58170 39374 58226
rect 39430 58170 39498 58226
rect 39554 58170 39622 58226
rect 39678 58170 39774 58226
rect 39154 58102 39774 58170
rect 39154 58046 39250 58102
rect 39306 58046 39374 58102
rect 39430 58046 39498 58102
rect 39554 58046 39622 58102
rect 39678 58046 39774 58102
rect 39154 57978 39774 58046
rect 39154 57922 39250 57978
rect 39306 57922 39374 57978
rect 39430 57922 39498 57978
rect 39554 57922 39622 57978
rect 39678 57922 39774 57978
rect 39154 40350 39774 57922
rect 39154 40294 39250 40350
rect 39306 40294 39374 40350
rect 39430 40294 39498 40350
rect 39554 40294 39622 40350
rect 39678 40294 39774 40350
rect 39154 40226 39774 40294
rect 39154 40170 39250 40226
rect 39306 40170 39374 40226
rect 39430 40170 39498 40226
rect 39554 40170 39622 40226
rect 39678 40170 39774 40226
rect 39154 40102 39774 40170
rect 39154 40046 39250 40102
rect 39306 40046 39374 40102
rect 39430 40046 39498 40102
rect 39554 40046 39622 40102
rect 39678 40046 39774 40102
rect 39154 39978 39774 40046
rect 39154 39922 39250 39978
rect 39306 39922 39374 39978
rect 39430 39922 39498 39978
rect 39554 39922 39622 39978
rect 39678 39922 39774 39978
rect 39154 22350 39774 39922
rect 39154 22294 39250 22350
rect 39306 22294 39374 22350
rect 39430 22294 39498 22350
rect 39554 22294 39622 22350
rect 39678 22294 39774 22350
rect 39154 22226 39774 22294
rect 39154 22170 39250 22226
rect 39306 22170 39374 22226
rect 39430 22170 39498 22226
rect 39554 22170 39622 22226
rect 39678 22170 39774 22226
rect 39154 22102 39774 22170
rect 39154 22046 39250 22102
rect 39306 22046 39374 22102
rect 39430 22046 39498 22102
rect 39554 22046 39622 22102
rect 39678 22046 39774 22102
rect 39154 21978 39774 22046
rect 39154 21922 39250 21978
rect 39306 21922 39374 21978
rect 39430 21922 39498 21978
rect 39554 21922 39622 21978
rect 39678 21922 39774 21978
rect 39154 4350 39774 21922
rect 39154 4294 39250 4350
rect 39306 4294 39374 4350
rect 39430 4294 39498 4350
rect 39554 4294 39622 4350
rect 39678 4294 39774 4350
rect 39154 4226 39774 4294
rect 39154 4170 39250 4226
rect 39306 4170 39374 4226
rect 39430 4170 39498 4226
rect 39554 4170 39622 4226
rect 39678 4170 39774 4226
rect 39154 4102 39774 4170
rect 39154 4046 39250 4102
rect 39306 4046 39374 4102
rect 39430 4046 39498 4102
rect 39554 4046 39622 4102
rect 39678 4046 39774 4102
rect 39154 3978 39774 4046
rect 39154 3922 39250 3978
rect 39306 3922 39374 3978
rect 39430 3922 39498 3978
rect 39554 3922 39622 3978
rect 39678 3922 39774 3978
rect 39154 -160 39774 3922
rect 39154 -216 39250 -160
rect 39306 -216 39374 -160
rect 39430 -216 39498 -160
rect 39554 -216 39622 -160
rect 39678 -216 39774 -160
rect 39154 -284 39774 -216
rect 39154 -340 39250 -284
rect 39306 -340 39374 -284
rect 39430 -340 39498 -284
rect 39554 -340 39622 -284
rect 39678 -340 39774 -284
rect 39154 -408 39774 -340
rect 39154 -464 39250 -408
rect 39306 -464 39374 -408
rect 39430 -464 39498 -408
rect 39554 -464 39622 -408
rect 39678 -464 39774 -408
rect 39154 -532 39774 -464
rect 39154 -588 39250 -532
rect 39306 -588 39374 -532
rect 39430 -588 39498 -532
rect 39554 -588 39622 -532
rect 39678 -588 39774 -532
rect 39154 -1644 39774 -588
rect 42874 82350 43494 99922
rect 44492 234388 44548 234398
rect 44492 96628 44548 234332
rect 57154 220350 57774 237922
rect 57154 220294 57250 220350
rect 57306 220294 57374 220350
rect 57430 220294 57498 220350
rect 57554 220294 57622 220350
rect 57678 220294 57774 220350
rect 57154 220226 57774 220294
rect 57154 220170 57250 220226
rect 57306 220170 57374 220226
rect 57430 220170 57498 220226
rect 57554 220170 57622 220226
rect 57678 220170 57774 220226
rect 57154 220102 57774 220170
rect 57154 220046 57250 220102
rect 57306 220046 57374 220102
rect 57430 220046 57498 220102
rect 57554 220046 57622 220102
rect 57678 220046 57774 220102
rect 57154 219978 57774 220046
rect 57154 219922 57250 219978
rect 57306 219922 57374 219978
rect 57430 219922 57498 219978
rect 57554 219922 57622 219978
rect 57678 219922 57774 219978
rect 57154 202350 57774 219922
rect 60874 598172 61494 598268
rect 60874 598116 60970 598172
rect 61026 598116 61094 598172
rect 61150 598116 61218 598172
rect 61274 598116 61342 598172
rect 61398 598116 61494 598172
rect 60874 598048 61494 598116
rect 60874 597992 60970 598048
rect 61026 597992 61094 598048
rect 61150 597992 61218 598048
rect 61274 597992 61342 598048
rect 61398 597992 61494 598048
rect 60874 597924 61494 597992
rect 60874 597868 60970 597924
rect 61026 597868 61094 597924
rect 61150 597868 61218 597924
rect 61274 597868 61342 597924
rect 61398 597868 61494 597924
rect 60874 597800 61494 597868
rect 60874 597744 60970 597800
rect 61026 597744 61094 597800
rect 61150 597744 61218 597800
rect 61274 597744 61342 597800
rect 61398 597744 61494 597800
rect 60874 586350 61494 597744
rect 78874 598172 79494 598268
rect 78874 598116 78970 598172
rect 79026 598116 79094 598172
rect 79150 598116 79218 598172
rect 79274 598116 79342 598172
rect 79398 598116 79494 598172
rect 78874 598048 79494 598116
rect 78874 597992 78970 598048
rect 79026 597992 79094 598048
rect 79150 597992 79218 598048
rect 79274 597992 79342 598048
rect 79398 597992 79494 598048
rect 78874 597924 79494 597992
rect 78874 597868 78970 597924
rect 79026 597868 79094 597924
rect 79150 597868 79218 597924
rect 79274 597868 79342 597924
rect 79398 597868 79494 597924
rect 78874 597800 79494 597868
rect 78874 597744 78970 597800
rect 79026 597744 79094 597800
rect 79150 597744 79218 597800
rect 79274 597744 79342 597800
rect 79398 597744 79494 597800
rect 77308 589764 77364 589774
rect 77308 588868 77364 589708
rect 77308 588802 77364 588812
rect 60874 586294 60970 586350
rect 61026 586294 61094 586350
rect 61150 586294 61218 586350
rect 61274 586294 61342 586350
rect 61398 586294 61494 586350
rect 60874 586226 61494 586294
rect 60874 586170 60970 586226
rect 61026 586170 61094 586226
rect 61150 586170 61218 586226
rect 61274 586170 61342 586226
rect 61398 586170 61494 586226
rect 60874 586102 61494 586170
rect 60874 586046 60970 586102
rect 61026 586046 61094 586102
rect 61150 586046 61218 586102
rect 61274 586046 61342 586102
rect 61398 586046 61494 586102
rect 60874 585978 61494 586046
rect 60874 585922 60970 585978
rect 61026 585922 61094 585978
rect 61150 585922 61218 585978
rect 61274 585922 61342 585978
rect 61398 585922 61494 585978
rect 60874 568350 61494 585922
rect 60874 568294 60970 568350
rect 61026 568294 61094 568350
rect 61150 568294 61218 568350
rect 61274 568294 61342 568350
rect 61398 568294 61494 568350
rect 60874 568226 61494 568294
rect 60874 568170 60970 568226
rect 61026 568170 61094 568226
rect 61150 568170 61218 568226
rect 61274 568170 61342 568226
rect 61398 568170 61494 568226
rect 60874 568102 61494 568170
rect 60874 568046 60970 568102
rect 61026 568046 61094 568102
rect 61150 568046 61218 568102
rect 61274 568046 61342 568102
rect 61398 568046 61494 568102
rect 60874 567978 61494 568046
rect 60874 567922 60970 567978
rect 61026 567922 61094 567978
rect 61150 567922 61218 567978
rect 61274 567922 61342 567978
rect 61398 567922 61494 567978
rect 60874 550350 61494 567922
rect 60874 550294 60970 550350
rect 61026 550294 61094 550350
rect 61150 550294 61218 550350
rect 61274 550294 61342 550350
rect 61398 550294 61494 550350
rect 60874 550226 61494 550294
rect 60874 550170 60970 550226
rect 61026 550170 61094 550226
rect 61150 550170 61218 550226
rect 61274 550170 61342 550226
rect 61398 550170 61494 550226
rect 60874 550102 61494 550170
rect 60874 550046 60970 550102
rect 61026 550046 61094 550102
rect 61150 550046 61218 550102
rect 61274 550046 61342 550102
rect 61398 550046 61494 550102
rect 60874 549978 61494 550046
rect 60874 549922 60970 549978
rect 61026 549922 61094 549978
rect 61150 549922 61218 549978
rect 61274 549922 61342 549978
rect 61398 549922 61494 549978
rect 60874 532350 61494 549922
rect 60874 532294 60970 532350
rect 61026 532294 61094 532350
rect 61150 532294 61218 532350
rect 61274 532294 61342 532350
rect 61398 532294 61494 532350
rect 60874 532226 61494 532294
rect 60874 532170 60970 532226
rect 61026 532170 61094 532226
rect 61150 532170 61218 532226
rect 61274 532170 61342 532226
rect 61398 532170 61494 532226
rect 60874 532102 61494 532170
rect 60874 532046 60970 532102
rect 61026 532046 61094 532102
rect 61150 532046 61218 532102
rect 61274 532046 61342 532102
rect 61398 532046 61494 532102
rect 60874 531978 61494 532046
rect 60874 531922 60970 531978
rect 61026 531922 61094 531978
rect 61150 531922 61218 531978
rect 61274 531922 61342 531978
rect 61398 531922 61494 531978
rect 60874 514350 61494 531922
rect 60874 514294 60970 514350
rect 61026 514294 61094 514350
rect 61150 514294 61218 514350
rect 61274 514294 61342 514350
rect 61398 514294 61494 514350
rect 60874 514226 61494 514294
rect 60874 514170 60970 514226
rect 61026 514170 61094 514226
rect 61150 514170 61218 514226
rect 61274 514170 61342 514226
rect 61398 514170 61494 514226
rect 60874 514102 61494 514170
rect 60874 514046 60970 514102
rect 61026 514046 61094 514102
rect 61150 514046 61218 514102
rect 61274 514046 61342 514102
rect 61398 514046 61494 514102
rect 60874 513978 61494 514046
rect 60874 513922 60970 513978
rect 61026 513922 61094 513978
rect 61150 513922 61218 513978
rect 61274 513922 61342 513978
rect 61398 513922 61494 513978
rect 60874 496350 61494 513922
rect 60874 496294 60970 496350
rect 61026 496294 61094 496350
rect 61150 496294 61218 496350
rect 61274 496294 61342 496350
rect 61398 496294 61494 496350
rect 60874 496226 61494 496294
rect 60874 496170 60970 496226
rect 61026 496170 61094 496226
rect 61150 496170 61218 496226
rect 61274 496170 61342 496226
rect 61398 496170 61494 496226
rect 60874 496102 61494 496170
rect 60874 496046 60970 496102
rect 61026 496046 61094 496102
rect 61150 496046 61218 496102
rect 61274 496046 61342 496102
rect 61398 496046 61494 496102
rect 60874 495978 61494 496046
rect 60874 495922 60970 495978
rect 61026 495922 61094 495978
rect 61150 495922 61218 495978
rect 61274 495922 61342 495978
rect 61398 495922 61494 495978
rect 60874 478350 61494 495922
rect 60874 478294 60970 478350
rect 61026 478294 61094 478350
rect 61150 478294 61218 478350
rect 61274 478294 61342 478350
rect 61398 478294 61494 478350
rect 60874 478226 61494 478294
rect 60874 478170 60970 478226
rect 61026 478170 61094 478226
rect 61150 478170 61218 478226
rect 61274 478170 61342 478226
rect 61398 478170 61494 478226
rect 60874 478102 61494 478170
rect 60874 478046 60970 478102
rect 61026 478046 61094 478102
rect 61150 478046 61218 478102
rect 61274 478046 61342 478102
rect 61398 478046 61494 478102
rect 60874 477978 61494 478046
rect 60874 477922 60970 477978
rect 61026 477922 61094 477978
rect 61150 477922 61218 477978
rect 61274 477922 61342 477978
rect 61398 477922 61494 477978
rect 60874 460350 61494 477922
rect 60874 460294 60970 460350
rect 61026 460294 61094 460350
rect 61150 460294 61218 460350
rect 61274 460294 61342 460350
rect 61398 460294 61494 460350
rect 60874 460226 61494 460294
rect 60874 460170 60970 460226
rect 61026 460170 61094 460226
rect 61150 460170 61218 460226
rect 61274 460170 61342 460226
rect 61398 460170 61494 460226
rect 60874 460102 61494 460170
rect 60874 460046 60970 460102
rect 61026 460046 61094 460102
rect 61150 460046 61218 460102
rect 61274 460046 61342 460102
rect 61398 460046 61494 460102
rect 60874 459978 61494 460046
rect 60874 459922 60970 459978
rect 61026 459922 61094 459978
rect 61150 459922 61218 459978
rect 61274 459922 61342 459978
rect 61398 459922 61494 459978
rect 60874 442350 61494 459922
rect 60874 442294 60970 442350
rect 61026 442294 61094 442350
rect 61150 442294 61218 442350
rect 61274 442294 61342 442350
rect 61398 442294 61494 442350
rect 60874 442226 61494 442294
rect 60874 442170 60970 442226
rect 61026 442170 61094 442226
rect 61150 442170 61218 442226
rect 61274 442170 61342 442226
rect 61398 442170 61494 442226
rect 60874 442102 61494 442170
rect 60874 442046 60970 442102
rect 61026 442046 61094 442102
rect 61150 442046 61218 442102
rect 61274 442046 61342 442102
rect 61398 442046 61494 442102
rect 60874 441978 61494 442046
rect 60874 441922 60970 441978
rect 61026 441922 61094 441978
rect 61150 441922 61218 441978
rect 61274 441922 61342 441978
rect 61398 441922 61494 441978
rect 60874 424350 61494 441922
rect 60874 424294 60970 424350
rect 61026 424294 61094 424350
rect 61150 424294 61218 424350
rect 61274 424294 61342 424350
rect 61398 424294 61494 424350
rect 60874 424226 61494 424294
rect 60874 424170 60970 424226
rect 61026 424170 61094 424226
rect 61150 424170 61218 424226
rect 61274 424170 61342 424226
rect 61398 424170 61494 424226
rect 60874 424102 61494 424170
rect 60874 424046 60970 424102
rect 61026 424046 61094 424102
rect 61150 424046 61218 424102
rect 61274 424046 61342 424102
rect 61398 424046 61494 424102
rect 60874 423978 61494 424046
rect 60874 423922 60970 423978
rect 61026 423922 61094 423978
rect 61150 423922 61218 423978
rect 61274 423922 61342 423978
rect 61398 423922 61494 423978
rect 60874 406350 61494 423922
rect 60874 406294 60970 406350
rect 61026 406294 61094 406350
rect 61150 406294 61218 406350
rect 61274 406294 61342 406350
rect 61398 406294 61494 406350
rect 60874 406226 61494 406294
rect 60874 406170 60970 406226
rect 61026 406170 61094 406226
rect 61150 406170 61218 406226
rect 61274 406170 61342 406226
rect 61398 406170 61494 406226
rect 60874 406102 61494 406170
rect 60874 406046 60970 406102
rect 61026 406046 61094 406102
rect 61150 406046 61218 406102
rect 61274 406046 61342 406102
rect 61398 406046 61494 406102
rect 60874 405978 61494 406046
rect 60874 405922 60970 405978
rect 61026 405922 61094 405978
rect 61150 405922 61218 405978
rect 61274 405922 61342 405978
rect 61398 405922 61494 405978
rect 60874 388350 61494 405922
rect 60874 388294 60970 388350
rect 61026 388294 61094 388350
rect 61150 388294 61218 388350
rect 61274 388294 61342 388350
rect 61398 388294 61494 388350
rect 60874 388226 61494 388294
rect 60874 388170 60970 388226
rect 61026 388170 61094 388226
rect 61150 388170 61218 388226
rect 61274 388170 61342 388226
rect 61398 388170 61494 388226
rect 60874 388102 61494 388170
rect 60874 388046 60970 388102
rect 61026 388046 61094 388102
rect 61150 388046 61218 388102
rect 61274 388046 61342 388102
rect 61398 388046 61494 388102
rect 60874 387978 61494 388046
rect 60874 387922 60970 387978
rect 61026 387922 61094 387978
rect 61150 387922 61218 387978
rect 61274 387922 61342 387978
rect 61398 387922 61494 387978
rect 60874 370350 61494 387922
rect 60874 370294 60970 370350
rect 61026 370294 61094 370350
rect 61150 370294 61218 370350
rect 61274 370294 61342 370350
rect 61398 370294 61494 370350
rect 60874 370226 61494 370294
rect 60874 370170 60970 370226
rect 61026 370170 61094 370226
rect 61150 370170 61218 370226
rect 61274 370170 61342 370226
rect 61398 370170 61494 370226
rect 60874 370102 61494 370170
rect 60874 370046 60970 370102
rect 61026 370046 61094 370102
rect 61150 370046 61218 370102
rect 61274 370046 61342 370102
rect 61398 370046 61494 370102
rect 60874 369978 61494 370046
rect 60874 369922 60970 369978
rect 61026 369922 61094 369978
rect 61150 369922 61218 369978
rect 61274 369922 61342 369978
rect 61398 369922 61494 369978
rect 60874 352350 61494 369922
rect 60874 352294 60970 352350
rect 61026 352294 61094 352350
rect 61150 352294 61218 352350
rect 61274 352294 61342 352350
rect 61398 352294 61494 352350
rect 60874 352226 61494 352294
rect 60874 352170 60970 352226
rect 61026 352170 61094 352226
rect 61150 352170 61218 352226
rect 61274 352170 61342 352226
rect 61398 352170 61494 352226
rect 60874 352102 61494 352170
rect 60874 352046 60970 352102
rect 61026 352046 61094 352102
rect 61150 352046 61218 352102
rect 61274 352046 61342 352102
rect 61398 352046 61494 352102
rect 60874 351978 61494 352046
rect 60874 351922 60970 351978
rect 61026 351922 61094 351978
rect 61150 351922 61218 351978
rect 61274 351922 61342 351978
rect 61398 351922 61494 351978
rect 60874 334350 61494 351922
rect 60874 334294 60970 334350
rect 61026 334294 61094 334350
rect 61150 334294 61218 334350
rect 61274 334294 61342 334350
rect 61398 334294 61494 334350
rect 60874 334226 61494 334294
rect 60874 334170 60970 334226
rect 61026 334170 61094 334226
rect 61150 334170 61218 334226
rect 61274 334170 61342 334226
rect 61398 334170 61494 334226
rect 60874 334102 61494 334170
rect 60874 334046 60970 334102
rect 61026 334046 61094 334102
rect 61150 334046 61218 334102
rect 61274 334046 61342 334102
rect 61398 334046 61494 334102
rect 60874 333978 61494 334046
rect 60874 333922 60970 333978
rect 61026 333922 61094 333978
rect 61150 333922 61218 333978
rect 61274 333922 61342 333978
rect 61398 333922 61494 333978
rect 60874 316350 61494 333922
rect 60874 316294 60970 316350
rect 61026 316294 61094 316350
rect 61150 316294 61218 316350
rect 61274 316294 61342 316350
rect 61398 316294 61494 316350
rect 60874 316226 61494 316294
rect 60874 316170 60970 316226
rect 61026 316170 61094 316226
rect 61150 316170 61218 316226
rect 61274 316170 61342 316226
rect 61398 316170 61494 316226
rect 60874 316102 61494 316170
rect 60874 316046 60970 316102
rect 61026 316046 61094 316102
rect 61150 316046 61218 316102
rect 61274 316046 61342 316102
rect 61398 316046 61494 316102
rect 60874 315978 61494 316046
rect 60874 315922 60970 315978
rect 61026 315922 61094 315978
rect 61150 315922 61218 315978
rect 61274 315922 61342 315978
rect 61398 315922 61494 315978
rect 60874 298350 61494 315922
rect 60874 298294 60970 298350
rect 61026 298294 61094 298350
rect 61150 298294 61218 298350
rect 61274 298294 61342 298350
rect 61398 298294 61494 298350
rect 60874 298226 61494 298294
rect 60874 298170 60970 298226
rect 61026 298170 61094 298226
rect 61150 298170 61218 298226
rect 61274 298170 61342 298226
rect 61398 298170 61494 298226
rect 60874 298102 61494 298170
rect 60874 298046 60970 298102
rect 61026 298046 61094 298102
rect 61150 298046 61218 298102
rect 61274 298046 61342 298102
rect 61398 298046 61494 298102
rect 60874 297978 61494 298046
rect 60874 297922 60970 297978
rect 61026 297922 61094 297978
rect 61150 297922 61218 297978
rect 61274 297922 61342 297978
rect 61398 297922 61494 297978
rect 60874 280350 61494 297922
rect 60874 280294 60970 280350
rect 61026 280294 61094 280350
rect 61150 280294 61218 280350
rect 61274 280294 61342 280350
rect 61398 280294 61494 280350
rect 60874 280226 61494 280294
rect 60874 280170 60970 280226
rect 61026 280170 61094 280226
rect 61150 280170 61218 280226
rect 61274 280170 61342 280226
rect 61398 280170 61494 280226
rect 60874 280102 61494 280170
rect 60874 280046 60970 280102
rect 61026 280046 61094 280102
rect 61150 280046 61218 280102
rect 61274 280046 61342 280102
rect 61398 280046 61494 280102
rect 60874 279978 61494 280046
rect 60874 279922 60970 279978
rect 61026 279922 61094 279978
rect 61150 279922 61218 279978
rect 61274 279922 61342 279978
rect 61398 279922 61494 279978
rect 60874 262350 61494 279922
rect 60874 262294 60970 262350
rect 61026 262294 61094 262350
rect 61150 262294 61218 262350
rect 61274 262294 61342 262350
rect 61398 262294 61494 262350
rect 60874 262226 61494 262294
rect 60874 262170 60970 262226
rect 61026 262170 61094 262226
rect 61150 262170 61218 262226
rect 61274 262170 61342 262226
rect 61398 262170 61494 262226
rect 60874 262102 61494 262170
rect 60874 262046 60970 262102
rect 61026 262046 61094 262102
rect 61150 262046 61218 262102
rect 61274 262046 61342 262102
rect 61398 262046 61494 262102
rect 60874 261978 61494 262046
rect 60874 261922 60970 261978
rect 61026 261922 61094 261978
rect 61150 261922 61218 261978
rect 61274 261922 61342 261978
rect 61398 261922 61494 261978
rect 60874 244350 61494 261922
rect 60874 244294 60970 244350
rect 61026 244294 61094 244350
rect 61150 244294 61218 244350
rect 61274 244294 61342 244350
rect 61398 244294 61494 244350
rect 60874 244226 61494 244294
rect 60874 244170 60970 244226
rect 61026 244170 61094 244226
rect 61150 244170 61218 244226
rect 61274 244170 61342 244226
rect 61398 244170 61494 244226
rect 60874 244102 61494 244170
rect 60874 244046 60970 244102
rect 61026 244046 61094 244102
rect 61150 244046 61218 244102
rect 61274 244046 61342 244102
rect 61398 244046 61494 244102
rect 60874 243978 61494 244046
rect 60874 243922 60970 243978
rect 61026 243922 61094 243978
rect 61150 243922 61218 243978
rect 61274 243922 61342 243978
rect 61398 243922 61494 243978
rect 60874 226350 61494 243922
rect 78874 586350 79494 597744
rect 78874 586294 78970 586350
rect 79026 586294 79094 586350
rect 79150 586294 79218 586350
rect 79274 586294 79342 586350
rect 79398 586294 79494 586350
rect 78874 586226 79494 586294
rect 78874 586170 78970 586226
rect 79026 586170 79094 586226
rect 79150 586170 79218 586226
rect 79274 586170 79342 586226
rect 79398 586170 79494 586226
rect 78874 586102 79494 586170
rect 78874 586046 78970 586102
rect 79026 586046 79094 586102
rect 79150 586046 79218 586102
rect 79274 586046 79342 586102
rect 79398 586046 79494 586102
rect 78874 585978 79494 586046
rect 78874 585922 78970 585978
rect 79026 585922 79094 585978
rect 79150 585922 79218 585978
rect 79274 585922 79342 585978
rect 79398 585922 79494 585978
rect 78874 568350 79494 585922
rect 78874 568294 78970 568350
rect 79026 568294 79094 568350
rect 79150 568294 79218 568350
rect 79274 568294 79342 568350
rect 79398 568294 79494 568350
rect 78874 568226 79494 568294
rect 78874 568170 78970 568226
rect 79026 568170 79094 568226
rect 79150 568170 79218 568226
rect 79274 568170 79342 568226
rect 79398 568170 79494 568226
rect 78874 568102 79494 568170
rect 78874 568046 78970 568102
rect 79026 568046 79094 568102
rect 79150 568046 79218 568102
rect 79274 568046 79342 568102
rect 79398 568046 79494 568102
rect 78874 567978 79494 568046
rect 78874 567922 78970 567978
rect 79026 567922 79094 567978
rect 79150 567922 79218 567978
rect 79274 567922 79342 567978
rect 79398 567922 79494 567978
rect 78874 550350 79494 567922
rect 78874 550294 78970 550350
rect 79026 550294 79094 550350
rect 79150 550294 79218 550350
rect 79274 550294 79342 550350
rect 79398 550294 79494 550350
rect 78874 550226 79494 550294
rect 78874 550170 78970 550226
rect 79026 550170 79094 550226
rect 79150 550170 79218 550226
rect 79274 550170 79342 550226
rect 79398 550170 79494 550226
rect 78874 550102 79494 550170
rect 78874 550046 78970 550102
rect 79026 550046 79094 550102
rect 79150 550046 79218 550102
rect 79274 550046 79342 550102
rect 79398 550046 79494 550102
rect 78874 549978 79494 550046
rect 78874 549922 78970 549978
rect 79026 549922 79094 549978
rect 79150 549922 79218 549978
rect 79274 549922 79342 549978
rect 79398 549922 79494 549978
rect 78874 532350 79494 549922
rect 78874 532294 78970 532350
rect 79026 532294 79094 532350
rect 79150 532294 79218 532350
rect 79274 532294 79342 532350
rect 79398 532294 79494 532350
rect 78874 532226 79494 532294
rect 78874 532170 78970 532226
rect 79026 532170 79094 532226
rect 79150 532170 79218 532226
rect 79274 532170 79342 532226
rect 79398 532170 79494 532226
rect 78874 532102 79494 532170
rect 78874 532046 78970 532102
rect 79026 532046 79094 532102
rect 79150 532046 79218 532102
rect 79274 532046 79342 532102
rect 79398 532046 79494 532102
rect 78874 531978 79494 532046
rect 78874 531922 78970 531978
rect 79026 531922 79094 531978
rect 79150 531922 79218 531978
rect 79274 531922 79342 531978
rect 79398 531922 79494 531978
rect 78874 514350 79494 531922
rect 78874 514294 78970 514350
rect 79026 514294 79094 514350
rect 79150 514294 79218 514350
rect 79274 514294 79342 514350
rect 79398 514294 79494 514350
rect 78874 514226 79494 514294
rect 78874 514170 78970 514226
rect 79026 514170 79094 514226
rect 79150 514170 79218 514226
rect 79274 514170 79342 514226
rect 79398 514170 79494 514226
rect 78874 514102 79494 514170
rect 78874 514046 78970 514102
rect 79026 514046 79094 514102
rect 79150 514046 79218 514102
rect 79274 514046 79342 514102
rect 79398 514046 79494 514102
rect 78874 513978 79494 514046
rect 78874 513922 78970 513978
rect 79026 513922 79094 513978
rect 79150 513922 79218 513978
rect 79274 513922 79342 513978
rect 79398 513922 79494 513978
rect 78874 496350 79494 513922
rect 78874 496294 78970 496350
rect 79026 496294 79094 496350
rect 79150 496294 79218 496350
rect 79274 496294 79342 496350
rect 79398 496294 79494 496350
rect 78874 496226 79494 496294
rect 78874 496170 78970 496226
rect 79026 496170 79094 496226
rect 79150 496170 79218 496226
rect 79274 496170 79342 496226
rect 79398 496170 79494 496226
rect 78874 496102 79494 496170
rect 78874 496046 78970 496102
rect 79026 496046 79094 496102
rect 79150 496046 79218 496102
rect 79274 496046 79342 496102
rect 79398 496046 79494 496102
rect 78874 495978 79494 496046
rect 78874 495922 78970 495978
rect 79026 495922 79094 495978
rect 79150 495922 79218 495978
rect 79274 495922 79342 495978
rect 79398 495922 79494 495978
rect 78874 478350 79494 495922
rect 78874 478294 78970 478350
rect 79026 478294 79094 478350
rect 79150 478294 79218 478350
rect 79274 478294 79342 478350
rect 79398 478294 79494 478350
rect 78874 478226 79494 478294
rect 78874 478170 78970 478226
rect 79026 478170 79094 478226
rect 79150 478170 79218 478226
rect 79274 478170 79342 478226
rect 79398 478170 79494 478226
rect 78874 478102 79494 478170
rect 78874 478046 78970 478102
rect 79026 478046 79094 478102
rect 79150 478046 79218 478102
rect 79274 478046 79342 478102
rect 79398 478046 79494 478102
rect 78874 477978 79494 478046
rect 78874 477922 78970 477978
rect 79026 477922 79094 477978
rect 79150 477922 79218 477978
rect 79274 477922 79342 477978
rect 79398 477922 79494 477978
rect 78874 460350 79494 477922
rect 78874 460294 78970 460350
rect 79026 460294 79094 460350
rect 79150 460294 79218 460350
rect 79274 460294 79342 460350
rect 79398 460294 79494 460350
rect 78874 460226 79494 460294
rect 78874 460170 78970 460226
rect 79026 460170 79094 460226
rect 79150 460170 79218 460226
rect 79274 460170 79342 460226
rect 79398 460170 79494 460226
rect 78874 460102 79494 460170
rect 78874 460046 78970 460102
rect 79026 460046 79094 460102
rect 79150 460046 79218 460102
rect 79274 460046 79342 460102
rect 79398 460046 79494 460102
rect 78874 459978 79494 460046
rect 78874 459922 78970 459978
rect 79026 459922 79094 459978
rect 79150 459922 79218 459978
rect 79274 459922 79342 459978
rect 79398 459922 79494 459978
rect 78874 442350 79494 459922
rect 78874 442294 78970 442350
rect 79026 442294 79094 442350
rect 79150 442294 79218 442350
rect 79274 442294 79342 442350
rect 79398 442294 79494 442350
rect 78874 442226 79494 442294
rect 78874 442170 78970 442226
rect 79026 442170 79094 442226
rect 79150 442170 79218 442226
rect 79274 442170 79342 442226
rect 79398 442170 79494 442226
rect 78874 442102 79494 442170
rect 78874 442046 78970 442102
rect 79026 442046 79094 442102
rect 79150 442046 79218 442102
rect 79274 442046 79342 442102
rect 79398 442046 79494 442102
rect 78874 441978 79494 442046
rect 78874 441922 78970 441978
rect 79026 441922 79094 441978
rect 79150 441922 79218 441978
rect 79274 441922 79342 441978
rect 79398 441922 79494 441978
rect 78874 424350 79494 441922
rect 78874 424294 78970 424350
rect 79026 424294 79094 424350
rect 79150 424294 79218 424350
rect 79274 424294 79342 424350
rect 79398 424294 79494 424350
rect 78874 424226 79494 424294
rect 78874 424170 78970 424226
rect 79026 424170 79094 424226
rect 79150 424170 79218 424226
rect 79274 424170 79342 424226
rect 79398 424170 79494 424226
rect 78874 424102 79494 424170
rect 78874 424046 78970 424102
rect 79026 424046 79094 424102
rect 79150 424046 79218 424102
rect 79274 424046 79342 424102
rect 79398 424046 79494 424102
rect 78874 423978 79494 424046
rect 78874 423922 78970 423978
rect 79026 423922 79094 423978
rect 79150 423922 79218 423978
rect 79274 423922 79342 423978
rect 79398 423922 79494 423978
rect 78874 406350 79494 423922
rect 78874 406294 78970 406350
rect 79026 406294 79094 406350
rect 79150 406294 79218 406350
rect 79274 406294 79342 406350
rect 79398 406294 79494 406350
rect 78874 406226 79494 406294
rect 78874 406170 78970 406226
rect 79026 406170 79094 406226
rect 79150 406170 79218 406226
rect 79274 406170 79342 406226
rect 79398 406170 79494 406226
rect 78874 406102 79494 406170
rect 78874 406046 78970 406102
rect 79026 406046 79094 406102
rect 79150 406046 79218 406102
rect 79274 406046 79342 406102
rect 79398 406046 79494 406102
rect 78874 405978 79494 406046
rect 78874 405922 78970 405978
rect 79026 405922 79094 405978
rect 79150 405922 79218 405978
rect 79274 405922 79342 405978
rect 79398 405922 79494 405978
rect 78874 388350 79494 405922
rect 78874 388294 78970 388350
rect 79026 388294 79094 388350
rect 79150 388294 79218 388350
rect 79274 388294 79342 388350
rect 79398 388294 79494 388350
rect 78874 388226 79494 388294
rect 78874 388170 78970 388226
rect 79026 388170 79094 388226
rect 79150 388170 79218 388226
rect 79274 388170 79342 388226
rect 79398 388170 79494 388226
rect 78874 388102 79494 388170
rect 78874 388046 78970 388102
rect 79026 388046 79094 388102
rect 79150 388046 79218 388102
rect 79274 388046 79342 388102
rect 79398 388046 79494 388102
rect 78874 387978 79494 388046
rect 78874 387922 78970 387978
rect 79026 387922 79094 387978
rect 79150 387922 79218 387978
rect 79274 387922 79342 387978
rect 79398 387922 79494 387978
rect 78874 370350 79494 387922
rect 78874 370294 78970 370350
rect 79026 370294 79094 370350
rect 79150 370294 79218 370350
rect 79274 370294 79342 370350
rect 79398 370294 79494 370350
rect 78874 370226 79494 370294
rect 78874 370170 78970 370226
rect 79026 370170 79094 370226
rect 79150 370170 79218 370226
rect 79274 370170 79342 370226
rect 79398 370170 79494 370226
rect 78874 370102 79494 370170
rect 78874 370046 78970 370102
rect 79026 370046 79094 370102
rect 79150 370046 79218 370102
rect 79274 370046 79342 370102
rect 79398 370046 79494 370102
rect 78874 369978 79494 370046
rect 78874 369922 78970 369978
rect 79026 369922 79094 369978
rect 79150 369922 79218 369978
rect 79274 369922 79342 369978
rect 79398 369922 79494 369978
rect 78874 352350 79494 369922
rect 78874 352294 78970 352350
rect 79026 352294 79094 352350
rect 79150 352294 79218 352350
rect 79274 352294 79342 352350
rect 79398 352294 79494 352350
rect 78874 352226 79494 352294
rect 78874 352170 78970 352226
rect 79026 352170 79094 352226
rect 79150 352170 79218 352226
rect 79274 352170 79342 352226
rect 79398 352170 79494 352226
rect 78874 352102 79494 352170
rect 78874 352046 78970 352102
rect 79026 352046 79094 352102
rect 79150 352046 79218 352102
rect 79274 352046 79342 352102
rect 79398 352046 79494 352102
rect 78874 351978 79494 352046
rect 78874 351922 78970 351978
rect 79026 351922 79094 351978
rect 79150 351922 79218 351978
rect 79274 351922 79342 351978
rect 79398 351922 79494 351978
rect 78874 334350 79494 351922
rect 78874 334294 78970 334350
rect 79026 334294 79094 334350
rect 79150 334294 79218 334350
rect 79274 334294 79342 334350
rect 79398 334294 79494 334350
rect 78874 334226 79494 334294
rect 78874 334170 78970 334226
rect 79026 334170 79094 334226
rect 79150 334170 79218 334226
rect 79274 334170 79342 334226
rect 79398 334170 79494 334226
rect 78874 334102 79494 334170
rect 78874 334046 78970 334102
rect 79026 334046 79094 334102
rect 79150 334046 79218 334102
rect 79274 334046 79342 334102
rect 79398 334046 79494 334102
rect 78874 333978 79494 334046
rect 78874 333922 78970 333978
rect 79026 333922 79094 333978
rect 79150 333922 79218 333978
rect 79274 333922 79342 333978
rect 79398 333922 79494 333978
rect 78874 316350 79494 333922
rect 78874 316294 78970 316350
rect 79026 316294 79094 316350
rect 79150 316294 79218 316350
rect 79274 316294 79342 316350
rect 79398 316294 79494 316350
rect 78874 316226 79494 316294
rect 78874 316170 78970 316226
rect 79026 316170 79094 316226
rect 79150 316170 79218 316226
rect 79274 316170 79342 316226
rect 79398 316170 79494 316226
rect 78874 316102 79494 316170
rect 78874 316046 78970 316102
rect 79026 316046 79094 316102
rect 79150 316046 79218 316102
rect 79274 316046 79342 316102
rect 79398 316046 79494 316102
rect 78874 315978 79494 316046
rect 78874 315922 78970 315978
rect 79026 315922 79094 315978
rect 79150 315922 79218 315978
rect 79274 315922 79342 315978
rect 79398 315922 79494 315978
rect 78874 298350 79494 315922
rect 78874 298294 78970 298350
rect 79026 298294 79094 298350
rect 79150 298294 79218 298350
rect 79274 298294 79342 298350
rect 79398 298294 79494 298350
rect 78874 298226 79494 298294
rect 78874 298170 78970 298226
rect 79026 298170 79094 298226
rect 79150 298170 79218 298226
rect 79274 298170 79342 298226
rect 79398 298170 79494 298226
rect 78874 298102 79494 298170
rect 78874 298046 78970 298102
rect 79026 298046 79094 298102
rect 79150 298046 79218 298102
rect 79274 298046 79342 298102
rect 79398 298046 79494 298102
rect 78874 297978 79494 298046
rect 78874 297922 78970 297978
rect 79026 297922 79094 297978
rect 79150 297922 79218 297978
rect 79274 297922 79342 297978
rect 79398 297922 79494 297978
rect 78874 280350 79494 297922
rect 78874 280294 78970 280350
rect 79026 280294 79094 280350
rect 79150 280294 79218 280350
rect 79274 280294 79342 280350
rect 79398 280294 79494 280350
rect 78874 280226 79494 280294
rect 78874 280170 78970 280226
rect 79026 280170 79094 280226
rect 79150 280170 79218 280226
rect 79274 280170 79342 280226
rect 79398 280170 79494 280226
rect 78874 280102 79494 280170
rect 78874 280046 78970 280102
rect 79026 280046 79094 280102
rect 79150 280046 79218 280102
rect 79274 280046 79342 280102
rect 79398 280046 79494 280102
rect 78874 279978 79494 280046
rect 78874 279922 78970 279978
rect 79026 279922 79094 279978
rect 79150 279922 79218 279978
rect 79274 279922 79342 279978
rect 79398 279922 79494 279978
rect 78874 262350 79494 279922
rect 78874 262294 78970 262350
rect 79026 262294 79094 262350
rect 79150 262294 79218 262350
rect 79274 262294 79342 262350
rect 79398 262294 79494 262350
rect 78874 262226 79494 262294
rect 78874 262170 78970 262226
rect 79026 262170 79094 262226
rect 79150 262170 79218 262226
rect 79274 262170 79342 262226
rect 79398 262170 79494 262226
rect 78874 262102 79494 262170
rect 78874 262046 78970 262102
rect 79026 262046 79094 262102
rect 79150 262046 79218 262102
rect 79274 262046 79342 262102
rect 79398 262046 79494 262102
rect 78874 261978 79494 262046
rect 78874 261922 78970 261978
rect 79026 261922 79094 261978
rect 79150 261922 79218 261978
rect 79274 261922 79342 261978
rect 79398 261922 79494 261978
rect 78874 244350 79494 261922
rect 78874 244294 78970 244350
rect 79026 244294 79094 244350
rect 79150 244294 79218 244350
rect 79274 244294 79342 244350
rect 79398 244294 79494 244350
rect 78874 244226 79494 244294
rect 78874 244170 78970 244226
rect 79026 244170 79094 244226
rect 79150 244170 79218 244226
rect 79274 244170 79342 244226
rect 79398 244170 79494 244226
rect 78874 244102 79494 244170
rect 78874 244046 78970 244102
rect 79026 244046 79094 244102
rect 79150 244046 79218 244102
rect 79274 244046 79342 244102
rect 79398 244046 79494 244102
rect 78874 243978 79494 244046
rect 78874 243922 78970 243978
rect 79026 243922 79094 243978
rect 79150 243922 79218 243978
rect 79274 243922 79342 243978
rect 79398 243922 79494 243978
rect 75154 238350 75774 242964
rect 75154 238294 75250 238350
rect 75306 238294 75374 238350
rect 75430 238294 75498 238350
rect 75554 238294 75622 238350
rect 75678 238294 75774 238350
rect 75154 238226 75774 238294
rect 75154 238170 75250 238226
rect 75306 238170 75374 238226
rect 75430 238170 75498 238226
rect 75554 238170 75622 238226
rect 75678 238170 75774 238226
rect 75154 238102 75774 238170
rect 75154 238046 75250 238102
rect 75306 238046 75374 238102
rect 75430 238046 75498 238102
rect 75554 238046 75622 238102
rect 75678 238046 75774 238102
rect 75154 237978 75774 238046
rect 75154 237922 75250 237978
rect 75306 237922 75374 237978
rect 75430 237922 75498 237978
rect 75554 237922 75622 237978
rect 75678 237922 75774 237978
rect 63868 229348 63924 229358
rect 63868 227668 63924 229292
rect 63868 227602 63924 227612
rect 60874 226294 60970 226350
rect 61026 226294 61094 226350
rect 61150 226294 61218 226350
rect 61274 226294 61342 226350
rect 61398 226294 61494 226350
rect 60874 226226 61494 226294
rect 60874 226170 60970 226226
rect 61026 226170 61094 226226
rect 61150 226170 61218 226226
rect 61274 226170 61342 226226
rect 61398 226170 61494 226226
rect 60874 226102 61494 226170
rect 60874 226046 60970 226102
rect 61026 226046 61094 226102
rect 61150 226046 61218 226102
rect 61274 226046 61342 226102
rect 61398 226046 61494 226102
rect 60874 225978 61494 226046
rect 60874 225922 60970 225978
rect 61026 225922 61094 225978
rect 61150 225922 61218 225978
rect 61274 225922 61342 225978
rect 61398 225922 61494 225978
rect 60874 219134 61494 225922
rect 64448 220350 64768 220384
rect 64448 220294 64518 220350
rect 64574 220294 64642 220350
rect 64698 220294 64768 220350
rect 64448 220226 64768 220294
rect 64448 220170 64518 220226
rect 64574 220170 64642 220226
rect 64698 220170 64768 220226
rect 64448 220102 64768 220170
rect 64448 220046 64518 220102
rect 64574 220046 64642 220102
rect 64698 220046 64768 220102
rect 64448 219978 64768 220046
rect 64448 219922 64518 219978
rect 64574 219922 64642 219978
rect 64698 219922 64768 219978
rect 64448 219888 64768 219922
rect 75154 220350 75774 237922
rect 75154 220294 75250 220350
rect 75306 220294 75374 220350
rect 75430 220294 75498 220350
rect 75554 220294 75622 220350
rect 75678 220294 75774 220350
rect 75154 220226 75774 220294
rect 75154 220170 75250 220226
rect 75306 220170 75374 220226
rect 75430 220170 75498 220226
rect 75554 220170 75622 220226
rect 75678 220170 75774 220226
rect 75154 220102 75774 220170
rect 75154 220046 75250 220102
rect 75306 220046 75374 220102
rect 75430 220046 75498 220102
rect 75554 220046 75622 220102
rect 75678 220046 75774 220102
rect 75154 219978 75774 220046
rect 75154 219922 75250 219978
rect 75306 219922 75374 219978
rect 75430 219922 75498 219978
rect 75554 219922 75622 219978
rect 75678 219922 75774 219978
rect 75154 219134 75774 219922
rect 78874 226350 79494 243922
rect 93154 597212 93774 598268
rect 93154 597156 93250 597212
rect 93306 597156 93374 597212
rect 93430 597156 93498 597212
rect 93554 597156 93622 597212
rect 93678 597156 93774 597212
rect 93154 597088 93774 597156
rect 93154 597032 93250 597088
rect 93306 597032 93374 597088
rect 93430 597032 93498 597088
rect 93554 597032 93622 597088
rect 93678 597032 93774 597088
rect 93154 596964 93774 597032
rect 93154 596908 93250 596964
rect 93306 596908 93374 596964
rect 93430 596908 93498 596964
rect 93554 596908 93622 596964
rect 93678 596908 93774 596964
rect 93154 596840 93774 596908
rect 93154 596784 93250 596840
rect 93306 596784 93374 596840
rect 93430 596784 93498 596840
rect 93554 596784 93622 596840
rect 93678 596784 93774 596840
rect 93154 580350 93774 596784
rect 93154 580294 93250 580350
rect 93306 580294 93374 580350
rect 93430 580294 93498 580350
rect 93554 580294 93622 580350
rect 93678 580294 93774 580350
rect 93154 580226 93774 580294
rect 93154 580170 93250 580226
rect 93306 580170 93374 580226
rect 93430 580170 93498 580226
rect 93554 580170 93622 580226
rect 93678 580170 93774 580226
rect 93154 580102 93774 580170
rect 93154 580046 93250 580102
rect 93306 580046 93374 580102
rect 93430 580046 93498 580102
rect 93554 580046 93622 580102
rect 93678 580046 93774 580102
rect 93154 579978 93774 580046
rect 93154 579922 93250 579978
rect 93306 579922 93374 579978
rect 93430 579922 93498 579978
rect 93554 579922 93622 579978
rect 93678 579922 93774 579978
rect 93154 562350 93774 579922
rect 93154 562294 93250 562350
rect 93306 562294 93374 562350
rect 93430 562294 93498 562350
rect 93554 562294 93622 562350
rect 93678 562294 93774 562350
rect 93154 562226 93774 562294
rect 93154 562170 93250 562226
rect 93306 562170 93374 562226
rect 93430 562170 93498 562226
rect 93554 562170 93622 562226
rect 93678 562170 93774 562226
rect 93154 562102 93774 562170
rect 93154 562046 93250 562102
rect 93306 562046 93374 562102
rect 93430 562046 93498 562102
rect 93554 562046 93622 562102
rect 93678 562046 93774 562102
rect 93154 561978 93774 562046
rect 93154 561922 93250 561978
rect 93306 561922 93374 561978
rect 93430 561922 93498 561978
rect 93554 561922 93622 561978
rect 93678 561922 93774 561978
rect 93154 544350 93774 561922
rect 93154 544294 93250 544350
rect 93306 544294 93374 544350
rect 93430 544294 93498 544350
rect 93554 544294 93622 544350
rect 93678 544294 93774 544350
rect 93154 544226 93774 544294
rect 93154 544170 93250 544226
rect 93306 544170 93374 544226
rect 93430 544170 93498 544226
rect 93554 544170 93622 544226
rect 93678 544170 93774 544226
rect 93154 544102 93774 544170
rect 93154 544046 93250 544102
rect 93306 544046 93374 544102
rect 93430 544046 93498 544102
rect 93554 544046 93622 544102
rect 93678 544046 93774 544102
rect 93154 543978 93774 544046
rect 93154 543922 93250 543978
rect 93306 543922 93374 543978
rect 93430 543922 93498 543978
rect 93554 543922 93622 543978
rect 93678 543922 93774 543978
rect 93154 526350 93774 543922
rect 93154 526294 93250 526350
rect 93306 526294 93374 526350
rect 93430 526294 93498 526350
rect 93554 526294 93622 526350
rect 93678 526294 93774 526350
rect 93154 526226 93774 526294
rect 93154 526170 93250 526226
rect 93306 526170 93374 526226
rect 93430 526170 93498 526226
rect 93554 526170 93622 526226
rect 93678 526170 93774 526226
rect 93154 526102 93774 526170
rect 93154 526046 93250 526102
rect 93306 526046 93374 526102
rect 93430 526046 93498 526102
rect 93554 526046 93622 526102
rect 93678 526046 93774 526102
rect 93154 525978 93774 526046
rect 93154 525922 93250 525978
rect 93306 525922 93374 525978
rect 93430 525922 93498 525978
rect 93554 525922 93622 525978
rect 93678 525922 93774 525978
rect 93154 508350 93774 525922
rect 93154 508294 93250 508350
rect 93306 508294 93374 508350
rect 93430 508294 93498 508350
rect 93554 508294 93622 508350
rect 93678 508294 93774 508350
rect 93154 508226 93774 508294
rect 93154 508170 93250 508226
rect 93306 508170 93374 508226
rect 93430 508170 93498 508226
rect 93554 508170 93622 508226
rect 93678 508170 93774 508226
rect 93154 508102 93774 508170
rect 93154 508046 93250 508102
rect 93306 508046 93374 508102
rect 93430 508046 93498 508102
rect 93554 508046 93622 508102
rect 93678 508046 93774 508102
rect 93154 507978 93774 508046
rect 93154 507922 93250 507978
rect 93306 507922 93374 507978
rect 93430 507922 93498 507978
rect 93554 507922 93622 507978
rect 93678 507922 93774 507978
rect 93154 490350 93774 507922
rect 93154 490294 93250 490350
rect 93306 490294 93374 490350
rect 93430 490294 93498 490350
rect 93554 490294 93622 490350
rect 93678 490294 93774 490350
rect 93154 490226 93774 490294
rect 93154 490170 93250 490226
rect 93306 490170 93374 490226
rect 93430 490170 93498 490226
rect 93554 490170 93622 490226
rect 93678 490170 93774 490226
rect 93154 490102 93774 490170
rect 93154 490046 93250 490102
rect 93306 490046 93374 490102
rect 93430 490046 93498 490102
rect 93554 490046 93622 490102
rect 93678 490046 93774 490102
rect 93154 489978 93774 490046
rect 93154 489922 93250 489978
rect 93306 489922 93374 489978
rect 93430 489922 93498 489978
rect 93554 489922 93622 489978
rect 93678 489922 93774 489978
rect 93154 472350 93774 489922
rect 93154 472294 93250 472350
rect 93306 472294 93374 472350
rect 93430 472294 93498 472350
rect 93554 472294 93622 472350
rect 93678 472294 93774 472350
rect 93154 472226 93774 472294
rect 93154 472170 93250 472226
rect 93306 472170 93374 472226
rect 93430 472170 93498 472226
rect 93554 472170 93622 472226
rect 93678 472170 93774 472226
rect 93154 472102 93774 472170
rect 93154 472046 93250 472102
rect 93306 472046 93374 472102
rect 93430 472046 93498 472102
rect 93554 472046 93622 472102
rect 93678 472046 93774 472102
rect 93154 471978 93774 472046
rect 93154 471922 93250 471978
rect 93306 471922 93374 471978
rect 93430 471922 93498 471978
rect 93554 471922 93622 471978
rect 93678 471922 93774 471978
rect 93154 454350 93774 471922
rect 93154 454294 93250 454350
rect 93306 454294 93374 454350
rect 93430 454294 93498 454350
rect 93554 454294 93622 454350
rect 93678 454294 93774 454350
rect 93154 454226 93774 454294
rect 93154 454170 93250 454226
rect 93306 454170 93374 454226
rect 93430 454170 93498 454226
rect 93554 454170 93622 454226
rect 93678 454170 93774 454226
rect 93154 454102 93774 454170
rect 93154 454046 93250 454102
rect 93306 454046 93374 454102
rect 93430 454046 93498 454102
rect 93554 454046 93622 454102
rect 93678 454046 93774 454102
rect 93154 453978 93774 454046
rect 93154 453922 93250 453978
rect 93306 453922 93374 453978
rect 93430 453922 93498 453978
rect 93554 453922 93622 453978
rect 93678 453922 93774 453978
rect 93154 436350 93774 453922
rect 93154 436294 93250 436350
rect 93306 436294 93374 436350
rect 93430 436294 93498 436350
rect 93554 436294 93622 436350
rect 93678 436294 93774 436350
rect 93154 436226 93774 436294
rect 93154 436170 93250 436226
rect 93306 436170 93374 436226
rect 93430 436170 93498 436226
rect 93554 436170 93622 436226
rect 93678 436170 93774 436226
rect 93154 436102 93774 436170
rect 93154 436046 93250 436102
rect 93306 436046 93374 436102
rect 93430 436046 93498 436102
rect 93554 436046 93622 436102
rect 93678 436046 93774 436102
rect 93154 435978 93774 436046
rect 93154 435922 93250 435978
rect 93306 435922 93374 435978
rect 93430 435922 93498 435978
rect 93554 435922 93622 435978
rect 93678 435922 93774 435978
rect 93154 418350 93774 435922
rect 93154 418294 93250 418350
rect 93306 418294 93374 418350
rect 93430 418294 93498 418350
rect 93554 418294 93622 418350
rect 93678 418294 93774 418350
rect 93154 418226 93774 418294
rect 93154 418170 93250 418226
rect 93306 418170 93374 418226
rect 93430 418170 93498 418226
rect 93554 418170 93622 418226
rect 93678 418170 93774 418226
rect 93154 418102 93774 418170
rect 93154 418046 93250 418102
rect 93306 418046 93374 418102
rect 93430 418046 93498 418102
rect 93554 418046 93622 418102
rect 93678 418046 93774 418102
rect 93154 417978 93774 418046
rect 93154 417922 93250 417978
rect 93306 417922 93374 417978
rect 93430 417922 93498 417978
rect 93554 417922 93622 417978
rect 93678 417922 93774 417978
rect 93154 400350 93774 417922
rect 93154 400294 93250 400350
rect 93306 400294 93374 400350
rect 93430 400294 93498 400350
rect 93554 400294 93622 400350
rect 93678 400294 93774 400350
rect 93154 400226 93774 400294
rect 93154 400170 93250 400226
rect 93306 400170 93374 400226
rect 93430 400170 93498 400226
rect 93554 400170 93622 400226
rect 93678 400170 93774 400226
rect 93154 400102 93774 400170
rect 93154 400046 93250 400102
rect 93306 400046 93374 400102
rect 93430 400046 93498 400102
rect 93554 400046 93622 400102
rect 93678 400046 93774 400102
rect 93154 399978 93774 400046
rect 93154 399922 93250 399978
rect 93306 399922 93374 399978
rect 93430 399922 93498 399978
rect 93554 399922 93622 399978
rect 93678 399922 93774 399978
rect 93154 382350 93774 399922
rect 93154 382294 93250 382350
rect 93306 382294 93374 382350
rect 93430 382294 93498 382350
rect 93554 382294 93622 382350
rect 93678 382294 93774 382350
rect 93154 382226 93774 382294
rect 93154 382170 93250 382226
rect 93306 382170 93374 382226
rect 93430 382170 93498 382226
rect 93554 382170 93622 382226
rect 93678 382170 93774 382226
rect 93154 382102 93774 382170
rect 93154 382046 93250 382102
rect 93306 382046 93374 382102
rect 93430 382046 93498 382102
rect 93554 382046 93622 382102
rect 93678 382046 93774 382102
rect 93154 381978 93774 382046
rect 93154 381922 93250 381978
rect 93306 381922 93374 381978
rect 93430 381922 93498 381978
rect 93554 381922 93622 381978
rect 93678 381922 93774 381978
rect 93154 364350 93774 381922
rect 93154 364294 93250 364350
rect 93306 364294 93374 364350
rect 93430 364294 93498 364350
rect 93554 364294 93622 364350
rect 93678 364294 93774 364350
rect 93154 364226 93774 364294
rect 93154 364170 93250 364226
rect 93306 364170 93374 364226
rect 93430 364170 93498 364226
rect 93554 364170 93622 364226
rect 93678 364170 93774 364226
rect 93154 364102 93774 364170
rect 93154 364046 93250 364102
rect 93306 364046 93374 364102
rect 93430 364046 93498 364102
rect 93554 364046 93622 364102
rect 93678 364046 93774 364102
rect 93154 363978 93774 364046
rect 93154 363922 93250 363978
rect 93306 363922 93374 363978
rect 93430 363922 93498 363978
rect 93554 363922 93622 363978
rect 93678 363922 93774 363978
rect 93154 346350 93774 363922
rect 93154 346294 93250 346350
rect 93306 346294 93374 346350
rect 93430 346294 93498 346350
rect 93554 346294 93622 346350
rect 93678 346294 93774 346350
rect 93154 346226 93774 346294
rect 93154 346170 93250 346226
rect 93306 346170 93374 346226
rect 93430 346170 93498 346226
rect 93554 346170 93622 346226
rect 93678 346170 93774 346226
rect 93154 346102 93774 346170
rect 93154 346046 93250 346102
rect 93306 346046 93374 346102
rect 93430 346046 93498 346102
rect 93554 346046 93622 346102
rect 93678 346046 93774 346102
rect 93154 345978 93774 346046
rect 93154 345922 93250 345978
rect 93306 345922 93374 345978
rect 93430 345922 93498 345978
rect 93554 345922 93622 345978
rect 93678 345922 93774 345978
rect 93154 328350 93774 345922
rect 93154 328294 93250 328350
rect 93306 328294 93374 328350
rect 93430 328294 93498 328350
rect 93554 328294 93622 328350
rect 93678 328294 93774 328350
rect 93154 328226 93774 328294
rect 93154 328170 93250 328226
rect 93306 328170 93374 328226
rect 93430 328170 93498 328226
rect 93554 328170 93622 328226
rect 93678 328170 93774 328226
rect 93154 328102 93774 328170
rect 93154 328046 93250 328102
rect 93306 328046 93374 328102
rect 93430 328046 93498 328102
rect 93554 328046 93622 328102
rect 93678 328046 93774 328102
rect 93154 327978 93774 328046
rect 93154 327922 93250 327978
rect 93306 327922 93374 327978
rect 93430 327922 93498 327978
rect 93554 327922 93622 327978
rect 93678 327922 93774 327978
rect 93154 310350 93774 327922
rect 93154 310294 93250 310350
rect 93306 310294 93374 310350
rect 93430 310294 93498 310350
rect 93554 310294 93622 310350
rect 93678 310294 93774 310350
rect 93154 310226 93774 310294
rect 93154 310170 93250 310226
rect 93306 310170 93374 310226
rect 93430 310170 93498 310226
rect 93554 310170 93622 310226
rect 93678 310170 93774 310226
rect 93154 310102 93774 310170
rect 93154 310046 93250 310102
rect 93306 310046 93374 310102
rect 93430 310046 93498 310102
rect 93554 310046 93622 310102
rect 93678 310046 93774 310102
rect 93154 309978 93774 310046
rect 93154 309922 93250 309978
rect 93306 309922 93374 309978
rect 93430 309922 93498 309978
rect 93554 309922 93622 309978
rect 93678 309922 93774 309978
rect 93154 292350 93774 309922
rect 93154 292294 93250 292350
rect 93306 292294 93374 292350
rect 93430 292294 93498 292350
rect 93554 292294 93622 292350
rect 93678 292294 93774 292350
rect 93154 292226 93774 292294
rect 93154 292170 93250 292226
rect 93306 292170 93374 292226
rect 93430 292170 93498 292226
rect 93554 292170 93622 292226
rect 93678 292170 93774 292226
rect 93154 292102 93774 292170
rect 93154 292046 93250 292102
rect 93306 292046 93374 292102
rect 93430 292046 93498 292102
rect 93554 292046 93622 292102
rect 93678 292046 93774 292102
rect 93154 291978 93774 292046
rect 93154 291922 93250 291978
rect 93306 291922 93374 291978
rect 93430 291922 93498 291978
rect 93554 291922 93622 291978
rect 93678 291922 93774 291978
rect 93154 274350 93774 291922
rect 93154 274294 93250 274350
rect 93306 274294 93374 274350
rect 93430 274294 93498 274350
rect 93554 274294 93622 274350
rect 93678 274294 93774 274350
rect 93154 274226 93774 274294
rect 93154 274170 93250 274226
rect 93306 274170 93374 274226
rect 93430 274170 93498 274226
rect 93554 274170 93622 274226
rect 93678 274170 93774 274226
rect 93154 274102 93774 274170
rect 93154 274046 93250 274102
rect 93306 274046 93374 274102
rect 93430 274046 93498 274102
rect 93554 274046 93622 274102
rect 93678 274046 93774 274102
rect 93154 273978 93774 274046
rect 93154 273922 93250 273978
rect 93306 273922 93374 273978
rect 93430 273922 93498 273978
rect 93554 273922 93622 273978
rect 93678 273922 93774 273978
rect 93154 256350 93774 273922
rect 93154 256294 93250 256350
rect 93306 256294 93374 256350
rect 93430 256294 93498 256350
rect 93554 256294 93622 256350
rect 93678 256294 93774 256350
rect 93154 256226 93774 256294
rect 93154 256170 93250 256226
rect 93306 256170 93374 256226
rect 93430 256170 93498 256226
rect 93554 256170 93622 256226
rect 93678 256170 93774 256226
rect 93154 256102 93774 256170
rect 93154 256046 93250 256102
rect 93306 256046 93374 256102
rect 93430 256046 93498 256102
rect 93554 256046 93622 256102
rect 93678 256046 93774 256102
rect 93154 255978 93774 256046
rect 93154 255922 93250 255978
rect 93306 255922 93374 255978
rect 93430 255922 93498 255978
rect 93554 255922 93622 255978
rect 93678 255922 93774 255978
rect 93154 238350 93774 255922
rect 93154 238294 93250 238350
rect 93306 238294 93374 238350
rect 93430 238294 93498 238350
rect 93554 238294 93622 238350
rect 93678 238294 93774 238350
rect 93154 238226 93774 238294
rect 93154 238170 93250 238226
rect 93306 238170 93374 238226
rect 93430 238170 93498 238226
rect 93554 238170 93622 238226
rect 93678 238170 93774 238226
rect 93154 238102 93774 238170
rect 93154 238046 93250 238102
rect 93306 238046 93374 238102
rect 93430 238046 93498 238102
rect 93554 238046 93622 238102
rect 93678 238046 93774 238102
rect 93154 237978 93774 238046
rect 93154 237922 93250 237978
rect 93306 237922 93374 237978
rect 93430 237922 93498 237978
rect 93554 237922 93622 237978
rect 93678 237922 93774 237978
rect 80892 229460 80948 229470
rect 80892 227892 80948 229404
rect 80892 227826 80948 227836
rect 78874 226294 78970 226350
rect 79026 226294 79094 226350
rect 79150 226294 79218 226350
rect 79274 226294 79342 226350
rect 79398 226294 79494 226350
rect 78874 226226 79494 226294
rect 78874 226170 78970 226226
rect 79026 226170 79094 226226
rect 79150 226170 79218 226226
rect 79274 226170 79342 226226
rect 79398 226170 79494 226226
rect 78874 226102 79494 226170
rect 78874 226046 78970 226102
rect 79026 226046 79094 226102
rect 79150 226046 79218 226102
rect 79274 226046 79342 226102
rect 79398 226046 79494 226102
rect 78874 225978 79494 226046
rect 78874 225922 78970 225978
rect 79026 225922 79094 225978
rect 79150 225922 79218 225978
rect 79274 225922 79342 225978
rect 79398 225922 79494 225978
rect 78874 219134 79494 225922
rect 79808 226350 80128 226384
rect 79808 226294 79878 226350
rect 79934 226294 80002 226350
rect 80058 226294 80128 226350
rect 79808 226226 80128 226294
rect 79808 226170 79878 226226
rect 79934 226170 80002 226226
rect 80058 226170 80128 226226
rect 79808 226102 80128 226170
rect 79808 226046 79878 226102
rect 79934 226046 80002 226102
rect 80058 226046 80128 226102
rect 79808 225978 80128 226046
rect 79808 225922 79878 225978
rect 79934 225922 80002 225978
rect 80058 225922 80128 225978
rect 79808 225888 80128 225922
rect 93154 220350 93774 237922
rect 96874 598172 97494 598268
rect 96874 598116 96970 598172
rect 97026 598116 97094 598172
rect 97150 598116 97218 598172
rect 97274 598116 97342 598172
rect 97398 598116 97494 598172
rect 96874 598048 97494 598116
rect 96874 597992 96970 598048
rect 97026 597992 97094 598048
rect 97150 597992 97218 598048
rect 97274 597992 97342 598048
rect 97398 597992 97494 598048
rect 96874 597924 97494 597992
rect 96874 597868 96970 597924
rect 97026 597868 97094 597924
rect 97150 597868 97218 597924
rect 97274 597868 97342 597924
rect 97398 597868 97494 597924
rect 96874 597800 97494 597868
rect 96874 597744 96970 597800
rect 97026 597744 97094 597800
rect 97150 597744 97218 597800
rect 97274 597744 97342 597800
rect 97398 597744 97494 597800
rect 96874 586350 97494 597744
rect 96874 586294 96970 586350
rect 97026 586294 97094 586350
rect 97150 586294 97218 586350
rect 97274 586294 97342 586350
rect 97398 586294 97494 586350
rect 96874 586226 97494 586294
rect 96874 586170 96970 586226
rect 97026 586170 97094 586226
rect 97150 586170 97218 586226
rect 97274 586170 97342 586226
rect 97398 586170 97494 586226
rect 96874 586102 97494 586170
rect 96874 586046 96970 586102
rect 97026 586046 97094 586102
rect 97150 586046 97218 586102
rect 97274 586046 97342 586102
rect 97398 586046 97494 586102
rect 96874 585978 97494 586046
rect 96874 585922 96970 585978
rect 97026 585922 97094 585978
rect 97150 585922 97218 585978
rect 97274 585922 97342 585978
rect 97398 585922 97494 585978
rect 96874 568350 97494 585922
rect 96874 568294 96970 568350
rect 97026 568294 97094 568350
rect 97150 568294 97218 568350
rect 97274 568294 97342 568350
rect 97398 568294 97494 568350
rect 96874 568226 97494 568294
rect 96874 568170 96970 568226
rect 97026 568170 97094 568226
rect 97150 568170 97218 568226
rect 97274 568170 97342 568226
rect 97398 568170 97494 568226
rect 96874 568102 97494 568170
rect 96874 568046 96970 568102
rect 97026 568046 97094 568102
rect 97150 568046 97218 568102
rect 97274 568046 97342 568102
rect 97398 568046 97494 568102
rect 96874 567978 97494 568046
rect 96874 567922 96970 567978
rect 97026 567922 97094 567978
rect 97150 567922 97218 567978
rect 97274 567922 97342 567978
rect 97398 567922 97494 567978
rect 96874 550350 97494 567922
rect 96874 550294 96970 550350
rect 97026 550294 97094 550350
rect 97150 550294 97218 550350
rect 97274 550294 97342 550350
rect 97398 550294 97494 550350
rect 96874 550226 97494 550294
rect 96874 550170 96970 550226
rect 97026 550170 97094 550226
rect 97150 550170 97218 550226
rect 97274 550170 97342 550226
rect 97398 550170 97494 550226
rect 96874 550102 97494 550170
rect 96874 550046 96970 550102
rect 97026 550046 97094 550102
rect 97150 550046 97218 550102
rect 97274 550046 97342 550102
rect 97398 550046 97494 550102
rect 96874 549978 97494 550046
rect 96874 549922 96970 549978
rect 97026 549922 97094 549978
rect 97150 549922 97218 549978
rect 97274 549922 97342 549978
rect 97398 549922 97494 549978
rect 96874 532350 97494 549922
rect 96874 532294 96970 532350
rect 97026 532294 97094 532350
rect 97150 532294 97218 532350
rect 97274 532294 97342 532350
rect 97398 532294 97494 532350
rect 96874 532226 97494 532294
rect 96874 532170 96970 532226
rect 97026 532170 97094 532226
rect 97150 532170 97218 532226
rect 97274 532170 97342 532226
rect 97398 532170 97494 532226
rect 96874 532102 97494 532170
rect 96874 532046 96970 532102
rect 97026 532046 97094 532102
rect 97150 532046 97218 532102
rect 97274 532046 97342 532102
rect 97398 532046 97494 532102
rect 96874 531978 97494 532046
rect 96874 531922 96970 531978
rect 97026 531922 97094 531978
rect 97150 531922 97218 531978
rect 97274 531922 97342 531978
rect 97398 531922 97494 531978
rect 96874 514350 97494 531922
rect 96874 514294 96970 514350
rect 97026 514294 97094 514350
rect 97150 514294 97218 514350
rect 97274 514294 97342 514350
rect 97398 514294 97494 514350
rect 96874 514226 97494 514294
rect 96874 514170 96970 514226
rect 97026 514170 97094 514226
rect 97150 514170 97218 514226
rect 97274 514170 97342 514226
rect 97398 514170 97494 514226
rect 96874 514102 97494 514170
rect 96874 514046 96970 514102
rect 97026 514046 97094 514102
rect 97150 514046 97218 514102
rect 97274 514046 97342 514102
rect 97398 514046 97494 514102
rect 96874 513978 97494 514046
rect 96874 513922 96970 513978
rect 97026 513922 97094 513978
rect 97150 513922 97218 513978
rect 97274 513922 97342 513978
rect 97398 513922 97494 513978
rect 96874 496350 97494 513922
rect 96874 496294 96970 496350
rect 97026 496294 97094 496350
rect 97150 496294 97218 496350
rect 97274 496294 97342 496350
rect 97398 496294 97494 496350
rect 96874 496226 97494 496294
rect 96874 496170 96970 496226
rect 97026 496170 97094 496226
rect 97150 496170 97218 496226
rect 97274 496170 97342 496226
rect 97398 496170 97494 496226
rect 96874 496102 97494 496170
rect 96874 496046 96970 496102
rect 97026 496046 97094 496102
rect 97150 496046 97218 496102
rect 97274 496046 97342 496102
rect 97398 496046 97494 496102
rect 96874 495978 97494 496046
rect 96874 495922 96970 495978
rect 97026 495922 97094 495978
rect 97150 495922 97218 495978
rect 97274 495922 97342 495978
rect 97398 495922 97494 495978
rect 96874 478350 97494 495922
rect 96874 478294 96970 478350
rect 97026 478294 97094 478350
rect 97150 478294 97218 478350
rect 97274 478294 97342 478350
rect 97398 478294 97494 478350
rect 96874 478226 97494 478294
rect 96874 478170 96970 478226
rect 97026 478170 97094 478226
rect 97150 478170 97218 478226
rect 97274 478170 97342 478226
rect 97398 478170 97494 478226
rect 96874 478102 97494 478170
rect 96874 478046 96970 478102
rect 97026 478046 97094 478102
rect 97150 478046 97218 478102
rect 97274 478046 97342 478102
rect 97398 478046 97494 478102
rect 96874 477978 97494 478046
rect 96874 477922 96970 477978
rect 97026 477922 97094 477978
rect 97150 477922 97218 477978
rect 97274 477922 97342 477978
rect 97398 477922 97494 477978
rect 96874 460350 97494 477922
rect 96874 460294 96970 460350
rect 97026 460294 97094 460350
rect 97150 460294 97218 460350
rect 97274 460294 97342 460350
rect 97398 460294 97494 460350
rect 96874 460226 97494 460294
rect 96874 460170 96970 460226
rect 97026 460170 97094 460226
rect 97150 460170 97218 460226
rect 97274 460170 97342 460226
rect 97398 460170 97494 460226
rect 96874 460102 97494 460170
rect 96874 460046 96970 460102
rect 97026 460046 97094 460102
rect 97150 460046 97218 460102
rect 97274 460046 97342 460102
rect 97398 460046 97494 460102
rect 96874 459978 97494 460046
rect 96874 459922 96970 459978
rect 97026 459922 97094 459978
rect 97150 459922 97218 459978
rect 97274 459922 97342 459978
rect 97398 459922 97494 459978
rect 96874 442350 97494 459922
rect 96874 442294 96970 442350
rect 97026 442294 97094 442350
rect 97150 442294 97218 442350
rect 97274 442294 97342 442350
rect 97398 442294 97494 442350
rect 96874 442226 97494 442294
rect 96874 442170 96970 442226
rect 97026 442170 97094 442226
rect 97150 442170 97218 442226
rect 97274 442170 97342 442226
rect 97398 442170 97494 442226
rect 96874 442102 97494 442170
rect 96874 442046 96970 442102
rect 97026 442046 97094 442102
rect 97150 442046 97218 442102
rect 97274 442046 97342 442102
rect 97398 442046 97494 442102
rect 96874 441978 97494 442046
rect 96874 441922 96970 441978
rect 97026 441922 97094 441978
rect 97150 441922 97218 441978
rect 97274 441922 97342 441978
rect 97398 441922 97494 441978
rect 96874 424350 97494 441922
rect 96874 424294 96970 424350
rect 97026 424294 97094 424350
rect 97150 424294 97218 424350
rect 97274 424294 97342 424350
rect 97398 424294 97494 424350
rect 96874 424226 97494 424294
rect 96874 424170 96970 424226
rect 97026 424170 97094 424226
rect 97150 424170 97218 424226
rect 97274 424170 97342 424226
rect 97398 424170 97494 424226
rect 96874 424102 97494 424170
rect 96874 424046 96970 424102
rect 97026 424046 97094 424102
rect 97150 424046 97218 424102
rect 97274 424046 97342 424102
rect 97398 424046 97494 424102
rect 96874 423978 97494 424046
rect 96874 423922 96970 423978
rect 97026 423922 97094 423978
rect 97150 423922 97218 423978
rect 97274 423922 97342 423978
rect 97398 423922 97494 423978
rect 96874 406350 97494 423922
rect 96874 406294 96970 406350
rect 97026 406294 97094 406350
rect 97150 406294 97218 406350
rect 97274 406294 97342 406350
rect 97398 406294 97494 406350
rect 96874 406226 97494 406294
rect 96874 406170 96970 406226
rect 97026 406170 97094 406226
rect 97150 406170 97218 406226
rect 97274 406170 97342 406226
rect 97398 406170 97494 406226
rect 96874 406102 97494 406170
rect 96874 406046 96970 406102
rect 97026 406046 97094 406102
rect 97150 406046 97218 406102
rect 97274 406046 97342 406102
rect 97398 406046 97494 406102
rect 96874 405978 97494 406046
rect 96874 405922 96970 405978
rect 97026 405922 97094 405978
rect 97150 405922 97218 405978
rect 97274 405922 97342 405978
rect 97398 405922 97494 405978
rect 96874 388350 97494 405922
rect 96874 388294 96970 388350
rect 97026 388294 97094 388350
rect 97150 388294 97218 388350
rect 97274 388294 97342 388350
rect 97398 388294 97494 388350
rect 96874 388226 97494 388294
rect 96874 388170 96970 388226
rect 97026 388170 97094 388226
rect 97150 388170 97218 388226
rect 97274 388170 97342 388226
rect 97398 388170 97494 388226
rect 96874 388102 97494 388170
rect 96874 388046 96970 388102
rect 97026 388046 97094 388102
rect 97150 388046 97218 388102
rect 97274 388046 97342 388102
rect 97398 388046 97494 388102
rect 96874 387978 97494 388046
rect 96874 387922 96970 387978
rect 97026 387922 97094 387978
rect 97150 387922 97218 387978
rect 97274 387922 97342 387978
rect 97398 387922 97494 387978
rect 96874 370350 97494 387922
rect 96874 370294 96970 370350
rect 97026 370294 97094 370350
rect 97150 370294 97218 370350
rect 97274 370294 97342 370350
rect 97398 370294 97494 370350
rect 96874 370226 97494 370294
rect 96874 370170 96970 370226
rect 97026 370170 97094 370226
rect 97150 370170 97218 370226
rect 97274 370170 97342 370226
rect 97398 370170 97494 370226
rect 96874 370102 97494 370170
rect 96874 370046 96970 370102
rect 97026 370046 97094 370102
rect 97150 370046 97218 370102
rect 97274 370046 97342 370102
rect 97398 370046 97494 370102
rect 96874 369978 97494 370046
rect 96874 369922 96970 369978
rect 97026 369922 97094 369978
rect 97150 369922 97218 369978
rect 97274 369922 97342 369978
rect 97398 369922 97494 369978
rect 96874 352350 97494 369922
rect 96874 352294 96970 352350
rect 97026 352294 97094 352350
rect 97150 352294 97218 352350
rect 97274 352294 97342 352350
rect 97398 352294 97494 352350
rect 96874 352226 97494 352294
rect 96874 352170 96970 352226
rect 97026 352170 97094 352226
rect 97150 352170 97218 352226
rect 97274 352170 97342 352226
rect 97398 352170 97494 352226
rect 96874 352102 97494 352170
rect 96874 352046 96970 352102
rect 97026 352046 97094 352102
rect 97150 352046 97218 352102
rect 97274 352046 97342 352102
rect 97398 352046 97494 352102
rect 96874 351978 97494 352046
rect 96874 351922 96970 351978
rect 97026 351922 97094 351978
rect 97150 351922 97218 351978
rect 97274 351922 97342 351978
rect 97398 351922 97494 351978
rect 96874 334350 97494 351922
rect 96874 334294 96970 334350
rect 97026 334294 97094 334350
rect 97150 334294 97218 334350
rect 97274 334294 97342 334350
rect 97398 334294 97494 334350
rect 96874 334226 97494 334294
rect 96874 334170 96970 334226
rect 97026 334170 97094 334226
rect 97150 334170 97218 334226
rect 97274 334170 97342 334226
rect 97398 334170 97494 334226
rect 96874 334102 97494 334170
rect 96874 334046 96970 334102
rect 97026 334046 97094 334102
rect 97150 334046 97218 334102
rect 97274 334046 97342 334102
rect 97398 334046 97494 334102
rect 96874 333978 97494 334046
rect 96874 333922 96970 333978
rect 97026 333922 97094 333978
rect 97150 333922 97218 333978
rect 97274 333922 97342 333978
rect 97398 333922 97494 333978
rect 96874 316350 97494 333922
rect 96874 316294 96970 316350
rect 97026 316294 97094 316350
rect 97150 316294 97218 316350
rect 97274 316294 97342 316350
rect 97398 316294 97494 316350
rect 96874 316226 97494 316294
rect 96874 316170 96970 316226
rect 97026 316170 97094 316226
rect 97150 316170 97218 316226
rect 97274 316170 97342 316226
rect 97398 316170 97494 316226
rect 96874 316102 97494 316170
rect 96874 316046 96970 316102
rect 97026 316046 97094 316102
rect 97150 316046 97218 316102
rect 97274 316046 97342 316102
rect 97398 316046 97494 316102
rect 96874 315978 97494 316046
rect 96874 315922 96970 315978
rect 97026 315922 97094 315978
rect 97150 315922 97218 315978
rect 97274 315922 97342 315978
rect 97398 315922 97494 315978
rect 96874 298350 97494 315922
rect 96874 298294 96970 298350
rect 97026 298294 97094 298350
rect 97150 298294 97218 298350
rect 97274 298294 97342 298350
rect 97398 298294 97494 298350
rect 96874 298226 97494 298294
rect 96874 298170 96970 298226
rect 97026 298170 97094 298226
rect 97150 298170 97218 298226
rect 97274 298170 97342 298226
rect 97398 298170 97494 298226
rect 96874 298102 97494 298170
rect 96874 298046 96970 298102
rect 97026 298046 97094 298102
rect 97150 298046 97218 298102
rect 97274 298046 97342 298102
rect 97398 298046 97494 298102
rect 96874 297978 97494 298046
rect 96874 297922 96970 297978
rect 97026 297922 97094 297978
rect 97150 297922 97218 297978
rect 97274 297922 97342 297978
rect 97398 297922 97494 297978
rect 96874 280350 97494 297922
rect 96874 280294 96970 280350
rect 97026 280294 97094 280350
rect 97150 280294 97218 280350
rect 97274 280294 97342 280350
rect 97398 280294 97494 280350
rect 96874 280226 97494 280294
rect 96874 280170 96970 280226
rect 97026 280170 97094 280226
rect 97150 280170 97218 280226
rect 97274 280170 97342 280226
rect 97398 280170 97494 280226
rect 96874 280102 97494 280170
rect 96874 280046 96970 280102
rect 97026 280046 97094 280102
rect 97150 280046 97218 280102
rect 97274 280046 97342 280102
rect 97398 280046 97494 280102
rect 96874 279978 97494 280046
rect 96874 279922 96970 279978
rect 97026 279922 97094 279978
rect 97150 279922 97218 279978
rect 97274 279922 97342 279978
rect 97398 279922 97494 279978
rect 96874 262350 97494 279922
rect 96874 262294 96970 262350
rect 97026 262294 97094 262350
rect 97150 262294 97218 262350
rect 97274 262294 97342 262350
rect 97398 262294 97494 262350
rect 96874 262226 97494 262294
rect 96874 262170 96970 262226
rect 97026 262170 97094 262226
rect 97150 262170 97218 262226
rect 97274 262170 97342 262226
rect 97398 262170 97494 262226
rect 96874 262102 97494 262170
rect 96874 262046 96970 262102
rect 97026 262046 97094 262102
rect 97150 262046 97218 262102
rect 97274 262046 97342 262102
rect 97398 262046 97494 262102
rect 96874 261978 97494 262046
rect 96874 261922 96970 261978
rect 97026 261922 97094 261978
rect 97150 261922 97218 261978
rect 97274 261922 97342 261978
rect 97398 261922 97494 261978
rect 96874 244350 97494 261922
rect 96874 244294 96970 244350
rect 97026 244294 97094 244350
rect 97150 244294 97218 244350
rect 97274 244294 97342 244350
rect 97398 244294 97494 244350
rect 96874 244226 97494 244294
rect 96874 244170 96970 244226
rect 97026 244170 97094 244226
rect 97150 244170 97218 244226
rect 97274 244170 97342 244226
rect 97398 244170 97494 244226
rect 96874 244102 97494 244170
rect 96874 244046 96970 244102
rect 97026 244046 97094 244102
rect 97150 244046 97218 244102
rect 97274 244046 97342 244102
rect 97398 244046 97494 244102
rect 96874 243978 97494 244046
rect 96874 243922 96970 243978
rect 97026 243922 97094 243978
rect 97150 243922 97218 243978
rect 97274 243922 97342 243978
rect 97398 243922 97494 243978
rect 96874 226350 97494 243922
rect 111154 597212 111774 598268
rect 111154 597156 111250 597212
rect 111306 597156 111374 597212
rect 111430 597156 111498 597212
rect 111554 597156 111622 597212
rect 111678 597156 111774 597212
rect 111154 597088 111774 597156
rect 111154 597032 111250 597088
rect 111306 597032 111374 597088
rect 111430 597032 111498 597088
rect 111554 597032 111622 597088
rect 111678 597032 111774 597088
rect 111154 596964 111774 597032
rect 111154 596908 111250 596964
rect 111306 596908 111374 596964
rect 111430 596908 111498 596964
rect 111554 596908 111622 596964
rect 111678 596908 111774 596964
rect 111154 596840 111774 596908
rect 111154 596784 111250 596840
rect 111306 596784 111374 596840
rect 111430 596784 111498 596840
rect 111554 596784 111622 596840
rect 111678 596784 111774 596840
rect 111154 580350 111774 596784
rect 111154 580294 111250 580350
rect 111306 580294 111374 580350
rect 111430 580294 111498 580350
rect 111554 580294 111622 580350
rect 111678 580294 111774 580350
rect 111154 580226 111774 580294
rect 111154 580170 111250 580226
rect 111306 580170 111374 580226
rect 111430 580170 111498 580226
rect 111554 580170 111622 580226
rect 111678 580170 111774 580226
rect 111154 580102 111774 580170
rect 111154 580046 111250 580102
rect 111306 580046 111374 580102
rect 111430 580046 111498 580102
rect 111554 580046 111622 580102
rect 111678 580046 111774 580102
rect 111154 579978 111774 580046
rect 111154 579922 111250 579978
rect 111306 579922 111374 579978
rect 111430 579922 111498 579978
rect 111554 579922 111622 579978
rect 111678 579922 111774 579978
rect 111154 562350 111774 579922
rect 111154 562294 111250 562350
rect 111306 562294 111374 562350
rect 111430 562294 111498 562350
rect 111554 562294 111622 562350
rect 111678 562294 111774 562350
rect 111154 562226 111774 562294
rect 111154 562170 111250 562226
rect 111306 562170 111374 562226
rect 111430 562170 111498 562226
rect 111554 562170 111622 562226
rect 111678 562170 111774 562226
rect 111154 562102 111774 562170
rect 111154 562046 111250 562102
rect 111306 562046 111374 562102
rect 111430 562046 111498 562102
rect 111554 562046 111622 562102
rect 111678 562046 111774 562102
rect 111154 561978 111774 562046
rect 111154 561922 111250 561978
rect 111306 561922 111374 561978
rect 111430 561922 111498 561978
rect 111554 561922 111622 561978
rect 111678 561922 111774 561978
rect 111154 544350 111774 561922
rect 111154 544294 111250 544350
rect 111306 544294 111374 544350
rect 111430 544294 111498 544350
rect 111554 544294 111622 544350
rect 111678 544294 111774 544350
rect 111154 544226 111774 544294
rect 111154 544170 111250 544226
rect 111306 544170 111374 544226
rect 111430 544170 111498 544226
rect 111554 544170 111622 544226
rect 111678 544170 111774 544226
rect 111154 544102 111774 544170
rect 111154 544046 111250 544102
rect 111306 544046 111374 544102
rect 111430 544046 111498 544102
rect 111554 544046 111622 544102
rect 111678 544046 111774 544102
rect 111154 543978 111774 544046
rect 111154 543922 111250 543978
rect 111306 543922 111374 543978
rect 111430 543922 111498 543978
rect 111554 543922 111622 543978
rect 111678 543922 111774 543978
rect 111154 526350 111774 543922
rect 111154 526294 111250 526350
rect 111306 526294 111374 526350
rect 111430 526294 111498 526350
rect 111554 526294 111622 526350
rect 111678 526294 111774 526350
rect 111154 526226 111774 526294
rect 111154 526170 111250 526226
rect 111306 526170 111374 526226
rect 111430 526170 111498 526226
rect 111554 526170 111622 526226
rect 111678 526170 111774 526226
rect 111154 526102 111774 526170
rect 111154 526046 111250 526102
rect 111306 526046 111374 526102
rect 111430 526046 111498 526102
rect 111554 526046 111622 526102
rect 111678 526046 111774 526102
rect 111154 525978 111774 526046
rect 111154 525922 111250 525978
rect 111306 525922 111374 525978
rect 111430 525922 111498 525978
rect 111554 525922 111622 525978
rect 111678 525922 111774 525978
rect 111154 508350 111774 525922
rect 111154 508294 111250 508350
rect 111306 508294 111374 508350
rect 111430 508294 111498 508350
rect 111554 508294 111622 508350
rect 111678 508294 111774 508350
rect 111154 508226 111774 508294
rect 111154 508170 111250 508226
rect 111306 508170 111374 508226
rect 111430 508170 111498 508226
rect 111554 508170 111622 508226
rect 111678 508170 111774 508226
rect 111154 508102 111774 508170
rect 111154 508046 111250 508102
rect 111306 508046 111374 508102
rect 111430 508046 111498 508102
rect 111554 508046 111622 508102
rect 111678 508046 111774 508102
rect 111154 507978 111774 508046
rect 111154 507922 111250 507978
rect 111306 507922 111374 507978
rect 111430 507922 111498 507978
rect 111554 507922 111622 507978
rect 111678 507922 111774 507978
rect 111154 490350 111774 507922
rect 111154 490294 111250 490350
rect 111306 490294 111374 490350
rect 111430 490294 111498 490350
rect 111554 490294 111622 490350
rect 111678 490294 111774 490350
rect 111154 490226 111774 490294
rect 111154 490170 111250 490226
rect 111306 490170 111374 490226
rect 111430 490170 111498 490226
rect 111554 490170 111622 490226
rect 111678 490170 111774 490226
rect 111154 490102 111774 490170
rect 111154 490046 111250 490102
rect 111306 490046 111374 490102
rect 111430 490046 111498 490102
rect 111554 490046 111622 490102
rect 111678 490046 111774 490102
rect 111154 489978 111774 490046
rect 111154 489922 111250 489978
rect 111306 489922 111374 489978
rect 111430 489922 111498 489978
rect 111554 489922 111622 489978
rect 111678 489922 111774 489978
rect 111154 472350 111774 489922
rect 111154 472294 111250 472350
rect 111306 472294 111374 472350
rect 111430 472294 111498 472350
rect 111554 472294 111622 472350
rect 111678 472294 111774 472350
rect 111154 472226 111774 472294
rect 111154 472170 111250 472226
rect 111306 472170 111374 472226
rect 111430 472170 111498 472226
rect 111554 472170 111622 472226
rect 111678 472170 111774 472226
rect 111154 472102 111774 472170
rect 111154 472046 111250 472102
rect 111306 472046 111374 472102
rect 111430 472046 111498 472102
rect 111554 472046 111622 472102
rect 111678 472046 111774 472102
rect 111154 471978 111774 472046
rect 111154 471922 111250 471978
rect 111306 471922 111374 471978
rect 111430 471922 111498 471978
rect 111554 471922 111622 471978
rect 111678 471922 111774 471978
rect 111154 454350 111774 471922
rect 111154 454294 111250 454350
rect 111306 454294 111374 454350
rect 111430 454294 111498 454350
rect 111554 454294 111622 454350
rect 111678 454294 111774 454350
rect 111154 454226 111774 454294
rect 111154 454170 111250 454226
rect 111306 454170 111374 454226
rect 111430 454170 111498 454226
rect 111554 454170 111622 454226
rect 111678 454170 111774 454226
rect 111154 454102 111774 454170
rect 111154 454046 111250 454102
rect 111306 454046 111374 454102
rect 111430 454046 111498 454102
rect 111554 454046 111622 454102
rect 111678 454046 111774 454102
rect 111154 453978 111774 454046
rect 111154 453922 111250 453978
rect 111306 453922 111374 453978
rect 111430 453922 111498 453978
rect 111554 453922 111622 453978
rect 111678 453922 111774 453978
rect 111154 436350 111774 453922
rect 111154 436294 111250 436350
rect 111306 436294 111374 436350
rect 111430 436294 111498 436350
rect 111554 436294 111622 436350
rect 111678 436294 111774 436350
rect 111154 436226 111774 436294
rect 111154 436170 111250 436226
rect 111306 436170 111374 436226
rect 111430 436170 111498 436226
rect 111554 436170 111622 436226
rect 111678 436170 111774 436226
rect 111154 436102 111774 436170
rect 111154 436046 111250 436102
rect 111306 436046 111374 436102
rect 111430 436046 111498 436102
rect 111554 436046 111622 436102
rect 111678 436046 111774 436102
rect 111154 435978 111774 436046
rect 111154 435922 111250 435978
rect 111306 435922 111374 435978
rect 111430 435922 111498 435978
rect 111554 435922 111622 435978
rect 111678 435922 111774 435978
rect 111154 418350 111774 435922
rect 111154 418294 111250 418350
rect 111306 418294 111374 418350
rect 111430 418294 111498 418350
rect 111554 418294 111622 418350
rect 111678 418294 111774 418350
rect 111154 418226 111774 418294
rect 111154 418170 111250 418226
rect 111306 418170 111374 418226
rect 111430 418170 111498 418226
rect 111554 418170 111622 418226
rect 111678 418170 111774 418226
rect 111154 418102 111774 418170
rect 111154 418046 111250 418102
rect 111306 418046 111374 418102
rect 111430 418046 111498 418102
rect 111554 418046 111622 418102
rect 111678 418046 111774 418102
rect 111154 417978 111774 418046
rect 111154 417922 111250 417978
rect 111306 417922 111374 417978
rect 111430 417922 111498 417978
rect 111554 417922 111622 417978
rect 111678 417922 111774 417978
rect 111154 400350 111774 417922
rect 111154 400294 111250 400350
rect 111306 400294 111374 400350
rect 111430 400294 111498 400350
rect 111554 400294 111622 400350
rect 111678 400294 111774 400350
rect 111154 400226 111774 400294
rect 111154 400170 111250 400226
rect 111306 400170 111374 400226
rect 111430 400170 111498 400226
rect 111554 400170 111622 400226
rect 111678 400170 111774 400226
rect 111154 400102 111774 400170
rect 111154 400046 111250 400102
rect 111306 400046 111374 400102
rect 111430 400046 111498 400102
rect 111554 400046 111622 400102
rect 111678 400046 111774 400102
rect 111154 399978 111774 400046
rect 111154 399922 111250 399978
rect 111306 399922 111374 399978
rect 111430 399922 111498 399978
rect 111554 399922 111622 399978
rect 111678 399922 111774 399978
rect 111154 382350 111774 399922
rect 111154 382294 111250 382350
rect 111306 382294 111374 382350
rect 111430 382294 111498 382350
rect 111554 382294 111622 382350
rect 111678 382294 111774 382350
rect 111154 382226 111774 382294
rect 111154 382170 111250 382226
rect 111306 382170 111374 382226
rect 111430 382170 111498 382226
rect 111554 382170 111622 382226
rect 111678 382170 111774 382226
rect 111154 382102 111774 382170
rect 111154 382046 111250 382102
rect 111306 382046 111374 382102
rect 111430 382046 111498 382102
rect 111554 382046 111622 382102
rect 111678 382046 111774 382102
rect 111154 381978 111774 382046
rect 111154 381922 111250 381978
rect 111306 381922 111374 381978
rect 111430 381922 111498 381978
rect 111554 381922 111622 381978
rect 111678 381922 111774 381978
rect 111154 364350 111774 381922
rect 111154 364294 111250 364350
rect 111306 364294 111374 364350
rect 111430 364294 111498 364350
rect 111554 364294 111622 364350
rect 111678 364294 111774 364350
rect 111154 364226 111774 364294
rect 111154 364170 111250 364226
rect 111306 364170 111374 364226
rect 111430 364170 111498 364226
rect 111554 364170 111622 364226
rect 111678 364170 111774 364226
rect 111154 364102 111774 364170
rect 111154 364046 111250 364102
rect 111306 364046 111374 364102
rect 111430 364046 111498 364102
rect 111554 364046 111622 364102
rect 111678 364046 111774 364102
rect 111154 363978 111774 364046
rect 111154 363922 111250 363978
rect 111306 363922 111374 363978
rect 111430 363922 111498 363978
rect 111554 363922 111622 363978
rect 111678 363922 111774 363978
rect 111154 346350 111774 363922
rect 111154 346294 111250 346350
rect 111306 346294 111374 346350
rect 111430 346294 111498 346350
rect 111554 346294 111622 346350
rect 111678 346294 111774 346350
rect 111154 346226 111774 346294
rect 111154 346170 111250 346226
rect 111306 346170 111374 346226
rect 111430 346170 111498 346226
rect 111554 346170 111622 346226
rect 111678 346170 111774 346226
rect 111154 346102 111774 346170
rect 111154 346046 111250 346102
rect 111306 346046 111374 346102
rect 111430 346046 111498 346102
rect 111554 346046 111622 346102
rect 111678 346046 111774 346102
rect 111154 345978 111774 346046
rect 111154 345922 111250 345978
rect 111306 345922 111374 345978
rect 111430 345922 111498 345978
rect 111554 345922 111622 345978
rect 111678 345922 111774 345978
rect 111154 328350 111774 345922
rect 111154 328294 111250 328350
rect 111306 328294 111374 328350
rect 111430 328294 111498 328350
rect 111554 328294 111622 328350
rect 111678 328294 111774 328350
rect 111154 328226 111774 328294
rect 111154 328170 111250 328226
rect 111306 328170 111374 328226
rect 111430 328170 111498 328226
rect 111554 328170 111622 328226
rect 111678 328170 111774 328226
rect 111154 328102 111774 328170
rect 111154 328046 111250 328102
rect 111306 328046 111374 328102
rect 111430 328046 111498 328102
rect 111554 328046 111622 328102
rect 111678 328046 111774 328102
rect 111154 327978 111774 328046
rect 111154 327922 111250 327978
rect 111306 327922 111374 327978
rect 111430 327922 111498 327978
rect 111554 327922 111622 327978
rect 111678 327922 111774 327978
rect 111154 310350 111774 327922
rect 111154 310294 111250 310350
rect 111306 310294 111374 310350
rect 111430 310294 111498 310350
rect 111554 310294 111622 310350
rect 111678 310294 111774 310350
rect 111154 310226 111774 310294
rect 111154 310170 111250 310226
rect 111306 310170 111374 310226
rect 111430 310170 111498 310226
rect 111554 310170 111622 310226
rect 111678 310170 111774 310226
rect 111154 310102 111774 310170
rect 111154 310046 111250 310102
rect 111306 310046 111374 310102
rect 111430 310046 111498 310102
rect 111554 310046 111622 310102
rect 111678 310046 111774 310102
rect 111154 309978 111774 310046
rect 111154 309922 111250 309978
rect 111306 309922 111374 309978
rect 111430 309922 111498 309978
rect 111554 309922 111622 309978
rect 111678 309922 111774 309978
rect 111154 292350 111774 309922
rect 111154 292294 111250 292350
rect 111306 292294 111374 292350
rect 111430 292294 111498 292350
rect 111554 292294 111622 292350
rect 111678 292294 111774 292350
rect 111154 292226 111774 292294
rect 111154 292170 111250 292226
rect 111306 292170 111374 292226
rect 111430 292170 111498 292226
rect 111554 292170 111622 292226
rect 111678 292170 111774 292226
rect 111154 292102 111774 292170
rect 111154 292046 111250 292102
rect 111306 292046 111374 292102
rect 111430 292046 111498 292102
rect 111554 292046 111622 292102
rect 111678 292046 111774 292102
rect 111154 291978 111774 292046
rect 111154 291922 111250 291978
rect 111306 291922 111374 291978
rect 111430 291922 111498 291978
rect 111554 291922 111622 291978
rect 111678 291922 111774 291978
rect 111154 274350 111774 291922
rect 111154 274294 111250 274350
rect 111306 274294 111374 274350
rect 111430 274294 111498 274350
rect 111554 274294 111622 274350
rect 111678 274294 111774 274350
rect 111154 274226 111774 274294
rect 111154 274170 111250 274226
rect 111306 274170 111374 274226
rect 111430 274170 111498 274226
rect 111554 274170 111622 274226
rect 111678 274170 111774 274226
rect 111154 274102 111774 274170
rect 111154 274046 111250 274102
rect 111306 274046 111374 274102
rect 111430 274046 111498 274102
rect 111554 274046 111622 274102
rect 111678 274046 111774 274102
rect 111154 273978 111774 274046
rect 111154 273922 111250 273978
rect 111306 273922 111374 273978
rect 111430 273922 111498 273978
rect 111554 273922 111622 273978
rect 111678 273922 111774 273978
rect 111154 256350 111774 273922
rect 111154 256294 111250 256350
rect 111306 256294 111374 256350
rect 111430 256294 111498 256350
rect 111554 256294 111622 256350
rect 111678 256294 111774 256350
rect 111154 256226 111774 256294
rect 111154 256170 111250 256226
rect 111306 256170 111374 256226
rect 111430 256170 111498 256226
rect 111554 256170 111622 256226
rect 111678 256170 111774 256226
rect 111154 256102 111774 256170
rect 111154 256046 111250 256102
rect 111306 256046 111374 256102
rect 111430 256046 111498 256102
rect 111554 256046 111622 256102
rect 111678 256046 111774 256102
rect 111154 255978 111774 256046
rect 111154 255922 111250 255978
rect 111306 255922 111374 255978
rect 111430 255922 111498 255978
rect 111554 255922 111622 255978
rect 111678 255922 111774 255978
rect 111154 238350 111774 255922
rect 129154 597212 129774 598268
rect 129154 597156 129250 597212
rect 129306 597156 129374 597212
rect 129430 597156 129498 597212
rect 129554 597156 129622 597212
rect 129678 597156 129774 597212
rect 129154 597088 129774 597156
rect 129154 597032 129250 597088
rect 129306 597032 129374 597088
rect 129430 597032 129498 597088
rect 129554 597032 129622 597088
rect 129678 597032 129774 597088
rect 129154 596964 129774 597032
rect 129154 596908 129250 596964
rect 129306 596908 129374 596964
rect 129430 596908 129498 596964
rect 129554 596908 129622 596964
rect 129678 596908 129774 596964
rect 129154 596840 129774 596908
rect 129154 596784 129250 596840
rect 129306 596784 129374 596840
rect 129430 596784 129498 596840
rect 129554 596784 129622 596840
rect 129678 596784 129774 596840
rect 129154 580350 129774 596784
rect 129154 580294 129250 580350
rect 129306 580294 129374 580350
rect 129430 580294 129498 580350
rect 129554 580294 129622 580350
rect 129678 580294 129774 580350
rect 129154 580226 129774 580294
rect 129154 580170 129250 580226
rect 129306 580170 129374 580226
rect 129430 580170 129498 580226
rect 129554 580170 129622 580226
rect 129678 580170 129774 580226
rect 129154 580102 129774 580170
rect 129154 580046 129250 580102
rect 129306 580046 129374 580102
rect 129430 580046 129498 580102
rect 129554 580046 129622 580102
rect 129678 580046 129774 580102
rect 129154 579978 129774 580046
rect 129154 579922 129250 579978
rect 129306 579922 129374 579978
rect 129430 579922 129498 579978
rect 129554 579922 129622 579978
rect 129678 579922 129774 579978
rect 129154 562350 129774 579922
rect 129154 562294 129250 562350
rect 129306 562294 129374 562350
rect 129430 562294 129498 562350
rect 129554 562294 129622 562350
rect 129678 562294 129774 562350
rect 129154 562226 129774 562294
rect 129154 562170 129250 562226
rect 129306 562170 129374 562226
rect 129430 562170 129498 562226
rect 129554 562170 129622 562226
rect 129678 562170 129774 562226
rect 129154 562102 129774 562170
rect 129154 562046 129250 562102
rect 129306 562046 129374 562102
rect 129430 562046 129498 562102
rect 129554 562046 129622 562102
rect 129678 562046 129774 562102
rect 129154 561978 129774 562046
rect 129154 561922 129250 561978
rect 129306 561922 129374 561978
rect 129430 561922 129498 561978
rect 129554 561922 129622 561978
rect 129678 561922 129774 561978
rect 129154 544350 129774 561922
rect 129154 544294 129250 544350
rect 129306 544294 129374 544350
rect 129430 544294 129498 544350
rect 129554 544294 129622 544350
rect 129678 544294 129774 544350
rect 129154 544226 129774 544294
rect 129154 544170 129250 544226
rect 129306 544170 129374 544226
rect 129430 544170 129498 544226
rect 129554 544170 129622 544226
rect 129678 544170 129774 544226
rect 129154 544102 129774 544170
rect 129154 544046 129250 544102
rect 129306 544046 129374 544102
rect 129430 544046 129498 544102
rect 129554 544046 129622 544102
rect 129678 544046 129774 544102
rect 129154 543978 129774 544046
rect 129154 543922 129250 543978
rect 129306 543922 129374 543978
rect 129430 543922 129498 543978
rect 129554 543922 129622 543978
rect 129678 543922 129774 543978
rect 129154 526350 129774 543922
rect 129154 526294 129250 526350
rect 129306 526294 129374 526350
rect 129430 526294 129498 526350
rect 129554 526294 129622 526350
rect 129678 526294 129774 526350
rect 129154 526226 129774 526294
rect 129154 526170 129250 526226
rect 129306 526170 129374 526226
rect 129430 526170 129498 526226
rect 129554 526170 129622 526226
rect 129678 526170 129774 526226
rect 129154 526102 129774 526170
rect 129154 526046 129250 526102
rect 129306 526046 129374 526102
rect 129430 526046 129498 526102
rect 129554 526046 129622 526102
rect 129678 526046 129774 526102
rect 129154 525978 129774 526046
rect 129154 525922 129250 525978
rect 129306 525922 129374 525978
rect 129430 525922 129498 525978
rect 129554 525922 129622 525978
rect 129678 525922 129774 525978
rect 129154 508350 129774 525922
rect 129154 508294 129250 508350
rect 129306 508294 129374 508350
rect 129430 508294 129498 508350
rect 129554 508294 129622 508350
rect 129678 508294 129774 508350
rect 129154 508226 129774 508294
rect 129154 508170 129250 508226
rect 129306 508170 129374 508226
rect 129430 508170 129498 508226
rect 129554 508170 129622 508226
rect 129678 508170 129774 508226
rect 129154 508102 129774 508170
rect 129154 508046 129250 508102
rect 129306 508046 129374 508102
rect 129430 508046 129498 508102
rect 129554 508046 129622 508102
rect 129678 508046 129774 508102
rect 129154 507978 129774 508046
rect 129154 507922 129250 507978
rect 129306 507922 129374 507978
rect 129430 507922 129498 507978
rect 129554 507922 129622 507978
rect 129678 507922 129774 507978
rect 129154 490350 129774 507922
rect 129154 490294 129250 490350
rect 129306 490294 129374 490350
rect 129430 490294 129498 490350
rect 129554 490294 129622 490350
rect 129678 490294 129774 490350
rect 129154 490226 129774 490294
rect 129154 490170 129250 490226
rect 129306 490170 129374 490226
rect 129430 490170 129498 490226
rect 129554 490170 129622 490226
rect 129678 490170 129774 490226
rect 129154 490102 129774 490170
rect 129154 490046 129250 490102
rect 129306 490046 129374 490102
rect 129430 490046 129498 490102
rect 129554 490046 129622 490102
rect 129678 490046 129774 490102
rect 129154 489978 129774 490046
rect 129154 489922 129250 489978
rect 129306 489922 129374 489978
rect 129430 489922 129498 489978
rect 129554 489922 129622 489978
rect 129678 489922 129774 489978
rect 129154 472350 129774 489922
rect 129154 472294 129250 472350
rect 129306 472294 129374 472350
rect 129430 472294 129498 472350
rect 129554 472294 129622 472350
rect 129678 472294 129774 472350
rect 129154 472226 129774 472294
rect 129154 472170 129250 472226
rect 129306 472170 129374 472226
rect 129430 472170 129498 472226
rect 129554 472170 129622 472226
rect 129678 472170 129774 472226
rect 129154 472102 129774 472170
rect 129154 472046 129250 472102
rect 129306 472046 129374 472102
rect 129430 472046 129498 472102
rect 129554 472046 129622 472102
rect 129678 472046 129774 472102
rect 129154 471978 129774 472046
rect 129154 471922 129250 471978
rect 129306 471922 129374 471978
rect 129430 471922 129498 471978
rect 129554 471922 129622 471978
rect 129678 471922 129774 471978
rect 129154 454350 129774 471922
rect 129154 454294 129250 454350
rect 129306 454294 129374 454350
rect 129430 454294 129498 454350
rect 129554 454294 129622 454350
rect 129678 454294 129774 454350
rect 129154 454226 129774 454294
rect 129154 454170 129250 454226
rect 129306 454170 129374 454226
rect 129430 454170 129498 454226
rect 129554 454170 129622 454226
rect 129678 454170 129774 454226
rect 129154 454102 129774 454170
rect 129154 454046 129250 454102
rect 129306 454046 129374 454102
rect 129430 454046 129498 454102
rect 129554 454046 129622 454102
rect 129678 454046 129774 454102
rect 129154 453978 129774 454046
rect 129154 453922 129250 453978
rect 129306 453922 129374 453978
rect 129430 453922 129498 453978
rect 129554 453922 129622 453978
rect 129678 453922 129774 453978
rect 129154 436350 129774 453922
rect 129154 436294 129250 436350
rect 129306 436294 129374 436350
rect 129430 436294 129498 436350
rect 129554 436294 129622 436350
rect 129678 436294 129774 436350
rect 129154 436226 129774 436294
rect 129154 436170 129250 436226
rect 129306 436170 129374 436226
rect 129430 436170 129498 436226
rect 129554 436170 129622 436226
rect 129678 436170 129774 436226
rect 129154 436102 129774 436170
rect 129154 436046 129250 436102
rect 129306 436046 129374 436102
rect 129430 436046 129498 436102
rect 129554 436046 129622 436102
rect 129678 436046 129774 436102
rect 129154 435978 129774 436046
rect 129154 435922 129250 435978
rect 129306 435922 129374 435978
rect 129430 435922 129498 435978
rect 129554 435922 129622 435978
rect 129678 435922 129774 435978
rect 129154 418350 129774 435922
rect 129154 418294 129250 418350
rect 129306 418294 129374 418350
rect 129430 418294 129498 418350
rect 129554 418294 129622 418350
rect 129678 418294 129774 418350
rect 129154 418226 129774 418294
rect 129154 418170 129250 418226
rect 129306 418170 129374 418226
rect 129430 418170 129498 418226
rect 129554 418170 129622 418226
rect 129678 418170 129774 418226
rect 129154 418102 129774 418170
rect 129154 418046 129250 418102
rect 129306 418046 129374 418102
rect 129430 418046 129498 418102
rect 129554 418046 129622 418102
rect 129678 418046 129774 418102
rect 129154 417978 129774 418046
rect 129154 417922 129250 417978
rect 129306 417922 129374 417978
rect 129430 417922 129498 417978
rect 129554 417922 129622 417978
rect 129678 417922 129774 417978
rect 129154 400350 129774 417922
rect 129154 400294 129250 400350
rect 129306 400294 129374 400350
rect 129430 400294 129498 400350
rect 129554 400294 129622 400350
rect 129678 400294 129774 400350
rect 129154 400226 129774 400294
rect 129154 400170 129250 400226
rect 129306 400170 129374 400226
rect 129430 400170 129498 400226
rect 129554 400170 129622 400226
rect 129678 400170 129774 400226
rect 129154 400102 129774 400170
rect 129154 400046 129250 400102
rect 129306 400046 129374 400102
rect 129430 400046 129498 400102
rect 129554 400046 129622 400102
rect 129678 400046 129774 400102
rect 129154 399978 129774 400046
rect 129154 399922 129250 399978
rect 129306 399922 129374 399978
rect 129430 399922 129498 399978
rect 129554 399922 129622 399978
rect 129678 399922 129774 399978
rect 129154 382350 129774 399922
rect 129154 382294 129250 382350
rect 129306 382294 129374 382350
rect 129430 382294 129498 382350
rect 129554 382294 129622 382350
rect 129678 382294 129774 382350
rect 129154 382226 129774 382294
rect 129154 382170 129250 382226
rect 129306 382170 129374 382226
rect 129430 382170 129498 382226
rect 129554 382170 129622 382226
rect 129678 382170 129774 382226
rect 129154 382102 129774 382170
rect 129154 382046 129250 382102
rect 129306 382046 129374 382102
rect 129430 382046 129498 382102
rect 129554 382046 129622 382102
rect 129678 382046 129774 382102
rect 129154 381978 129774 382046
rect 129154 381922 129250 381978
rect 129306 381922 129374 381978
rect 129430 381922 129498 381978
rect 129554 381922 129622 381978
rect 129678 381922 129774 381978
rect 129154 364350 129774 381922
rect 129154 364294 129250 364350
rect 129306 364294 129374 364350
rect 129430 364294 129498 364350
rect 129554 364294 129622 364350
rect 129678 364294 129774 364350
rect 129154 364226 129774 364294
rect 129154 364170 129250 364226
rect 129306 364170 129374 364226
rect 129430 364170 129498 364226
rect 129554 364170 129622 364226
rect 129678 364170 129774 364226
rect 129154 364102 129774 364170
rect 129154 364046 129250 364102
rect 129306 364046 129374 364102
rect 129430 364046 129498 364102
rect 129554 364046 129622 364102
rect 129678 364046 129774 364102
rect 129154 363978 129774 364046
rect 129154 363922 129250 363978
rect 129306 363922 129374 363978
rect 129430 363922 129498 363978
rect 129554 363922 129622 363978
rect 129678 363922 129774 363978
rect 129154 346350 129774 363922
rect 129154 346294 129250 346350
rect 129306 346294 129374 346350
rect 129430 346294 129498 346350
rect 129554 346294 129622 346350
rect 129678 346294 129774 346350
rect 129154 346226 129774 346294
rect 129154 346170 129250 346226
rect 129306 346170 129374 346226
rect 129430 346170 129498 346226
rect 129554 346170 129622 346226
rect 129678 346170 129774 346226
rect 129154 346102 129774 346170
rect 129154 346046 129250 346102
rect 129306 346046 129374 346102
rect 129430 346046 129498 346102
rect 129554 346046 129622 346102
rect 129678 346046 129774 346102
rect 129154 345978 129774 346046
rect 129154 345922 129250 345978
rect 129306 345922 129374 345978
rect 129430 345922 129498 345978
rect 129554 345922 129622 345978
rect 129678 345922 129774 345978
rect 129154 328350 129774 345922
rect 129154 328294 129250 328350
rect 129306 328294 129374 328350
rect 129430 328294 129498 328350
rect 129554 328294 129622 328350
rect 129678 328294 129774 328350
rect 129154 328226 129774 328294
rect 129154 328170 129250 328226
rect 129306 328170 129374 328226
rect 129430 328170 129498 328226
rect 129554 328170 129622 328226
rect 129678 328170 129774 328226
rect 129154 328102 129774 328170
rect 129154 328046 129250 328102
rect 129306 328046 129374 328102
rect 129430 328046 129498 328102
rect 129554 328046 129622 328102
rect 129678 328046 129774 328102
rect 129154 327978 129774 328046
rect 129154 327922 129250 327978
rect 129306 327922 129374 327978
rect 129430 327922 129498 327978
rect 129554 327922 129622 327978
rect 129678 327922 129774 327978
rect 129154 310350 129774 327922
rect 129154 310294 129250 310350
rect 129306 310294 129374 310350
rect 129430 310294 129498 310350
rect 129554 310294 129622 310350
rect 129678 310294 129774 310350
rect 129154 310226 129774 310294
rect 129154 310170 129250 310226
rect 129306 310170 129374 310226
rect 129430 310170 129498 310226
rect 129554 310170 129622 310226
rect 129678 310170 129774 310226
rect 129154 310102 129774 310170
rect 129154 310046 129250 310102
rect 129306 310046 129374 310102
rect 129430 310046 129498 310102
rect 129554 310046 129622 310102
rect 129678 310046 129774 310102
rect 129154 309978 129774 310046
rect 129154 309922 129250 309978
rect 129306 309922 129374 309978
rect 129430 309922 129498 309978
rect 129554 309922 129622 309978
rect 129678 309922 129774 309978
rect 129154 292350 129774 309922
rect 129154 292294 129250 292350
rect 129306 292294 129374 292350
rect 129430 292294 129498 292350
rect 129554 292294 129622 292350
rect 129678 292294 129774 292350
rect 129154 292226 129774 292294
rect 129154 292170 129250 292226
rect 129306 292170 129374 292226
rect 129430 292170 129498 292226
rect 129554 292170 129622 292226
rect 129678 292170 129774 292226
rect 129154 292102 129774 292170
rect 129154 292046 129250 292102
rect 129306 292046 129374 292102
rect 129430 292046 129498 292102
rect 129554 292046 129622 292102
rect 129678 292046 129774 292102
rect 129154 291978 129774 292046
rect 129154 291922 129250 291978
rect 129306 291922 129374 291978
rect 129430 291922 129498 291978
rect 129554 291922 129622 291978
rect 129678 291922 129774 291978
rect 129154 274350 129774 291922
rect 129154 274294 129250 274350
rect 129306 274294 129374 274350
rect 129430 274294 129498 274350
rect 129554 274294 129622 274350
rect 129678 274294 129774 274350
rect 129154 274226 129774 274294
rect 129154 274170 129250 274226
rect 129306 274170 129374 274226
rect 129430 274170 129498 274226
rect 129554 274170 129622 274226
rect 129678 274170 129774 274226
rect 129154 274102 129774 274170
rect 129154 274046 129250 274102
rect 129306 274046 129374 274102
rect 129430 274046 129498 274102
rect 129554 274046 129622 274102
rect 129678 274046 129774 274102
rect 129154 273978 129774 274046
rect 129154 273922 129250 273978
rect 129306 273922 129374 273978
rect 129430 273922 129498 273978
rect 129554 273922 129622 273978
rect 129678 273922 129774 273978
rect 129154 256350 129774 273922
rect 129154 256294 129250 256350
rect 129306 256294 129374 256350
rect 129430 256294 129498 256350
rect 129554 256294 129622 256350
rect 129678 256294 129774 256350
rect 129154 256226 129774 256294
rect 129154 256170 129250 256226
rect 129306 256170 129374 256226
rect 129430 256170 129498 256226
rect 129554 256170 129622 256226
rect 129678 256170 129774 256226
rect 129154 256102 129774 256170
rect 129154 256046 129250 256102
rect 129306 256046 129374 256102
rect 129430 256046 129498 256102
rect 129554 256046 129622 256102
rect 129678 256046 129774 256102
rect 129154 255978 129774 256046
rect 129154 255922 129250 255978
rect 129306 255922 129374 255978
rect 129430 255922 129498 255978
rect 129554 255922 129622 255978
rect 129678 255922 129774 255978
rect 111154 238294 111250 238350
rect 111306 238294 111374 238350
rect 111430 238294 111498 238350
rect 111554 238294 111622 238350
rect 111678 238294 111774 238350
rect 111154 238226 111774 238294
rect 111154 238170 111250 238226
rect 111306 238170 111374 238226
rect 111430 238170 111498 238226
rect 111554 238170 111622 238226
rect 111678 238170 111774 238226
rect 111154 238102 111774 238170
rect 111154 238046 111250 238102
rect 111306 238046 111374 238102
rect 111430 238046 111498 238102
rect 111554 238046 111622 238102
rect 111678 238046 111774 238102
rect 111154 237978 111774 238046
rect 111154 237922 111250 237978
rect 111306 237922 111374 237978
rect 111430 237922 111498 237978
rect 111554 237922 111622 237978
rect 111678 237922 111774 237978
rect 96874 226294 96970 226350
rect 97026 226294 97094 226350
rect 97150 226294 97218 226350
rect 97274 226294 97342 226350
rect 97398 226294 97494 226350
rect 96874 226226 97494 226294
rect 96874 226170 96970 226226
rect 97026 226170 97094 226226
rect 97150 226170 97218 226226
rect 97274 226170 97342 226226
rect 97398 226170 97494 226226
rect 96874 226102 97494 226170
rect 96874 226046 96970 226102
rect 97026 226046 97094 226102
rect 97150 226046 97218 226102
rect 97274 226046 97342 226102
rect 97398 226046 97494 226102
rect 96874 225978 97494 226046
rect 96874 225922 96970 225978
rect 97026 225922 97094 225978
rect 97150 225922 97218 225978
rect 97274 225922 97342 225978
rect 97398 225922 97494 225978
rect 93154 220294 93250 220350
rect 93306 220294 93374 220350
rect 93430 220294 93498 220350
rect 93554 220294 93622 220350
rect 93678 220294 93774 220350
rect 93154 220226 93774 220294
rect 93154 220170 93250 220226
rect 93306 220170 93374 220226
rect 93430 220170 93498 220226
rect 93554 220170 93622 220226
rect 93678 220170 93774 220226
rect 93154 220102 93774 220170
rect 93154 220046 93250 220102
rect 93306 220046 93374 220102
rect 93430 220046 93498 220102
rect 93554 220046 93622 220102
rect 93678 220046 93774 220102
rect 93154 219978 93774 220046
rect 93154 219922 93250 219978
rect 93306 219922 93374 219978
rect 93430 219922 93498 219978
rect 93554 219922 93622 219978
rect 93678 219922 93774 219978
rect 93154 219134 93774 219922
rect 95168 220350 95488 220384
rect 95168 220294 95238 220350
rect 95294 220294 95362 220350
rect 95418 220294 95488 220350
rect 95168 220226 95488 220294
rect 95168 220170 95238 220226
rect 95294 220170 95362 220226
rect 95418 220170 95488 220226
rect 95168 220102 95488 220170
rect 95168 220046 95238 220102
rect 95294 220046 95362 220102
rect 95418 220046 95488 220102
rect 95168 219978 95488 220046
rect 95168 219922 95238 219978
rect 95294 219922 95362 219978
rect 95418 219922 95488 219978
rect 95168 219888 95488 219922
rect 96874 219134 97494 225922
rect 110528 226350 110848 226384
rect 110528 226294 110598 226350
rect 110654 226294 110722 226350
rect 110778 226294 110848 226350
rect 110528 226226 110848 226294
rect 110528 226170 110598 226226
rect 110654 226170 110722 226226
rect 110778 226170 110848 226226
rect 110528 226102 110848 226170
rect 110528 226046 110598 226102
rect 110654 226046 110722 226102
rect 110778 226046 110848 226102
rect 110528 225978 110848 226046
rect 110528 225922 110598 225978
rect 110654 225922 110722 225978
rect 110778 225922 110848 225978
rect 110528 225888 110848 225922
rect 111154 220350 111774 237922
rect 111154 220294 111250 220350
rect 111306 220294 111374 220350
rect 111430 220294 111498 220350
rect 111554 220294 111622 220350
rect 111678 220294 111774 220350
rect 111154 220226 111774 220294
rect 111154 220170 111250 220226
rect 111306 220170 111374 220226
rect 111430 220170 111498 220226
rect 111554 220170 111622 220226
rect 111678 220170 111774 220226
rect 111154 220102 111774 220170
rect 111154 220046 111250 220102
rect 111306 220046 111374 220102
rect 111430 220046 111498 220102
rect 111554 220046 111622 220102
rect 111678 220046 111774 220102
rect 111154 219978 111774 220046
rect 111154 219922 111250 219978
rect 111306 219922 111374 219978
rect 111430 219922 111498 219978
rect 111554 219922 111622 219978
rect 111678 219922 111774 219978
rect 111154 219134 111774 219922
rect 114874 226350 115494 242964
rect 114874 226294 114970 226350
rect 115026 226294 115094 226350
rect 115150 226294 115218 226350
rect 115274 226294 115342 226350
rect 115398 226294 115494 226350
rect 114874 226226 115494 226294
rect 114874 226170 114970 226226
rect 115026 226170 115094 226226
rect 115150 226170 115218 226226
rect 115274 226170 115342 226226
rect 115398 226170 115494 226226
rect 114874 226102 115494 226170
rect 114874 226046 114970 226102
rect 115026 226046 115094 226102
rect 115150 226046 115218 226102
rect 115274 226046 115342 226102
rect 115398 226046 115494 226102
rect 114874 225978 115494 226046
rect 114874 225922 114970 225978
rect 115026 225922 115094 225978
rect 115150 225922 115218 225978
rect 115274 225922 115342 225978
rect 115398 225922 115494 225978
rect 114874 219134 115494 225922
rect 129154 238350 129774 255922
rect 129154 238294 129250 238350
rect 129306 238294 129374 238350
rect 129430 238294 129498 238350
rect 129554 238294 129622 238350
rect 129678 238294 129774 238350
rect 129154 238226 129774 238294
rect 129154 238170 129250 238226
rect 129306 238170 129374 238226
rect 129430 238170 129498 238226
rect 129554 238170 129622 238226
rect 129678 238170 129774 238226
rect 129154 238102 129774 238170
rect 129154 238046 129250 238102
rect 129306 238046 129374 238102
rect 129430 238046 129498 238102
rect 129554 238046 129622 238102
rect 129678 238046 129774 238102
rect 129154 237978 129774 238046
rect 129154 237922 129250 237978
rect 129306 237922 129374 237978
rect 129430 237922 129498 237978
rect 129554 237922 129622 237978
rect 129678 237922 129774 237978
rect 125888 220350 126208 220384
rect 125888 220294 125958 220350
rect 126014 220294 126082 220350
rect 126138 220294 126208 220350
rect 125888 220226 126208 220294
rect 125888 220170 125958 220226
rect 126014 220170 126082 220226
rect 126138 220170 126208 220226
rect 125888 220102 126208 220170
rect 125888 220046 125958 220102
rect 126014 220046 126082 220102
rect 126138 220046 126208 220102
rect 125888 219978 126208 220046
rect 125888 219922 125958 219978
rect 126014 219922 126082 219978
rect 126138 219922 126208 219978
rect 125888 219888 126208 219922
rect 129154 220350 129774 237922
rect 129154 220294 129250 220350
rect 129306 220294 129374 220350
rect 129430 220294 129498 220350
rect 129554 220294 129622 220350
rect 129678 220294 129774 220350
rect 129154 220226 129774 220294
rect 129154 220170 129250 220226
rect 129306 220170 129374 220226
rect 129430 220170 129498 220226
rect 129554 220170 129622 220226
rect 129678 220170 129774 220226
rect 129154 220102 129774 220170
rect 129154 220046 129250 220102
rect 129306 220046 129374 220102
rect 129430 220046 129498 220102
rect 129554 220046 129622 220102
rect 129678 220046 129774 220102
rect 129154 219978 129774 220046
rect 129154 219922 129250 219978
rect 129306 219922 129374 219978
rect 129430 219922 129498 219978
rect 129554 219922 129622 219978
rect 129678 219922 129774 219978
rect 129154 219134 129774 219922
rect 132874 598172 133494 598268
rect 132874 598116 132970 598172
rect 133026 598116 133094 598172
rect 133150 598116 133218 598172
rect 133274 598116 133342 598172
rect 133398 598116 133494 598172
rect 132874 598048 133494 598116
rect 132874 597992 132970 598048
rect 133026 597992 133094 598048
rect 133150 597992 133218 598048
rect 133274 597992 133342 598048
rect 133398 597992 133494 598048
rect 132874 597924 133494 597992
rect 132874 597868 132970 597924
rect 133026 597868 133094 597924
rect 133150 597868 133218 597924
rect 133274 597868 133342 597924
rect 133398 597868 133494 597924
rect 132874 597800 133494 597868
rect 132874 597744 132970 597800
rect 133026 597744 133094 597800
rect 133150 597744 133218 597800
rect 133274 597744 133342 597800
rect 133398 597744 133494 597800
rect 132874 586350 133494 597744
rect 132874 586294 132970 586350
rect 133026 586294 133094 586350
rect 133150 586294 133218 586350
rect 133274 586294 133342 586350
rect 133398 586294 133494 586350
rect 132874 586226 133494 586294
rect 132874 586170 132970 586226
rect 133026 586170 133094 586226
rect 133150 586170 133218 586226
rect 133274 586170 133342 586226
rect 133398 586170 133494 586226
rect 132874 586102 133494 586170
rect 132874 586046 132970 586102
rect 133026 586046 133094 586102
rect 133150 586046 133218 586102
rect 133274 586046 133342 586102
rect 133398 586046 133494 586102
rect 132874 585978 133494 586046
rect 132874 585922 132970 585978
rect 133026 585922 133094 585978
rect 133150 585922 133218 585978
rect 133274 585922 133342 585978
rect 133398 585922 133494 585978
rect 132874 568350 133494 585922
rect 132874 568294 132970 568350
rect 133026 568294 133094 568350
rect 133150 568294 133218 568350
rect 133274 568294 133342 568350
rect 133398 568294 133494 568350
rect 132874 568226 133494 568294
rect 132874 568170 132970 568226
rect 133026 568170 133094 568226
rect 133150 568170 133218 568226
rect 133274 568170 133342 568226
rect 133398 568170 133494 568226
rect 132874 568102 133494 568170
rect 132874 568046 132970 568102
rect 133026 568046 133094 568102
rect 133150 568046 133218 568102
rect 133274 568046 133342 568102
rect 133398 568046 133494 568102
rect 132874 567978 133494 568046
rect 132874 567922 132970 567978
rect 133026 567922 133094 567978
rect 133150 567922 133218 567978
rect 133274 567922 133342 567978
rect 133398 567922 133494 567978
rect 132874 550350 133494 567922
rect 132874 550294 132970 550350
rect 133026 550294 133094 550350
rect 133150 550294 133218 550350
rect 133274 550294 133342 550350
rect 133398 550294 133494 550350
rect 132874 550226 133494 550294
rect 132874 550170 132970 550226
rect 133026 550170 133094 550226
rect 133150 550170 133218 550226
rect 133274 550170 133342 550226
rect 133398 550170 133494 550226
rect 132874 550102 133494 550170
rect 132874 550046 132970 550102
rect 133026 550046 133094 550102
rect 133150 550046 133218 550102
rect 133274 550046 133342 550102
rect 133398 550046 133494 550102
rect 132874 549978 133494 550046
rect 132874 549922 132970 549978
rect 133026 549922 133094 549978
rect 133150 549922 133218 549978
rect 133274 549922 133342 549978
rect 133398 549922 133494 549978
rect 132874 532350 133494 549922
rect 132874 532294 132970 532350
rect 133026 532294 133094 532350
rect 133150 532294 133218 532350
rect 133274 532294 133342 532350
rect 133398 532294 133494 532350
rect 132874 532226 133494 532294
rect 132874 532170 132970 532226
rect 133026 532170 133094 532226
rect 133150 532170 133218 532226
rect 133274 532170 133342 532226
rect 133398 532170 133494 532226
rect 132874 532102 133494 532170
rect 132874 532046 132970 532102
rect 133026 532046 133094 532102
rect 133150 532046 133218 532102
rect 133274 532046 133342 532102
rect 133398 532046 133494 532102
rect 132874 531978 133494 532046
rect 132874 531922 132970 531978
rect 133026 531922 133094 531978
rect 133150 531922 133218 531978
rect 133274 531922 133342 531978
rect 133398 531922 133494 531978
rect 132874 514350 133494 531922
rect 132874 514294 132970 514350
rect 133026 514294 133094 514350
rect 133150 514294 133218 514350
rect 133274 514294 133342 514350
rect 133398 514294 133494 514350
rect 132874 514226 133494 514294
rect 132874 514170 132970 514226
rect 133026 514170 133094 514226
rect 133150 514170 133218 514226
rect 133274 514170 133342 514226
rect 133398 514170 133494 514226
rect 132874 514102 133494 514170
rect 132874 514046 132970 514102
rect 133026 514046 133094 514102
rect 133150 514046 133218 514102
rect 133274 514046 133342 514102
rect 133398 514046 133494 514102
rect 132874 513978 133494 514046
rect 132874 513922 132970 513978
rect 133026 513922 133094 513978
rect 133150 513922 133218 513978
rect 133274 513922 133342 513978
rect 133398 513922 133494 513978
rect 132874 496350 133494 513922
rect 132874 496294 132970 496350
rect 133026 496294 133094 496350
rect 133150 496294 133218 496350
rect 133274 496294 133342 496350
rect 133398 496294 133494 496350
rect 132874 496226 133494 496294
rect 132874 496170 132970 496226
rect 133026 496170 133094 496226
rect 133150 496170 133218 496226
rect 133274 496170 133342 496226
rect 133398 496170 133494 496226
rect 132874 496102 133494 496170
rect 132874 496046 132970 496102
rect 133026 496046 133094 496102
rect 133150 496046 133218 496102
rect 133274 496046 133342 496102
rect 133398 496046 133494 496102
rect 132874 495978 133494 496046
rect 132874 495922 132970 495978
rect 133026 495922 133094 495978
rect 133150 495922 133218 495978
rect 133274 495922 133342 495978
rect 133398 495922 133494 495978
rect 132874 478350 133494 495922
rect 132874 478294 132970 478350
rect 133026 478294 133094 478350
rect 133150 478294 133218 478350
rect 133274 478294 133342 478350
rect 133398 478294 133494 478350
rect 132874 478226 133494 478294
rect 132874 478170 132970 478226
rect 133026 478170 133094 478226
rect 133150 478170 133218 478226
rect 133274 478170 133342 478226
rect 133398 478170 133494 478226
rect 132874 478102 133494 478170
rect 132874 478046 132970 478102
rect 133026 478046 133094 478102
rect 133150 478046 133218 478102
rect 133274 478046 133342 478102
rect 133398 478046 133494 478102
rect 132874 477978 133494 478046
rect 132874 477922 132970 477978
rect 133026 477922 133094 477978
rect 133150 477922 133218 477978
rect 133274 477922 133342 477978
rect 133398 477922 133494 477978
rect 132874 460350 133494 477922
rect 132874 460294 132970 460350
rect 133026 460294 133094 460350
rect 133150 460294 133218 460350
rect 133274 460294 133342 460350
rect 133398 460294 133494 460350
rect 132874 460226 133494 460294
rect 132874 460170 132970 460226
rect 133026 460170 133094 460226
rect 133150 460170 133218 460226
rect 133274 460170 133342 460226
rect 133398 460170 133494 460226
rect 132874 460102 133494 460170
rect 132874 460046 132970 460102
rect 133026 460046 133094 460102
rect 133150 460046 133218 460102
rect 133274 460046 133342 460102
rect 133398 460046 133494 460102
rect 132874 459978 133494 460046
rect 132874 459922 132970 459978
rect 133026 459922 133094 459978
rect 133150 459922 133218 459978
rect 133274 459922 133342 459978
rect 133398 459922 133494 459978
rect 132874 442350 133494 459922
rect 132874 442294 132970 442350
rect 133026 442294 133094 442350
rect 133150 442294 133218 442350
rect 133274 442294 133342 442350
rect 133398 442294 133494 442350
rect 132874 442226 133494 442294
rect 132874 442170 132970 442226
rect 133026 442170 133094 442226
rect 133150 442170 133218 442226
rect 133274 442170 133342 442226
rect 133398 442170 133494 442226
rect 132874 442102 133494 442170
rect 132874 442046 132970 442102
rect 133026 442046 133094 442102
rect 133150 442046 133218 442102
rect 133274 442046 133342 442102
rect 133398 442046 133494 442102
rect 132874 441978 133494 442046
rect 132874 441922 132970 441978
rect 133026 441922 133094 441978
rect 133150 441922 133218 441978
rect 133274 441922 133342 441978
rect 133398 441922 133494 441978
rect 132874 424350 133494 441922
rect 132874 424294 132970 424350
rect 133026 424294 133094 424350
rect 133150 424294 133218 424350
rect 133274 424294 133342 424350
rect 133398 424294 133494 424350
rect 132874 424226 133494 424294
rect 132874 424170 132970 424226
rect 133026 424170 133094 424226
rect 133150 424170 133218 424226
rect 133274 424170 133342 424226
rect 133398 424170 133494 424226
rect 132874 424102 133494 424170
rect 132874 424046 132970 424102
rect 133026 424046 133094 424102
rect 133150 424046 133218 424102
rect 133274 424046 133342 424102
rect 133398 424046 133494 424102
rect 132874 423978 133494 424046
rect 132874 423922 132970 423978
rect 133026 423922 133094 423978
rect 133150 423922 133218 423978
rect 133274 423922 133342 423978
rect 133398 423922 133494 423978
rect 132874 406350 133494 423922
rect 132874 406294 132970 406350
rect 133026 406294 133094 406350
rect 133150 406294 133218 406350
rect 133274 406294 133342 406350
rect 133398 406294 133494 406350
rect 132874 406226 133494 406294
rect 132874 406170 132970 406226
rect 133026 406170 133094 406226
rect 133150 406170 133218 406226
rect 133274 406170 133342 406226
rect 133398 406170 133494 406226
rect 132874 406102 133494 406170
rect 132874 406046 132970 406102
rect 133026 406046 133094 406102
rect 133150 406046 133218 406102
rect 133274 406046 133342 406102
rect 133398 406046 133494 406102
rect 132874 405978 133494 406046
rect 132874 405922 132970 405978
rect 133026 405922 133094 405978
rect 133150 405922 133218 405978
rect 133274 405922 133342 405978
rect 133398 405922 133494 405978
rect 132874 388350 133494 405922
rect 132874 388294 132970 388350
rect 133026 388294 133094 388350
rect 133150 388294 133218 388350
rect 133274 388294 133342 388350
rect 133398 388294 133494 388350
rect 132874 388226 133494 388294
rect 132874 388170 132970 388226
rect 133026 388170 133094 388226
rect 133150 388170 133218 388226
rect 133274 388170 133342 388226
rect 133398 388170 133494 388226
rect 132874 388102 133494 388170
rect 132874 388046 132970 388102
rect 133026 388046 133094 388102
rect 133150 388046 133218 388102
rect 133274 388046 133342 388102
rect 133398 388046 133494 388102
rect 132874 387978 133494 388046
rect 132874 387922 132970 387978
rect 133026 387922 133094 387978
rect 133150 387922 133218 387978
rect 133274 387922 133342 387978
rect 133398 387922 133494 387978
rect 132874 370350 133494 387922
rect 132874 370294 132970 370350
rect 133026 370294 133094 370350
rect 133150 370294 133218 370350
rect 133274 370294 133342 370350
rect 133398 370294 133494 370350
rect 132874 370226 133494 370294
rect 132874 370170 132970 370226
rect 133026 370170 133094 370226
rect 133150 370170 133218 370226
rect 133274 370170 133342 370226
rect 133398 370170 133494 370226
rect 132874 370102 133494 370170
rect 132874 370046 132970 370102
rect 133026 370046 133094 370102
rect 133150 370046 133218 370102
rect 133274 370046 133342 370102
rect 133398 370046 133494 370102
rect 132874 369978 133494 370046
rect 132874 369922 132970 369978
rect 133026 369922 133094 369978
rect 133150 369922 133218 369978
rect 133274 369922 133342 369978
rect 133398 369922 133494 369978
rect 132874 352350 133494 369922
rect 132874 352294 132970 352350
rect 133026 352294 133094 352350
rect 133150 352294 133218 352350
rect 133274 352294 133342 352350
rect 133398 352294 133494 352350
rect 132874 352226 133494 352294
rect 132874 352170 132970 352226
rect 133026 352170 133094 352226
rect 133150 352170 133218 352226
rect 133274 352170 133342 352226
rect 133398 352170 133494 352226
rect 132874 352102 133494 352170
rect 132874 352046 132970 352102
rect 133026 352046 133094 352102
rect 133150 352046 133218 352102
rect 133274 352046 133342 352102
rect 133398 352046 133494 352102
rect 132874 351978 133494 352046
rect 132874 351922 132970 351978
rect 133026 351922 133094 351978
rect 133150 351922 133218 351978
rect 133274 351922 133342 351978
rect 133398 351922 133494 351978
rect 132874 334350 133494 351922
rect 132874 334294 132970 334350
rect 133026 334294 133094 334350
rect 133150 334294 133218 334350
rect 133274 334294 133342 334350
rect 133398 334294 133494 334350
rect 132874 334226 133494 334294
rect 132874 334170 132970 334226
rect 133026 334170 133094 334226
rect 133150 334170 133218 334226
rect 133274 334170 133342 334226
rect 133398 334170 133494 334226
rect 132874 334102 133494 334170
rect 132874 334046 132970 334102
rect 133026 334046 133094 334102
rect 133150 334046 133218 334102
rect 133274 334046 133342 334102
rect 133398 334046 133494 334102
rect 132874 333978 133494 334046
rect 132874 333922 132970 333978
rect 133026 333922 133094 333978
rect 133150 333922 133218 333978
rect 133274 333922 133342 333978
rect 133398 333922 133494 333978
rect 132874 316350 133494 333922
rect 132874 316294 132970 316350
rect 133026 316294 133094 316350
rect 133150 316294 133218 316350
rect 133274 316294 133342 316350
rect 133398 316294 133494 316350
rect 132874 316226 133494 316294
rect 132874 316170 132970 316226
rect 133026 316170 133094 316226
rect 133150 316170 133218 316226
rect 133274 316170 133342 316226
rect 133398 316170 133494 316226
rect 132874 316102 133494 316170
rect 132874 316046 132970 316102
rect 133026 316046 133094 316102
rect 133150 316046 133218 316102
rect 133274 316046 133342 316102
rect 133398 316046 133494 316102
rect 132874 315978 133494 316046
rect 132874 315922 132970 315978
rect 133026 315922 133094 315978
rect 133150 315922 133218 315978
rect 133274 315922 133342 315978
rect 133398 315922 133494 315978
rect 132874 298350 133494 315922
rect 132874 298294 132970 298350
rect 133026 298294 133094 298350
rect 133150 298294 133218 298350
rect 133274 298294 133342 298350
rect 133398 298294 133494 298350
rect 132874 298226 133494 298294
rect 132874 298170 132970 298226
rect 133026 298170 133094 298226
rect 133150 298170 133218 298226
rect 133274 298170 133342 298226
rect 133398 298170 133494 298226
rect 132874 298102 133494 298170
rect 132874 298046 132970 298102
rect 133026 298046 133094 298102
rect 133150 298046 133218 298102
rect 133274 298046 133342 298102
rect 133398 298046 133494 298102
rect 132874 297978 133494 298046
rect 132874 297922 132970 297978
rect 133026 297922 133094 297978
rect 133150 297922 133218 297978
rect 133274 297922 133342 297978
rect 133398 297922 133494 297978
rect 132874 280350 133494 297922
rect 132874 280294 132970 280350
rect 133026 280294 133094 280350
rect 133150 280294 133218 280350
rect 133274 280294 133342 280350
rect 133398 280294 133494 280350
rect 132874 280226 133494 280294
rect 132874 280170 132970 280226
rect 133026 280170 133094 280226
rect 133150 280170 133218 280226
rect 133274 280170 133342 280226
rect 133398 280170 133494 280226
rect 132874 280102 133494 280170
rect 132874 280046 132970 280102
rect 133026 280046 133094 280102
rect 133150 280046 133218 280102
rect 133274 280046 133342 280102
rect 133398 280046 133494 280102
rect 132874 279978 133494 280046
rect 132874 279922 132970 279978
rect 133026 279922 133094 279978
rect 133150 279922 133218 279978
rect 133274 279922 133342 279978
rect 133398 279922 133494 279978
rect 132874 262350 133494 279922
rect 132874 262294 132970 262350
rect 133026 262294 133094 262350
rect 133150 262294 133218 262350
rect 133274 262294 133342 262350
rect 133398 262294 133494 262350
rect 132874 262226 133494 262294
rect 132874 262170 132970 262226
rect 133026 262170 133094 262226
rect 133150 262170 133218 262226
rect 133274 262170 133342 262226
rect 133398 262170 133494 262226
rect 132874 262102 133494 262170
rect 132874 262046 132970 262102
rect 133026 262046 133094 262102
rect 133150 262046 133218 262102
rect 133274 262046 133342 262102
rect 133398 262046 133494 262102
rect 132874 261978 133494 262046
rect 132874 261922 132970 261978
rect 133026 261922 133094 261978
rect 133150 261922 133218 261978
rect 133274 261922 133342 261978
rect 133398 261922 133494 261978
rect 132874 244350 133494 261922
rect 132874 244294 132970 244350
rect 133026 244294 133094 244350
rect 133150 244294 133218 244350
rect 133274 244294 133342 244350
rect 133398 244294 133494 244350
rect 132874 244226 133494 244294
rect 132874 244170 132970 244226
rect 133026 244170 133094 244226
rect 133150 244170 133218 244226
rect 133274 244170 133342 244226
rect 133398 244170 133494 244226
rect 132874 244102 133494 244170
rect 132874 244046 132970 244102
rect 133026 244046 133094 244102
rect 133150 244046 133218 244102
rect 133274 244046 133342 244102
rect 133398 244046 133494 244102
rect 132874 243978 133494 244046
rect 132874 243922 132970 243978
rect 133026 243922 133094 243978
rect 133150 243922 133218 243978
rect 133274 243922 133342 243978
rect 133398 243922 133494 243978
rect 132874 226350 133494 243922
rect 147154 597212 147774 598268
rect 147154 597156 147250 597212
rect 147306 597156 147374 597212
rect 147430 597156 147498 597212
rect 147554 597156 147622 597212
rect 147678 597156 147774 597212
rect 147154 597088 147774 597156
rect 147154 597032 147250 597088
rect 147306 597032 147374 597088
rect 147430 597032 147498 597088
rect 147554 597032 147622 597088
rect 147678 597032 147774 597088
rect 147154 596964 147774 597032
rect 147154 596908 147250 596964
rect 147306 596908 147374 596964
rect 147430 596908 147498 596964
rect 147554 596908 147622 596964
rect 147678 596908 147774 596964
rect 147154 596840 147774 596908
rect 147154 596784 147250 596840
rect 147306 596784 147374 596840
rect 147430 596784 147498 596840
rect 147554 596784 147622 596840
rect 147678 596784 147774 596840
rect 147154 580350 147774 596784
rect 147154 580294 147250 580350
rect 147306 580294 147374 580350
rect 147430 580294 147498 580350
rect 147554 580294 147622 580350
rect 147678 580294 147774 580350
rect 147154 580226 147774 580294
rect 147154 580170 147250 580226
rect 147306 580170 147374 580226
rect 147430 580170 147498 580226
rect 147554 580170 147622 580226
rect 147678 580170 147774 580226
rect 147154 580102 147774 580170
rect 147154 580046 147250 580102
rect 147306 580046 147374 580102
rect 147430 580046 147498 580102
rect 147554 580046 147622 580102
rect 147678 580046 147774 580102
rect 147154 579978 147774 580046
rect 147154 579922 147250 579978
rect 147306 579922 147374 579978
rect 147430 579922 147498 579978
rect 147554 579922 147622 579978
rect 147678 579922 147774 579978
rect 147154 562350 147774 579922
rect 147154 562294 147250 562350
rect 147306 562294 147374 562350
rect 147430 562294 147498 562350
rect 147554 562294 147622 562350
rect 147678 562294 147774 562350
rect 147154 562226 147774 562294
rect 147154 562170 147250 562226
rect 147306 562170 147374 562226
rect 147430 562170 147498 562226
rect 147554 562170 147622 562226
rect 147678 562170 147774 562226
rect 147154 562102 147774 562170
rect 147154 562046 147250 562102
rect 147306 562046 147374 562102
rect 147430 562046 147498 562102
rect 147554 562046 147622 562102
rect 147678 562046 147774 562102
rect 147154 561978 147774 562046
rect 147154 561922 147250 561978
rect 147306 561922 147374 561978
rect 147430 561922 147498 561978
rect 147554 561922 147622 561978
rect 147678 561922 147774 561978
rect 147154 544350 147774 561922
rect 147154 544294 147250 544350
rect 147306 544294 147374 544350
rect 147430 544294 147498 544350
rect 147554 544294 147622 544350
rect 147678 544294 147774 544350
rect 147154 544226 147774 544294
rect 147154 544170 147250 544226
rect 147306 544170 147374 544226
rect 147430 544170 147498 544226
rect 147554 544170 147622 544226
rect 147678 544170 147774 544226
rect 147154 544102 147774 544170
rect 147154 544046 147250 544102
rect 147306 544046 147374 544102
rect 147430 544046 147498 544102
rect 147554 544046 147622 544102
rect 147678 544046 147774 544102
rect 147154 543978 147774 544046
rect 147154 543922 147250 543978
rect 147306 543922 147374 543978
rect 147430 543922 147498 543978
rect 147554 543922 147622 543978
rect 147678 543922 147774 543978
rect 147154 526350 147774 543922
rect 147154 526294 147250 526350
rect 147306 526294 147374 526350
rect 147430 526294 147498 526350
rect 147554 526294 147622 526350
rect 147678 526294 147774 526350
rect 147154 526226 147774 526294
rect 147154 526170 147250 526226
rect 147306 526170 147374 526226
rect 147430 526170 147498 526226
rect 147554 526170 147622 526226
rect 147678 526170 147774 526226
rect 147154 526102 147774 526170
rect 147154 526046 147250 526102
rect 147306 526046 147374 526102
rect 147430 526046 147498 526102
rect 147554 526046 147622 526102
rect 147678 526046 147774 526102
rect 147154 525978 147774 526046
rect 147154 525922 147250 525978
rect 147306 525922 147374 525978
rect 147430 525922 147498 525978
rect 147554 525922 147622 525978
rect 147678 525922 147774 525978
rect 147154 508350 147774 525922
rect 147154 508294 147250 508350
rect 147306 508294 147374 508350
rect 147430 508294 147498 508350
rect 147554 508294 147622 508350
rect 147678 508294 147774 508350
rect 147154 508226 147774 508294
rect 147154 508170 147250 508226
rect 147306 508170 147374 508226
rect 147430 508170 147498 508226
rect 147554 508170 147622 508226
rect 147678 508170 147774 508226
rect 147154 508102 147774 508170
rect 147154 508046 147250 508102
rect 147306 508046 147374 508102
rect 147430 508046 147498 508102
rect 147554 508046 147622 508102
rect 147678 508046 147774 508102
rect 147154 507978 147774 508046
rect 147154 507922 147250 507978
rect 147306 507922 147374 507978
rect 147430 507922 147498 507978
rect 147554 507922 147622 507978
rect 147678 507922 147774 507978
rect 147154 490350 147774 507922
rect 147154 490294 147250 490350
rect 147306 490294 147374 490350
rect 147430 490294 147498 490350
rect 147554 490294 147622 490350
rect 147678 490294 147774 490350
rect 147154 490226 147774 490294
rect 147154 490170 147250 490226
rect 147306 490170 147374 490226
rect 147430 490170 147498 490226
rect 147554 490170 147622 490226
rect 147678 490170 147774 490226
rect 147154 490102 147774 490170
rect 147154 490046 147250 490102
rect 147306 490046 147374 490102
rect 147430 490046 147498 490102
rect 147554 490046 147622 490102
rect 147678 490046 147774 490102
rect 147154 489978 147774 490046
rect 147154 489922 147250 489978
rect 147306 489922 147374 489978
rect 147430 489922 147498 489978
rect 147554 489922 147622 489978
rect 147678 489922 147774 489978
rect 147154 472350 147774 489922
rect 147154 472294 147250 472350
rect 147306 472294 147374 472350
rect 147430 472294 147498 472350
rect 147554 472294 147622 472350
rect 147678 472294 147774 472350
rect 147154 472226 147774 472294
rect 147154 472170 147250 472226
rect 147306 472170 147374 472226
rect 147430 472170 147498 472226
rect 147554 472170 147622 472226
rect 147678 472170 147774 472226
rect 147154 472102 147774 472170
rect 147154 472046 147250 472102
rect 147306 472046 147374 472102
rect 147430 472046 147498 472102
rect 147554 472046 147622 472102
rect 147678 472046 147774 472102
rect 147154 471978 147774 472046
rect 147154 471922 147250 471978
rect 147306 471922 147374 471978
rect 147430 471922 147498 471978
rect 147554 471922 147622 471978
rect 147678 471922 147774 471978
rect 147154 454350 147774 471922
rect 147154 454294 147250 454350
rect 147306 454294 147374 454350
rect 147430 454294 147498 454350
rect 147554 454294 147622 454350
rect 147678 454294 147774 454350
rect 147154 454226 147774 454294
rect 147154 454170 147250 454226
rect 147306 454170 147374 454226
rect 147430 454170 147498 454226
rect 147554 454170 147622 454226
rect 147678 454170 147774 454226
rect 147154 454102 147774 454170
rect 147154 454046 147250 454102
rect 147306 454046 147374 454102
rect 147430 454046 147498 454102
rect 147554 454046 147622 454102
rect 147678 454046 147774 454102
rect 147154 453978 147774 454046
rect 147154 453922 147250 453978
rect 147306 453922 147374 453978
rect 147430 453922 147498 453978
rect 147554 453922 147622 453978
rect 147678 453922 147774 453978
rect 147154 436350 147774 453922
rect 147154 436294 147250 436350
rect 147306 436294 147374 436350
rect 147430 436294 147498 436350
rect 147554 436294 147622 436350
rect 147678 436294 147774 436350
rect 147154 436226 147774 436294
rect 147154 436170 147250 436226
rect 147306 436170 147374 436226
rect 147430 436170 147498 436226
rect 147554 436170 147622 436226
rect 147678 436170 147774 436226
rect 147154 436102 147774 436170
rect 147154 436046 147250 436102
rect 147306 436046 147374 436102
rect 147430 436046 147498 436102
rect 147554 436046 147622 436102
rect 147678 436046 147774 436102
rect 147154 435978 147774 436046
rect 147154 435922 147250 435978
rect 147306 435922 147374 435978
rect 147430 435922 147498 435978
rect 147554 435922 147622 435978
rect 147678 435922 147774 435978
rect 147154 418350 147774 435922
rect 147154 418294 147250 418350
rect 147306 418294 147374 418350
rect 147430 418294 147498 418350
rect 147554 418294 147622 418350
rect 147678 418294 147774 418350
rect 147154 418226 147774 418294
rect 147154 418170 147250 418226
rect 147306 418170 147374 418226
rect 147430 418170 147498 418226
rect 147554 418170 147622 418226
rect 147678 418170 147774 418226
rect 147154 418102 147774 418170
rect 147154 418046 147250 418102
rect 147306 418046 147374 418102
rect 147430 418046 147498 418102
rect 147554 418046 147622 418102
rect 147678 418046 147774 418102
rect 147154 417978 147774 418046
rect 147154 417922 147250 417978
rect 147306 417922 147374 417978
rect 147430 417922 147498 417978
rect 147554 417922 147622 417978
rect 147678 417922 147774 417978
rect 147154 400350 147774 417922
rect 147154 400294 147250 400350
rect 147306 400294 147374 400350
rect 147430 400294 147498 400350
rect 147554 400294 147622 400350
rect 147678 400294 147774 400350
rect 147154 400226 147774 400294
rect 147154 400170 147250 400226
rect 147306 400170 147374 400226
rect 147430 400170 147498 400226
rect 147554 400170 147622 400226
rect 147678 400170 147774 400226
rect 147154 400102 147774 400170
rect 147154 400046 147250 400102
rect 147306 400046 147374 400102
rect 147430 400046 147498 400102
rect 147554 400046 147622 400102
rect 147678 400046 147774 400102
rect 147154 399978 147774 400046
rect 147154 399922 147250 399978
rect 147306 399922 147374 399978
rect 147430 399922 147498 399978
rect 147554 399922 147622 399978
rect 147678 399922 147774 399978
rect 147154 382350 147774 399922
rect 147154 382294 147250 382350
rect 147306 382294 147374 382350
rect 147430 382294 147498 382350
rect 147554 382294 147622 382350
rect 147678 382294 147774 382350
rect 147154 382226 147774 382294
rect 147154 382170 147250 382226
rect 147306 382170 147374 382226
rect 147430 382170 147498 382226
rect 147554 382170 147622 382226
rect 147678 382170 147774 382226
rect 147154 382102 147774 382170
rect 147154 382046 147250 382102
rect 147306 382046 147374 382102
rect 147430 382046 147498 382102
rect 147554 382046 147622 382102
rect 147678 382046 147774 382102
rect 147154 381978 147774 382046
rect 147154 381922 147250 381978
rect 147306 381922 147374 381978
rect 147430 381922 147498 381978
rect 147554 381922 147622 381978
rect 147678 381922 147774 381978
rect 147154 364350 147774 381922
rect 147154 364294 147250 364350
rect 147306 364294 147374 364350
rect 147430 364294 147498 364350
rect 147554 364294 147622 364350
rect 147678 364294 147774 364350
rect 147154 364226 147774 364294
rect 147154 364170 147250 364226
rect 147306 364170 147374 364226
rect 147430 364170 147498 364226
rect 147554 364170 147622 364226
rect 147678 364170 147774 364226
rect 147154 364102 147774 364170
rect 147154 364046 147250 364102
rect 147306 364046 147374 364102
rect 147430 364046 147498 364102
rect 147554 364046 147622 364102
rect 147678 364046 147774 364102
rect 147154 363978 147774 364046
rect 147154 363922 147250 363978
rect 147306 363922 147374 363978
rect 147430 363922 147498 363978
rect 147554 363922 147622 363978
rect 147678 363922 147774 363978
rect 147154 346350 147774 363922
rect 147154 346294 147250 346350
rect 147306 346294 147374 346350
rect 147430 346294 147498 346350
rect 147554 346294 147622 346350
rect 147678 346294 147774 346350
rect 147154 346226 147774 346294
rect 147154 346170 147250 346226
rect 147306 346170 147374 346226
rect 147430 346170 147498 346226
rect 147554 346170 147622 346226
rect 147678 346170 147774 346226
rect 147154 346102 147774 346170
rect 147154 346046 147250 346102
rect 147306 346046 147374 346102
rect 147430 346046 147498 346102
rect 147554 346046 147622 346102
rect 147678 346046 147774 346102
rect 147154 345978 147774 346046
rect 147154 345922 147250 345978
rect 147306 345922 147374 345978
rect 147430 345922 147498 345978
rect 147554 345922 147622 345978
rect 147678 345922 147774 345978
rect 147154 328350 147774 345922
rect 147154 328294 147250 328350
rect 147306 328294 147374 328350
rect 147430 328294 147498 328350
rect 147554 328294 147622 328350
rect 147678 328294 147774 328350
rect 147154 328226 147774 328294
rect 147154 328170 147250 328226
rect 147306 328170 147374 328226
rect 147430 328170 147498 328226
rect 147554 328170 147622 328226
rect 147678 328170 147774 328226
rect 147154 328102 147774 328170
rect 147154 328046 147250 328102
rect 147306 328046 147374 328102
rect 147430 328046 147498 328102
rect 147554 328046 147622 328102
rect 147678 328046 147774 328102
rect 147154 327978 147774 328046
rect 147154 327922 147250 327978
rect 147306 327922 147374 327978
rect 147430 327922 147498 327978
rect 147554 327922 147622 327978
rect 147678 327922 147774 327978
rect 147154 310350 147774 327922
rect 147154 310294 147250 310350
rect 147306 310294 147374 310350
rect 147430 310294 147498 310350
rect 147554 310294 147622 310350
rect 147678 310294 147774 310350
rect 147154 310226 147774 310294
rect 147154 310170 147250 310226
rect 147306 310170 147374 310226
rect 147430 310170 147498 310226
rect 147554 310170 147622 310226
rect 147678 310170 147774 310226
rect 147154 310102 147774 310170
rect 147154 310046 147250 310102
rect 147306 310046 147374 310102
rect 147430 310046 147498 310102
rect 147554 310046 147622 310102
rect 147678 310046 147774 310102
rect 147154 309978 147774 310046
rect 147154 309922 147250 309978
rect 147306 309922 147374 309978
rect 147430 309922 147498 309978
rect 147554 309922 147622 309978
rect 147678 309922 147774 309978
rect 147154 292350 147774 309922
rect 147154 292294 147250 292350
rect 147306 292294 147374 292350
rect 147430 292294 147498 292350
rect 147554 292294 147622 292350
rect 147678 292294 147774 292350
rect 147154 292226 147774 292294
rect 147154 292170 147250 292226
rect 147306 292170 147374 292226
rect 147430 292170 147498 292226
rect 147554 292170 147622 292226
rect 147678 292170 147774 292226
rect 147154 292102 147774 292170
rect 147154 292046 147250 292102
rect 147306 292046 147374 292102
rect 147430 292046 147498 292102
rect 147554 292046 147622 292102
rect 147678 292046 147774 292102
rect 147154 291978 147774 292046
rect 147154 291922 147250 291978
rect 147306 291922 147374 291978
rect 147430 291922 147498 291978
rect 147554 291922 147622 291978
rect 147678 291922 147774 291978
rect 147154 274350 147774 291922
rect 147154 274294 147250 274350
rect 147306 274294 147374 274350
rect 147430 274294 147498 274350
rect 147554 274294 147622 274350
rect 147678 274294 147774 274350
rect 147154 274226 147774 274294
rect 147154 274170 147250 274226
rect 147306 274170 147374 274226
rect 147430 274170 147498 274226
rect 147554 274170 147622 274226
rect 147678 274170 147774 274226
rect 147154 274102 147774 274170
rect 147154 274046 147250 274102
rect 147306 274046 147374 274102
rect 147430 274046 147498 274102
rect 147554 274046 147622 274102
rect 147678 274046 147774 274102
rect 147154 273978 147774 274046
rect 147154 273922 147250 273978
rect 147306 273922 147374 273978
rect 147430 273922 147498 273978
rect 147554 273922 147622 273978
rect 147678 273922 147774 273978
rect 147154 256350 147774 273922
rect 147154 256294 147250 256350
rect 147306 256294 147374 256350
rect 147430 256294 147498 256350
rect 147554 256294 147622 256350
rect 147678 256294 147774 256350
rect 147154 256226 147774 256294
rect 147154 256170 147250 256226
rect 147306 256170 147374 256226
rect 147430 256170 147498 256226
rect 147554 256170 147622 256226
rect 147678 256170 147774 256226
rect 147154 256102 147774 256170
rect 147154 256046 147250 256102
rect 147306 256046 147374 256102
rect 147430 256046 147498 256102
rect 147554 256046 147622 256102
rect 147678 256046 147774 256102
rect 147154 255978 147774 256046
rect 147154 255922 147250 255978
rect 147306 255922 147374 255978
rect 147430 255922 147498 255978
rect 147554 255922 147622 255978
rect 147678 255922 147774 255978
rect 147154 238350 147774 255922
rect 147154 238294 147250 238350
rect 147306 238294 147374 238350
rect 147430 238294 147498 238350
rect 147554 238294 147622 238350
rect 147678 238294 147774 238350
rect 147154 238226 147774 238294
rect 147154 238170 147250 238226
rect 147306 238170 147374 238226
rect 147430 238170 147498 238226
rect 147554 238170 147622 238226
rect 147678 238170 147774 238226
rect 147154 238102 147774 238170
rect 147154 238046 147250 238102
rect 147306 238046 147374 238102
rect 147430 238046 147498 238102
rect 147554 238046 147622 238102
rect 147678 238046 147774 238102
rect 147154 237978 147774 238046
rect 147154 237922 147250 237978
rect 147306 237922 147374 237978
rect 147430 237922 147498 237978
rect 147554 237922 147622 237978
rect 147678 237922 147774 237978
rect 132874 226294 132970 226350
rect 133026 226294 133094 226350
rect 133150 226294 133218 226350
rect 133274 226294 133342 226350
rect 133398 226294 133494 226350
rect 132874 226226 133494 226294
rect 132874 226170 132970 226226
rect 133026 226170 133094 226226
rect 133150 226170 133218 226226
rect 133274 226170 133342 226226
rect 133398 226170 133494 226226
rect 132874 226102 133494 226170
rect 132874 226046 132970 226102
rect 133026 226046 133094 226102
rect 133150 226046 133218 226102
rect 133274 226046 133342 226102
rect 133398 226046 133494 226102
rect 132874 225978 133494 226046
rect 132874 225922 132970 225978
rect 133026 225922 133094 225978
rect 133150 225922 133218 225978
rect 133274 225922 133342 225978
rect 133398 225922 133494 225978
rect 132874 219134 133494 225922
rect 141248 226350 141568 226384
rect 141248 226294 141318 226350
rect 141374 226294 141442 226350
rect 141498 226294 141568 226350
rect 141248 226226 141568 226294
rect 141248 226170 141318 226226
rect 141374 226170 141442 226226
rect 141498 226170 141568 226226
rect 141248 226102 141568 226170
rect 141248 226046 141318 226102
rect 141374 226046 141442 226102
rect 141498 226046 141568 226102
rect 141248 225978 141568 226046
rect 141248 225922 141318 225978
rect 141374 225922 141442 225978
rect 141498 225922 141568 225978
rect 141248 225888 141568 225922
rect 147154 220350 147774 237922
rect 147154 220294 147250 220350
rect 147306 220294 147374 220350
rect 147430 220294 147498 220350
rect 147554 220294 147622 220350
rect 147678 220294 147774 220350
rect 147154 220226 147774 220294
rect 147154 220170 147250 220226
rect 147306 220170 147374 220226
rect 147430 220170 147498 220226
rect 147554 220170 147622 220226
rect 147678 220170 147774 220226
rect 147154 220102 147774 220170
rect 147154 220046 147250 220102
rect 147306 220046 147374 220102
rect 147430 220046 147498 220102
rect 147554 220046 147622 220102
rect 147678 220046 147774 220102
rect 147154 219978 147774 220046
rect 147154 219922 147250 219978
rect 147306 219922 147374 219978
rect 147430 219922 147498 219978
rect 147554 219922 147622 219978
rect 147678 219922 147774 219978
rect 147154 219134 147774 219922
rect 150874 598172 151494 598268
rect 150874 598116 150970 598172
rect 151026 598116 151094 598172
rect 151150 598116 151218 598172
rect 151274 598116 151342 598172
rect 151398 598116 151494 598172
rect 150874 598048 151494 598116
rect 150874 597992 150970 598048
rect 151026 597992 151094 598048
rect 151150 597992 151218 598048
rect 151274 597992 151342 598048
rect 151398 597992 151494 598048
rect 150874 597924 151494 597992
rect 150874 597868 150970 597924
rect 151026 597868 151094 597924
rect 151150 597868 151218 597924
rect 151274 597868 151342 597924
rect 151398 597868 151494 597924
rect 150874 597800 151494 597868
rect 150874 597744 150970 597800
rect 151026 597744 151094 597800
rect 151150 597744 151218 597800
rect 151274 597744 151342 597800
rect 151398 597744 151494 597800
rect 150874 586350 151494 597744
rect 150874 586294 150970 586350
rect 151026 586294 151094 586350
rect 151150 586294 151218 586350
rect 151274 586294 151342 586350
rect 151398 586294 151494 586350
rect 150874 586226 151494 586294
rect 150874 586170 150970 586226
rect 151026 586170 151094 586226
rect 151150 586170 151218 586226
rect 151274 586170 151342 586226
rect 151398 586170 151494 586226
rect 150874 586102 151494 586170
rect 150874 586046 150970 586102
rect 151026 586046 151094 586102
rect 151150 586046 151218 586102
rect 151274 586046 151342 586102
rect 151398 586046 151494 586102
rect 150874 585978 151494 586046
rect 150874 585922 150970 585978
rect 151026 585922 151094 585978
rect 151150 585922 151218 585978
rect 151274 585922 151342 585978
rect 151398 585922 151494 585978
rect 150874 568350 151494 585922
rect 150874 568294 150970 568350
rect 151026 568294 151094 568350
rect 151150 568294 151218 568350
rect 151274 568294 151342 568350
rect 151398 568294 151494 568350
rect 150874 568226 151494 568294
rect 150874 568170 150970 568226
rect 151026 568170 151094 568226
rect 151150 568170 151218 568226
rect 151274 568170 151342 568226
rect 151398 568170 151494 568226
rect 150874 568102 151494 568170
rect 150874 568046 150970 568102
rect 151026 568046 151094 568102
rect 151150 568046 151218 568102
rect 151274 568046 151342 568102
rect 151398 568046 151494 568102
rect 150874 567978 151494 568046
rect 150874 567922 150970 567978
rect 151026 567922 151094 567978
rect 151150 567922 151218 567978
rect 151274 567922 151342 567978
rect 151398 567922 151494 567978
rect 150874 550350 151494 567922
rect 150874 550294 150970 550350
rect 151026 550294 151094 550350
rect 151150 550294 151218 550350
rect 151274 550294 151342 550350
rect 151398 550294 151494 550350
rect 150874 550226 151494 550294
rect 150874 550170 150970 550226
rect 151026 550170 151094 550226
rect 151150 550170 151218 550226
rect 151274 550170 151342 550226
rect 151398 550170 151494 550226
rect 150874 550102 151494 550170
rect 150874 550046 150970 550102
rect 151026 550046 151094 550102
rect 151150 550046 151218 550102
rect 151274 550046 151342 550102
rect 151398 550046 151494 550102
rect 150874 549978 151494 550046
rect 150874 549922 150970 549978
rect 151026 549922 151094 549978
rect 151150 549922 151218 549978
rect 151274 549922 151342 549978
rect 151398 549922 151494 549978
rect 150874 532350 151494 549922
rect 150874 532294 150970 532350
rect 151026 532294 151094 532350
rect 151150 532294 151218 532350
rect 151274 532294 151342 532350
rect 151398 532294 151494 532350
rect 150874 532226 151494 532294
rect 150874 532170 150970 532226
rect 151026 532170 151094 532226
rect 151150 532170 151218 532226
rect 151274 532170 151342 532226
rect 151398 532170 151494 532226
rect 150874 532102 151494 532170
rect 150874 532046 150970 532102
rect 151026 532046 151094 532102
rect 151150 532046 151218 532102
rect 151274 532046 151342 532102
rect 151398 532046 151494 532102
rect 150874 531978 151494 532046
rect 150874 531922 150970 531978
rect 151026 531922 151094 531978
rect 151150 531922 151218 531978
rect 151274 531922 151342 531978
rect 151398 531922 151494 531978
rect 150874 514350 151494 531922
rect 150874 514294 150970 514350
rect 151026 514294 151094 514350
rect 151150 514294 151218 514350
rect 151274 514294 151342 514350
rect 151398 514294 151494 514350
rect 150874 514226 151494 514294
rect 150874 514170 150970 514226
rect 151026 514170 151094 514226
rect 151150 514170 151218 514226
rect 151274 514170 151342 514226
rect 151398 514170 151494 514226
rect 150874 514102 151494 514170
rect 150874 514046 150970 514102
rect 151026 514046 151094 514102
rect 151150 514046 151218 514102
rect 151274 514046 151342 514102
rect 151398 514046 151494 514102
rect 150874 513978 151494 514046
rect 150874 513922 150970 513978
rect 151026 513922 151094 513978
rect 151150 513922 151218 513978
rect 151274 513922 151342 513978
rect 151398 513922 151494 513978
rect 150874 496350 151494 513922
rect 150874 496294 150970 496350
rect 151026 496294 151094 496350
rect 151150 496294 151218 496350
rect 151274 496294 151342 496350
rect 151398 496294 151494 496350
rect 150874 496226 151494 496294
rect 150874 496170 150970 496226
rect 151026 496170 151094 496226
rect 151150 496170 151218 496226
rect 151274 496170 151342 496226
rect 151398 496170 151494 496226
rect 150874 496102 151494 496170
rect 150874 496046 150970 496102
rect 151026 496046 151094 496102
rect 151150 496046 151218 496102
rect 151274 496046 151342 496102
rect 151398 496046 151494 496102
rect 150874 495978 151494 496046
rect 150874 495922 150970 495978
rect 151026 495922 151094 495978
rect 151150 495922 151218 495978
rect 151274 495922 151342 495978
rect 151398 495922 151494 495978
rect 150874 478350 151494 495922
rect 150874 478294 150970 478350
rect 151026 478294 151094 478350
rect 151150 478294 151218 478350
rect 151274 478294 151342 478350
rect 151398 478294 151494 478350
rect 150874 478226 151494 478294
rect 150874 478170 150970 478226
rect 151026 478170 151094 478226
rect 151150 478170 151218 478226
rect 151274 478170 151342 478226
rect 151398 478170 151494 478226
rect 150874 478102 151494 478170
rect 150874 478046 150970 478102
rect 151026 478046 151094 478102
rect 151150 478046 151218 478102
rect 151274 478046 151342 478102
rect 151398 478046 151494 478102
rect 150874 477978 151494 478046
rect 150874 477922 150970 477978
rect 151026 477922 151094 477978
rect 151150 477922 151218 477978
rect 151274 477922 151342 477978
rect 151398 477922 151494 477978
rect 150874 460350 151494 477922
rect 150874 460294 150970 460350
rect 151026 460294 151094 460350
rect 151150 460294 151218 460350
rect 151274 460294 151342 460350
rect 151398 460294 151494 460350
rect 150874 460226 151494 460294
rect 150874 460170 150970 460226
rect 151026 460170 151094 460226
rect 151150 460170 151218 460226
rect 151274 460170 151342 460226
rect 151398 460170 151494 460226
rect 150874 460102 151494 460170
rect 150874 460046 150970 460102
rect 151026 460046 151094 460102
rect 151150 460046 151218 460102
rect 151274 460046 151342 460102
rect 151398 460046 151494 460102
rect 150874 459978 151494 460046
rect 150874 459922 150970 459978
rect 151026 459922 151094 459978
rect 151150 459922 151218 459978
rect 151274 459922 151342 459978
rect 151398 459922 151494 459978
rect 150874 442350 151494 459922
rect 150874 442294 150970 442350
rect 151026 442294 151094 442350
rect 151150 442294 151218 442350
rect 151274 442294 151342 442350
rect 151398 442294 151494 442350
rect 150874 442226 151494 442294
rect 150874 442170 150970 442226
rect 151026 442170 151094 442226
rect 151150 442170 151218 442226
rect 151274 442170 151342 442226
rect 151398 442170 151494 442226
rect 150874 442102 151494 442170
rect 150874 442046 150970 442102
rect 151026 442046 151094 442102
rect 151150 442046 151218 442102
rect 151274 442046 151342 442102
rect 151398 442046 151494 442102
rect 150874 441978 151494 442046
rect 150874 441922 150970 441978
rect 151026 441922 151094 441978
rect 151150 441922 151218 441978
rect 151274 441922 151342 441978
rect 151398 441922 151494 441978
rect 150874 424350 151494 441922
rect 150874 424294 150970 424350
rect 151026 424294 151094 424350
rect 151150 424294 151218 424350
rect 151274 424294 151342 424350
rect 151398 424294 151494 424350
rect 150874 424226 151494 424294
rect 150874 424170 150970 424226
rect 151026 424170 151094 424226
rect 151150 424170 151218 424226
rect 151274 424170 151342 424226
rect 151398 424170 151494 424226
rect 150874 424102 151494 424170
rect 150874 424046 150970 424102
rect 151026 424046 151094 424102
rect 151150 424046 151218 424102
rect 151274 424046 151342 424102
rect 151398 424046 151494 424102
rect 150874 423978 151494 424046
rect 150874 423922 150970 423978
rect 151026 423922 151094 423978
rect 151150 423922 151218 423978
rect 151274 423922 151342 423978
rect 151398 423922 151494 423978
rect 150874 406350 151494 423922
rect 150874 406294 150970 406350
rect 151026 406294 151094 406350
rect 151150 406294 151218 406350
rect 151274 406294 151342 406350
rect 151398 406294 151494 406350
rect 150874 406226 151494 406294
rect 150874 406170 150970 406226
rect 151026 406170 151094 406226
rect 151150 406170 151218 406226
rect 151274 406170 151342 406226
rect 151398 406170 151494 406226
rect 150874 406102 151494 406170
rect 150874 406046 150970 406102
rect 151026 406046 151094 406102
rect 151150 406046 151218 406102
rect 151274 406046 151342 406102
rect 151398 406046 151494 406102
rect 150874 405978 151494 406046
rect 150874 405922 150970 405978
rect 151026 405922 151094 405978
rect 151150 405922 151218 405978
rect 151274 405922 151342 405978
rect 151398 405922 151494 405978
rect 150874 388350 151494 405922
rect 150874 388294 150970 388350
rect 151026 388294 151094 388350
rect 151150 388294 151218 388350
rect 151274 388294 151342 388350
rect 151398 388294 151494 388350
rect 150874 388226 151494 388294
rect 150874 388170 150970 388226
rect 151026 388170 151094 388226
rect 151150 388170 151218 388226
rect 151274 388170 151342 388226
rect 151398 388170 151494 388226
rect 150874 388102 151494 388170
rect 150874 388046 150970 388102
rect 151026 388046 151094 388102
rect 151150 388046 151218 388102
rect 151274 388046 151342 388102
rect 151398 388046 151494 388102
rect 150874 387978 151494 388046
rect 150874 387922 150970 387978
rect 151026 387922 151094 387978
rect 151150 387922 151218 387978
rect 151274 387922 151342 387978
rect 151398 387922 151494 387978
rect 150874 370350 151494 387922
rect 150874 370294 150970 370350
rect 151026 370294 151094 370350
rect 151150 370294 151218 370350
rect 151274 370294 151342 370350
rect 151398 370294 151494 370350
rect 150874 370226 151494 370294
rect 150874 370170 150970 370226
rect 151026 370170 151094 370226
rect 151150 370170 151218 370226
rect 151274 370170 151342 370226
rect 151398 370170 151494 370226
rect 150874 370102 151494 370170
rect 150874 370046 150970 370102
rect 151026 370046 151094 370102
rect 151150 370046 151218 370102
rect 151274 370046 151342 370102
rect 151398 370046 151494 370102
rect 150874 369978 151494 370046
rect 150874 369922 150970 369978
rect 151026 369922 151094 369978
rect 151150 369922 151218 369978
rect 151274 369922 151342 369978
rect 151398 369922 151494 369978
rect 150874 352350 151494 369922
rect 150874 352294 150970 352350
rect 151026 352294 151094 352350
rect 151150 352294 151218 352350
rect 151274 352294 151342 352350
rect 151398 352294 151494 352350
rect 150874 352226 151494 352294
rect 150874 352170 150970 352226
rect 151026 352170 151094 352226
rect 151150 352170 151218 352226
rect 151274 352170 151342 352226
rect 151398 352170 151494 352226
rect 150874 352102 151494 352170
rect 150874 352046 150970 352102
rect 151026 352046 151094 352102
rect 151150 352046 151218 352102
rect 151274 352046 151342 352102
rect 151398 352046 151494 352102
rect 150874 351978 151494 352046
rect 150874 351922 150970 351978
rect 151026 351922 151094 351978
rect 151150 351922 151218 351978
rect 151274 351922 151342 351978
rect 151398 351922 151494 351978
rect 150874 334350 151494 351922
rect 150874 334294 150970 334350
rect 151026 334294 151094 334350
rect 151150 334294 151218 334350
rect 151274 334294 151342 334350
rect 151398 334294 151494 334350
rect 150874 334226 151494 334294
rect 150874 334170 150970 334226
rect 151026 334170 151094 334226
rect 151150 334170 151218 334226
rect 151274 334170 151342 334226
rect 151398 334170 151494 334226
rect 150874 334102 151494 334170
rect 150874 334046 150970 334102
rect 151026 334046 151094 334102
rect 151150 334046 151218 334102
rect 151274 334046 151342 334102
rect 151398 334046 151494 334102
rect 150874 333978 151494 334046
rect 150874 333922 150970 333978
rect 151026 333922 151094 333978
rect 151150 333922 151218 333978
rect 151274 333922 151342 333978
rect 151398 333922 151494 333978
rect 150874 316350 151494 333922
rect 150874 316294 150970 316350
rect 151026 316294 151094 316350
rect 151150 316294 151218 316350
rect 151274 316294 151342 316350
rect 151398 316294 151494 316350
rect 150874 316226 151494 316294
rect 150874 316170 150970 316226
rect 151026 316170 151094 316226
rect 151150 316170 151218 316226
rect 151274 316170 151342 316226
rect 151398 316170 151494 316226
rect 150874 316102 151494 316170
rect 150874 316046 150970 316102
rect 151026 316046 151094 316102
rect 151150 316046 151218 316102
rect 151274 316046 151342 316102
rect 151398 316046 151494 316102
rect 150874 315978 151494 316046
rect 150874 315922 150970 315978
rect 151026 315922 151094 315978
rect 151150 315922 151218 315978
rect 151274 315922 151342 315978
rect 151398 315922 151494 315978
rect 150874 298350 151494 315922
rect 150874 298294 150970 298350
rect 151026 298294 151094 298350
rect 151150 298294 151218 298350
rect 151274 298294 151342 298350
rect 151398 298294 151494 298350
rect 150874 298226 151494 298294
rect 150874 298170 150970 298226
rect 151026 298170 151094 298226
rect 151150 298170 151218 298226
rect 151274 298170 151342 298226
rect 151398 298170 151494 298226
rect 150874 298102 151494 298170
rect 150874 298046 150970 298102
rect 151026 298046 151094 298102
rect 151150 298046 151218 298102
rect 151274 298046 151342 298102
rect 151398 298046 151494 298102
rect 150874 297978 151494 298046
rect 150874 297922 150970 297978
rect 151026 297922 151094 297978
rect 151150 297922 151218 297978
rect 151274 297922 151342 297978
rect 151398 297922 151494 297978
rect 150874 280350 151494 297922
rect 150874 280294 150970 280350
rect 151026 280294 151094 280350
rect 151150 280294 151218 280350
rect 151274 280294 151342 280350
rect 151398 280294 151494 280350
rect 150874 280226 151494 280294
rect 150874 280170 150970 280226
rect 151026 280170 151094 280226
rect 151150 280170 151218 280226
rect 151274 280170 151342 280226
rect 151398 280170 151494 280226
rect 150874 280102 151494 280170
rect 150874 280046 150970 280102
rect 151026 280046 151094 280102
rect 151150 280046 151218 280102
rect 151274 280046 151342 280102
rect 151398 280046 151494 280102
rect 150874 279978 151494 280046
rect 150874 279922 150970 279978
rect 151026 279922 151094 279978
rect 151150 279922 151218 279978
rect 151274 279922 151342 279978
rect 151398 279922 151494 279978
rect 150874 262350 151494 279922
rect 150874 262294 150970 262350
rect 151026 262294 151094 262350
rect 151150 262294 151218 262350
rect 151274 262294 151342 262350
rect 151398 262294 151494 262350
rect 150874 262226 151494 262294
rect 150874 262170 150970 262226
rect 151026 262170 151094 262226
rect 151150 262170 151218 262226
rect 151274 262170 151342 262226
rect 151398 262170 151494 262226
rect 150874 262102 151494 262170
rect 150874 262046 150970 262102
rect 151026 262046 151094 262102
rect 151150 262046 151218 262102
rect 151274 262046 151342 262102
rect 151398 262046 151494 262102
rect 150874 261978 151494 262046
rect 150874 261922 150970 261978
rect 151026 261922 151094 261978
rect 151150 261922 151218 261978
rect 151274 261922 151342 261978
rect 151398 261922 151494 261978
rect 150874 244350 151494 261922
rect 150874 244294 150970 244350
rect 151026 244294 151094 244350
rect 151150 244294 151218 244350
rect 151274 244294 151342 244350
rect 151398 244294 151494 244350
rect 150874 244226 151494 244294
rect 150874 244170 150970 244226
rect 151026 244170 151094 244226
rect 151150 244170 151218 244226
rect 151274 244170 151342 244226
rect 151398 244170 151494 244226
rect 150874 244102 151494 244170
rect 150874 244046 150970 244102
rect 151026 244046 151094 244102
rect 151150 244046 151218 244102
rect 151274 244046 151342 244102
rect 151398 244046 151494 244102
rect 150874 243978 151494 244046
rect 150874 243922 150970 243978
rect 151026 243922 151094 243978
rect 151150 243922 151218 243978
rect 151274 243922 151342 243978
rect 151398 243922 151494 243978
rect 150874 226350 151494 243922
rect 168874 598172 169494 598268
rect 168874 598116 168970 598172
rect 169026 598116 169094 598172
rect 169150 598116 169218 598172
rect 169274 598116 169342 598172
rect 169398 598116 169494 598172
rect 168874 598048 169494 598116
rect 168874 597992 168970 598048
rect 169026 597992 169094 598048
rect 169150 597992 169218 598048
rect 169274 597992 169342 598048
rect 169398 597992 169494 598048
rect 168874 597924 169494 597992
rect 168874 597868 168970 597924
rect 169026 597868 169094 597924
rect 169150 597868 169218 597924
rect 169274 597868 169342 597924
rect 169398 597868 169494 597924
rect 168874 597800 169494 597868
rect 168874 597744 168970 597800
rect 169026 597744 169094 597800
rect 169150 597744 169218 597800
rect 169274 597744 169342 597800
rect 169398 597744 169494 597800
rect 168874 586350 169494 597744
rect 168874 586294 168970 586350
rect 169026 586294 169094 586350
rect 169150 586294 169218 586350
rect 169274 586294 169342 586350
rect 169398 586294 169494 586350
rect 168874 586226 169494 586294
rect 168874 586170 168970 586226
rect 169026 586170 169094 586226
rect 169150 586170 169218 586226
rect 169274 586170 169342 586226
rect 169398 586170 169494 586226
rect 168874 586102 169494 586170
rect 168874 586046 168970 586102
rect 169026 586046 169094 586102
rect 169150 586046 169218 586102
rect 169274 586046 169342 586102
rect 169398 586046 169494 586102
rect 168874 585978 169494 586046
rect 168874 585922 168970 585978
rect 169026 585922 169094 585978
rect 169150 585922 169218 585978
rect 169274 585922 169342 585978
rect 169398 585922 169494 585978
rect 168874 568350 169494 585922
rect 168874 568294 168970 568350
rect 169026 568294 169094 568350
rect 169150 568294 169218 568350
rect 169274 568294 169342 568350
rect 169398 568294 169494 568350
rect 168874 568226 169494 568294
rect 168874 568170 168970 568226
rect 169026 568170 169094 568226
rect 169150 568170 169218 568226
rect 169274 568170 169342 568226
rect 169398 568170 169494 568226
rect 168874 568102 169494 568170
rect 168874 568046 168970 568102
rect 169026 568046 169094 568102
rect 169150 568046 169218 568102
rect 169274 568046 169342 568102
rect 169398 568046 169494 568102
rect 168874 567978 169494 568046
rect 168874 567922 168970 567978
rect 169026 567922 169094 567978
rect 169150 567922 169218 567978
rect 169274 567922 169342 567978
rect 169398 567922 169494 567978
rect 168874 550350 169494 567922
rect 168874 550294 168970 550350
rect 169026 550294 169094 550350
rect 169150 550294 169218 550350
rect 169274 550294 169342 550350
rect 169398 550294 169494 550350
rect 168874 550226 169494 550294
rect 168874 550170 168970 550226
rect 169026 550170 169094 550226
rect 169150 550170 169218 550226
rect 169274 550170 169342 550226
rect 169398 550170 169494 550226
rect 168874 550102 169494 550170
rect 168874 550046 168970 550102
rect 169026 550046 169094 550102
rect 169150 550046 169218 550102
rect 169274 550046 169342 550102
rect 169398 550046 169494 550102
rect 168874 549978 169494 550046
rect 168874 549922 168970 549978
rect 169026 549922 169094 549978
rect 169150 549922 169218 549978
rect 169274 549922 169342 549978
rect 169398 549922 169494 549978
rect 168874 532350 169494 549922
rect 168874 532294 168970 532350
rect 169026 532294 169094 532350
rect 169150 532294 169218 532350
rect 169274 532294 169342 532350
rect 169398 532294 169494 532350
rect 168874 532226 169494 532294
rect 168874 532170 168970 532226
rect 169026 532170 169094 532226
rect 169150 532170 169218 532226
rect 169274 532170 169342 532226
rect 169398 532170 169494 532226
rect 168874 532102 169494 532170
rect 168874 532046 168970 532102
rect 169026 532046 169094 532102
rect 169150 532046 169218 532102
rect 169274 532046 169342 532102
rect 169398 532046 169494 532102
rect 168874 531978 169494 532046
rect 168874 531922 168970 531978
rect 169026 531922 169094 531978
rect 169150 531922 169218 531978
rect 169274 531922 169342 531978
rect 169398 531922 169494 531978
rect 168874 514350 169494 531922
rect 168874 514294 168970 514350
rect 169026 514294 169094 514350
rect 169150 514294 169218 514350
rect 169274 514294 169342 514350
rect 169398 514294 169494 514350
rect 168874 514226 169494 514294
rect 168874 514170 168970 514226
rect 169026 514170 169094 514226
rect 169150 514170 169218 514226
rect 169274 514170 169342 514226
rect 169398 514170 169494 514226
rect 168874 514102 169494 514170
rect 168874 514046 168970 514102
rect 169026 514046 169094 514102
rect 169150 514046 169218 514102
rect 169274 514046 169342 514102
rect 169398 514046 169494 514102
rect 168874 513978 169494 514046
rect 168874 513922 168970 513978
rect 169026 513922 169094 513978
rect 169150 513922 169218 513978
rect 169274 513922 169342 513978
rect 169398 513922 169494 513978
rect 168874 496350 169494 513922
rect 168874 496294 168970 496350
rect 169026 496294 169094 496350
rect 169150 496294 169218 496350
rect 169274 496294 169342 496350
rect 169398 496294 169494 496350
rect 168874 496226 169494 496294
rect 168874 496170 168970 496226
rect 169026 496170 169094 496226
rect 169150 496170 169218 496226
rect 169274 496170 169342 496226
rect 169398 496170 169494 496226
rect 168874 496102 169494 496170
rect 168874 496046 168970 496102
rect 169026 496046 169094 496102
rect 169150 496046 169218 496102
rect 169274 496046 169342 496102
rect 169398 496046 169494 496102
rect 168874 495978 169494 496046
rect 168874 495922 168970 495978
rect 169026 495922 169094 495978
rect 169150 495922 169218 495978
rect 169274 495922 169342 495978
rect 169398 495922 169494 495978
rect 168874 478350 169494 495922
rect 168874 478294 168970 478350
rect 169026 478294 169094 478350
rect 169150 478294 169218 478350
rect 169274 478294 169342 478350
rect 169398 478294 169494 478350
rect 168874 478226 169494 478294
rect 168874 478170 168970 478226
rect 169026 478170 169094 478226
rect 169150 478170 169218 478226
rect 169274 478170 169342 478226
rect 169398 478170 169494 478226
rect 168874 478102 169494 478170
rect 168874 478046 168970 478102
rect 169026 478046 169094 478102
rect 169150 478046 169218 478102
rect 169274 478046 169342 478102
rect 169398 478046 169494 478102
rect 168874 477978 169494 478046
rect 168874 477922 168970 477978
rect 169026 477922 169094 477978
rect 169150 477922 169218 477978
rect 169274 477922 169342 477978
rect 169398 477922 169494 477978
rect 168874 460350 169494 477922
rect 168874 460294 168970 460350
rect 169026 460294 169094 460350
rect 169150 460294 169218 460350
rect 169274 460294 169342 460350
rect 169398 460294 169494 460350
rect 168874 460226 169494 460294
rect 168874 460170 168970 460226
rect 169026 460170 169094 460226
rect 169150 460170 169218 460226
rect 169274 460170 169342 460226
rect 169398 460170 169494 460226
rect 168874 460102 169494 460170
rect 168874 460046 168970 460102
rect 169026 460046 169094 460102
rect 169150 460046 169218 460102
rect 169274 460046 169342 460102
rect 169398 460046 169494 460102
rect 168874 459978 169494 460046
rect 168874 459922 168970 459978
rect 169026 459922 169094 459978
rect 169150 459922 169218 459978
rect 169274 459922 169342 459978
rect 169398 459922 169494 459978
rect 168874 442350 169494 459922
rect 168874 442294 168970 442350
rect 169026 442294 169094 442350
rect 169150 442294 169218 442350
rect 169274 442294 169342 442350
rect 169398 442294 169494 442350
rect 168874 442226 169494 442294
rect 168874 442170 168970 442226
rect 169026 442170 169094 442226
rect 169150 442170 169218 442226
rect 169274 442170 169342 442226
rect 169398 442170 169494 442226
rect 168874 442102 169494 442170
rect 168874 442046 168970 442102
rect 169026 442046 169094 442102
rect 169150 442046 169218 442102
rect 169274 442046 169342 442102
rect 169398 442046 169494 442102
rect 168874 441978 169494 442046
rect 168874 441922 168970 441978
rect 169026 441922 169094 441978
rect 169150 441922 169218 441978
rect 169274 441922 169342 441978
rect 169398 441922 169494 441978
rect 168874 424350 169494 441922
rect 168874 424294 168970 424350
rect 169026 424294 169094 424350
rect 169150 424294 169218 424350
rect 169274 424294 169342 424350
rect 169398 424294 169494 424350
rect 168874 424226 169494 424294
rect 168874 424170 168970 424226
rect 169026 424170 169094 424226
rect 169150 424170 169218 424226
rect 169274 424170 169342 424226
rect 169398 424170 169494 424226
rect 168874 424102 169494 424170
rect 168874 424046 168970 424102
rect 169026 424046 169094 424102
rect 169150 424046 169218 424102
rect 169274 424046 169342 424102
rect 169398 424046 169494 424102
rect 168874 423978 169494 424046
rect 168874 423922 168970 423978
rect 169026 423922 169094 423978
rect 169150 423922 169218 423978
rect 169274 423922 169342 423978
rect 169398 423922 169494 423978
rect 168874 406350 169494 423922
rect 168874 406294 168970 406350
rect 169026 406294 169094 406350
rect 169150 406294 169218 406350
rect 169274 406294 169342 406350
rect 169398 406294 169494 406350
rect 168874 406226 169494 406294
rect 168874 406170 168970 406226
rect 169026 406170 169094 406226
rect 169150 406170 169218 406226
rect 169274 406170 169342 406226
rect 169398 406170 169494 406226
rect 168874 406102 169494 406170
rect 168874 406046 168970 406102
rect 169026 406046 169094 406102
rect 169150 406046 169218 406102
rect 169274 406046 169342 406102
rect 169398 406046 169494 406102
rect 168874 405978 169494 406046
rect 168874 405922 168970 405978
rect 169026 405922 169094 405978
rect 169150 405922 169218 405978
rect 169274 405922 169342 405978
rect 169398 405922 169494 405978
rect 168874 388350 169494 405922
rect 168874 388294 168970 388350
rect 169026 388294 169094 388350
rect 169150 388294 169218 388350
rect 169274 388294 169342 388350
rect 169398 388294 169494 388350
rect 168874 388226 169494 388294
rect 168874 388170 168970 388226
rect 169026 388170 169094 388226
rect 169150 388170 169218 388226
rect 169274 388170 169342 388226
rect 169398 388170 169494 388226
rect 168874 388102 169494 388170
rect 168874 388046 168970 388102
rect 169026 388046 169094 388102
rect 169150 388046 169218 388102
rect 169274 388046 169342 388102
rect 169398 388046 169494 388102
rect 168874 387978 169494 388046
rect 168874 387922 168970 387978
rect 169026 387922 169094 387978
rect 169150 387922 169218 387978
rect 169274 387922 169342 387978
rect 169398 387922 169494 387978
rect 168874 370350 169494 387922
rect 168874 370294 168970 370350
rect 169026 370294 169094 370350
rect 169150 370294 169218 370350
rect 169274 370294 169342 370350
rect 169398 370294 169494 370350
rect 168874 370226 169494 370294
rect 168874 370170 168970 370226
rect 169026 370170 169094 370226
rect 169150 370170 169218 370226
rect 169274 370170 169342 370226
rect 169398 370170 169494 370226
rect 168874 370102 169494 370170
rect 168874 370046 168970 370102
rect 169026 370046 169094 370102
rect 169150 370046 169218 370102
rect 169274 370046 169342 370102
rect 169398 370046 169494 370102
rect 168874 369978 169494 370046
rect 168874 369922 168970 369978
rect 169026 369922 169094 369978
rect 169150 369922 169218 369978
rect 169274 369922 169342 369978
rect 169398 369922 169494 369978
rect 168874 352350 169494 369922
rect 168874 352294 168970 352350
rect 169026 352294 169094 352350
rect 169150 352294 169218 352350
rect 169274 352294 169342 352350
rect 169398 352294 169494 352350
rect 168874 352226 169494 352294
rect 168874 352170 168970 352226
rect 169026 352170 169094 352226
rect 169150 352170 169218 352226
rect 169274 352170 169342 352226
rect 169398 352170 169494 352226
rect 168874 352102 169494 352170
rect 168874 352046 168970 352102
rect 169026 352046 169094 352102
rect 169150 352046 169218 352102
rect 169274 352046 169342 352102
rect 169398 352046 169494 352102
rect 168874 351978 169494 352046
rect 168874 351922 168970 351978
rect 169026 351922 169094 351978
rect 169150 351922 169218 351978
rect 169274 351922 169342 351978
rect 169398 351922 169494 351978
rect 168874 334350 169494 351922
rect 168874 334294 168970 334350
rect 169026 334294 169094 334350
rect 169150 334294 169218 334350
rect 169274 334294 169342 334350
rect 169398 334294 169494 334350
rect 168874 334226 169494 334294
rect 168874 334170 168970 334226
rect 169026 334170 169094 334226
rect 169150 334170 169218 334226
rect 169274 334170 169342 334226
rect 169398 334170 169494 334226
rect 168874 334102 169494 334170
rect 168874 334046 168970 334102
rect 169026 334046 169094 334102
rect 169150 334046 169218 334102
rect 169274 334046 169342 334102
rect 169398 334046 169494 334102
rect 168874 333978 169494 334046
rect 168874 333922 168970 333978
rect 169026 333922 169094 333978
rect 169150 333922 169218 333978
rect 169274 333922 169342 333978
rect 169398 333922 169494 333978
rect 168874 316350 169494 333922
rect 168874 316294 168970 316350
rect 169026 316294 169094 316350
rect 169150 316294 169218 316350
rect 169274 316294 169342 316350
rect 169398 316294 169494 316350
rect 168874 316226 169494 316294
rect 168874 316170 168970 316226
rect 169026 316170 169094 316226
rect 169150 316170 169218 316226
rect 169274 316170 169342 316226
rect 169398 316170 169494 316226
rect 168874 316102 169494 316170
rect 168874 316046 168970 316102
rect 169026 316046 169094 316102
rect 169150 316046 169218 316102
rect 169274 316046 169342 316102
rect 169398 316046 169494 316102
rect 168874 315978 169494 316046
rect 168874 315922 168970 315978
rect 169026 315922 169094 315978
rect 169150 315922 169218 315978
rect 169274 315922 169342 315978
rect 169398 315922 169494 315978
rect 168874 298350 169494 315922
rect 168874 298294 168970 298350
rect 169026 298294 169094 298350
rect 169150 298294 169218 298350
rect 169274 298294 169342 298350
rect 169398 298294 169494 298350
rect 168874 298226 169494 298294
rect 168874 298170 168970 298226
rect 169026 298170 169094 298226
rect 169150 298170 169218 298226
rect 169274 298170 169342 298226
rect 169398 298170 169494 298226
rect 168874 298102 169494 298170
rect 168874 298046 168970 298102
rect 169026 298046 169094 298102
rect 169150 298046 169218 298102
rect 169274 298046 169342 298102
rect 169398 298046 169494 298102
rect 168874 297978 169494 298046
rect 168874 297922 168970 297978
rect 169026 297922 169094 297978
rect 169150 297922 169218 297978
rect 169274 297922 169342 297978
rect 169398 297922 169494 297978
rect 168874 280350 169494 297922
rect 168874 280294 168970 280350
rect 169026 280294 169094 280350
rect 169150 280294 169218 280350
rect 169274 280294 169342 280350
rect 169398 280294 169494 280350
rect 168874 280226 169494 280294
rect 168874 280170 168970 280226
rect 169026 280170 169094 280226
rect 169150 280170 169218 280226
rect 169274 280170 169342 280226
rect 169398 280170 169494 280226
rect 168874 280102 169494 280170
rect 168874 280046 168970 280102
rect 169026 280046 169094 280102
rect 169150 280046 169218 280102
rect 169274 280046 169342 280102
rect 169398 280046 169494 280102
rect 168874 279978 169494 280046
rect 168874 279922 168970 279978
rect 169026 279922 169094 279978
rect 169150 279922 169218 279978
rect 169274 279922 169342 279978
rect 169398 279922 169494 279978
rect 168874 262350 169494 279922
rect 168874 262294 168970 262350
rect 169026 262294 169094 262350
rect 169150 262294 169218 262350
rect 169274 262294 169342 262350
rect 169398 262294 169494 262350
rect 168874 262226 169494 262294
rect 168874 262170 168970 262226
rect 169026 262170 169094 262226
rect 169150 262170 169218 262226
rect 169274 262170 169342 262226
rect 169398 262170 169494 262226
rect 168874 262102 169494 262170
rect 168874 262046 168970 262102
rect 169026 262046 169094 262102
rect 169150 262046 169218 262102
rect 169274 262046 169342 262102
rect 169398 262046 169494 262102
rect 168874 261978 169494 262046
rect 168874 261922 168970 261978
rect 169026 261922 169094 261978
rect 169150 261922 169218 261978
rect 169274 261922 169342 261978
rect 169398 261922 169494 261978
rect 168874 244350 169494 261922
rect 168874 244294 168970 244350
rect 169026 244294 169094 244350
rect 169150 244294 169218 244350
rect 169274 244294 169342 244350
rect 169398 244294 169494 244350
rect 168874 244226 169494 244294
rect 168874 244170 168970 244226
rect 169026 244170 169094 244226
rect 169150 244170 169218 244226
rect 169274 244170 169342 244226
rect 169398 244170 169494 244226
rect 168874 244102 169494 244170
rect 168874 244046 168970 244102
rect 169026 244046 169094 244102
rect 169150 244046 169218 244102
rect 169274 244046 169342 244102
rect 169398 244046 169494 244102
rect 168874 243978 169494 244046
rect 168874 243922 168970 243978
rect 169026 243922 169094 243978
rect 169150 243922 169218 243978
rect 169274 243922 169342 243978
rect 169398 243922 169494 243978
rect 150874 226294 150970 226350
rect 151026 226294 151094 226350
rect 151150 226294 151218 226350
rect 151274 226294 151342 226350
rect 151398 226294 151494 226350
rect 150874 226226 151494 226294
rect 150874 226170 150970 226226
rect 151026 226170 151094 226226
rect 151150 226170 151218 226226
rect 151274 226170 151342 226226
rect 151398 226170 151494 226226
rect 150874 226102 151494 226170
rect 150874 226046 150970 226102
rect 151026 226046 151094 226102
rect 151150 226046 151218 226102
rect 151274 226046 151342 226102
rect 151398 226046 151494 226102
rect 150874 225978 151494 226046
rect 150874 225922 150970 225978
rect 151026 225922 151094 225978
rect 151150 225922 151218 225978
rect 151274 225922 151342 225978
rect 151398 225922 151494 225978
rect 150874 219134 151494 225922
rect 165154 238350 165774 242964
rect 165154 238294 165250 238350
rect 165306 238294 165374 238350
rect 165430 238294 165498 238350
rect 165554 238294 165622 238350
rect 165678 238294 165774 238350
rect 165154 238226 165774 238294
rect 165154 238170 165250 238226
rect 165306 238170 165374 238226
rect 165430 238170 165498 238226
rect 165554 238170 165622 238226
rect 165678 238170 165774 238226
rect 165154 238102 165774 238170
rect 165154 238046 165250 238102
rect 165306 238046 165374 238102
rect 165430 238046 165498 238102
rect 165554 238046 165622 238102
rect 165678 238046 165774 238102
rect 165154 237978 165774 238046
rect 165154 237922 165250 237978
rect 165306 237922 165374 237978
rect 165430 237922 165498 237978
rect 165554 237922 165622 237978
rect 165678 237922 165774 237978
rect 156608 220350 156928 220384
rect 156608 220294 156678 220350
rect 156734 220294 156802 220350
rect 156858 220294 156928 220350
rect 156608 220226 156928 220294
rect 156608 220170 156678 220226
rect 156734 220170 156802 220226
rect 156858 220170 156928 220226
rect 156608 220102 156928 220170
rect 156608 220046 156678 220102
rect 156734 220046 156802 220102
rect 156858 220046 156928 220102
rect 156608 219978 156928 220046
rect 156608 219922 156678 219978
rect 156734 219922 156802 219978
rect 156858 219922 156928 219978
rect 156608 219888 156928 219922
rect 165154 220350 165774 237922
rect 165154 220294 165250 220350
rect 165306 220294 165374 220350
rect 165430 220294 165498 220350
rect 165554 220294 165622 220350
rect 165678 220294 165774 220350
rect 165154 220226 165774 220294
rect 165154 220170 165250 220226
rect 165306 220170 165374 220226
rect 165430 220170 165498 220226
rect 165554 220170 165622 220226
rect 165678 220170 165774 220226
rect 165154 220102 165774 220170
rect 165154 220046 165250 220102
rect 165306 220046 165374 220102
rect 165430 220046 165498 220102
rect 165554 220046 165622 220102
rect 165678 220046 165774 220102
rect 165154 219978 165774 220046
rect 165154 219922 165250 219978
rect 165306 219922 165374 219978
rect 165430 219922 165498 219978
rect 165554 219922 165622 219978
rect 165678 219922 165774 219978
rect 165154 219134 165774 219922
rect 168874 226350 169494 243922
rect 183154 597212 183774 598268
rect 183154 597156 183250 597212
rect 183306 597156 183374 597212
rect 183430 597156 183498 597212
rect 183554 597156 183622 597212
rect 183678 597156 183774 597212
rect 183154 597088 183774 597156
rect 183154 597032 183250 597088
rect 183306 597032 183374 597088
rect 183430 597032 183498 597088
rect 183554 597032 183622 597088
rect 183678 597032 183774 597088
rect 183154 596964 183774 597032
rect 183154 596908 183250 596964
rect 183306 596908 183374 596964
rect 183430 596908 183498 596964
rect 183554 596908 183622 596964
rect 183678 596908 183774 596964
rect 183154 596840 183774 596908
rect 183154 596784 183250 596840
rect 183306 596784 183374 596840
rect 183430 596784 183498 596840
rect 183554 596784 183622 596840
rect 183678 596784 183774 596840
rect 183154 580350 183774 596784
rect 183154 580294 183250 580350
rect 183306 580294 183374 580350
rect 183430 580294 183498 580350
rect 183554 580294 183622 580350
rect 183678 580294 183774 580350
rect 183154 580226 183774 580294
rect 183154 580170 183250 580226
rect 183306 580170 183374 580226
rect 183430 580170 183498 580226
rect 183554 580170 183622 580226
rect 183678 580170 183774 580226
rect 183154 580102 183774 580170
rect 183154 580046 183250 580102
rect 183306 580046 183374 580102
rect 183430 580046 183498 580102
rect 183554 580046 183622 580102
rect 183678 580046 183774 580102
rect 183154 579978 183774 580046
rect 183154 579922 183250 579978
rect 183306 579922 183374 579978
rect 183430 579922 183498 579978
rect 183554 579922 183622 579978
rect 183678 579922 183774 579978
rect 183154 562350 183774 579922
rect 183154 562294 183250 562350
rect 183306 562294 183374 562350
rect 183430 562294 183498 562350
rect 183554 562294 183622 562350
rect 183678 562294 183774 562350
rect 183154 562226 183774 562294
rect 183154 562170 183250 562226
rect 183306 562170 183374 562226
rect 183430 562170 183498 562226
rect 183554 562170 183622 562226
rect 183678 562170 183774 562226
rect 183154 562102 183774 562170
rect 183154 562046 183250 562102
rect 183306 562046 183374 562102
rect 183430 562046 183498 562102
rect 183554 562046 183622 562102
rect 183678 562046 183774 562102
rect 183154 561978 183774 562046
rect 183154 561922 183250 561978
rect 183306 561922 183374 561978
rect 183430 561922 183498 561978
rect 183554 561922 183622 561978
rect 183678 561922 183774 561978
rect 183154 544350 183774 561922
rect 183154 544294 183250 544350
rect 183306 544294 183374 544350
rect 183430 544294 183498 544350
rect 183554 544294 183622 544350
rect 183678 544294 183774 544350
rect 183154 544226 183774 544294
rect 183154 544170 183250 544226
rect 183306 544170 183374 544226
rect 183430 544170 183498 544226
rect 183554 544170 183622 544226
rect 183678 544170 183774 544226
rect 183154 544102 183774 544170
rect 183154 544046 183250 544102
rect 183306 544046 183374 544102
rect 183430 544046 183498 544102
rect 183554 544046 183622 544102
rect 183678 544046 183774 544102
rect 183154 543978 183774 544046
rect 183154 543922 183250 543978
rect 183306 543922 183374 543978
rect 183430 543922 183498 543978
rect 183554 543922 183622 543978
rect 183678 543922 183774 543978
rect 183154 526350 183774 543922
rect 183154 526294 183250 526350
rect 183306 526294 183374 526350
rect 183430 526294 183498 526350
rect 183554 526294 183622 526350
rect 183678 526294 183774 526350
rect 183154 526226 183774 526294
rect 183154 526170 183250 526226
rect 183306 526170 183374 526226
rect 183430 526170 183498 526226
rect 183554 526170 183622 526226
rect 183678 526170 183774 526226
rect 183154 526102 183774 526170
rect 183154 526046 183250 526102
rect 183306 526046 183374 526102
rect 183430 526046 183498 526102
rect 183554 526046 183622 526102
rect 183678 526046 183774 526102
rect 183154 525978 183774 526046
rect 183154 525922 183250 525978
rect 183306 525922 183374 525978
rect 183430 525922 183498 525978
rect 183554 525922 183622 525978
rect 183678 525922 183774 525978
rect 183154 508350 183774 525922
rect 183154 508294 183250 508350
rect 183306 508294 183374 508350
rect 183430 508294 183498 508350
rect 183554 508294 183622 508350
rect 183678 508294 183774 508350
rect 183154 508226 183774 508294
rect 183154 508170 183250 508226
rect 183306 508170 183374 508226
rect 183430 508170 183498 508226
rect 183554 508170 183622 508226
rect 183678 508170 183774 508226
rect 183154 508102 183774 508170
rect 183154 508046 183250 508102
rect 183306 508046 183374 508102
rect 183430 508046 183498 508102
rect 183554 508046 183622 508102
rect 183678 508046 183774 508102
rect 183154 507978 183774 508046
rect 183154 507922 183250 507978
rect 183306 507922 183374 507978
rect 183430 507922 183498 507978
rect 183554 507922 183622 507978
rect 183678 507922 183774 507978
rect 183154 490350 183774 507922
rect 183154 490294 183250 490350
rect 183306 490294 183374 490350
rect 183430 490294 183498 490350
rect 183554 490294 183622 490350
rect 183678 490294 183774 490350
rect 183154 490226 183774 490294
rect 183154 490170 183250 490226
rect 183306 490170 183374 490226
rect 183430 490170 183498 490226
rect 183554 490170 183622 490226
rect 183678 490170 183774 490226
rect 183154 490102 183774 490170
rect 183154 490046 183250 490102
rect 183306 490046 183374 490102
rect 183430 490046 183498 490102
rect 183554 490046 183622 490102
rect 183678 490046 183774 490102
rect 183154 489978 183774 490046
rect 183154 489922 183250 489978
rect 183306 489922 183374 489978
rect 183430 489922 183498 489978
rect 183554 489922 183622 489978
rect 183678 489922 183774 489978
rect 183154 472350 183774 489922
rect 183154 472294 183250 472350
rect 183306 472294 183374 472350
rect 183430 472294 183498 472350
rect 183554 472294 183622 472350
rect 183678 472294 183774 472350
rect 183154 472226 183774 472294
rect 183154 472170 183250 472226
rect 183306 472170 183374 472226
rect 183430 472170 183498 472226
rect 183554 472170 183622 472226
rect 183678 472170 183774 472226
rect 183154 472102 183774 472170
rect 183154 472046 183250 472102
rect 183306 472046 183374 472102
rect 183430 472046 183498 472102
rect 183554 472046 183622 472102
rect 183678 472046 183774 472102
rect 183154 471978 183774 472046
rect 183154 471922 183250 471978
rect 183306 471922 183374 471978
rect 183430 471922 183498 471978
rect 183554 471922 183622 471978
rect 183678 471922 183774 471978
rect 183154 454350 183774 471922
rect 183154 454294 183250 454350
rect 183306 454294 183374 454350
rect 183430 454294 183498 454350
rect 183554 454294 183622 454350
rect 183678 454294 183774 454350
rect 183154 454226 183774 454294
rect 183154 454170 183250 454226
rect 183306 454170 183374 454226
rect 183430 454170 183498 454226
rect 183554 454170 183622 454226
rect 183678 454170 183774 454226
rect 183154 454102 183774 454170
rect 183154 454046 183250 454102
rect 183306 454046 183374 454102
rect 183430 454046 183498 454102
rect 183554 454046 183622 454102
rect 183678 454046 183774 454102
rect 183154 453978 183774 454046
rect 183154 453922 183250 453978
rect 183306 453922 183374 453978
rect 183430 453922 183498 453978
rect 183554 453922 183622 453978
rect 183678 453922 183774 453978
rect 183154 436350 183774 453922
rect 183154 436294 183250 436350
rect 183306 436294 183374 436350
rect 183430 436294 183498 436350
rect 183554 436294 183622 436350
rect 183678 436294 183774 436350
rect 183154 436226 183774 436294
rect 183154 436170 183250 436226
rect 183306 436170 183374 436226
rect 183430 436170 183498 436226
rect 183554 436170 183622 436226
rect 183678 436170 183774 436226
rect 183154 436102 183774 436170
rect 183154 436046 183250 436102
rect 183306 436046 183374 436102
rect 183430 436046 183498 436102
rect 183554 436046 183622 436102
rect 183678 436046 183774 436102
rect 183154 435978 183774 436046
rect 183154 435922 183250 435978
rect 183306 435922 183374 435978
rect 183430 435922 183498 435978
rect 183554 435922 183622 435978
rect 183678 435922 183774 435978
rect 183154 418350 183774 435922
rect 183154 418294 183250 418350
rect 183306 418294 183374 418350
rect 183430 418294 183498 418350
rect 183554 418294 183622 418350
rect 183678 418294 183774 418350
rect 183154 418226 183774 418294
rect 183154 418170 183250 418226
rect 183306 418170 183374 418226
rect 183430 418170 183498 418226
rect 183554 418170 183622 418226
rect 183678 418170 183774 418226
rect 183154 418102 183774 418170
rect 183154 418046 183250 418102
rect 183306 418046 183374 418102
rect 183430 418046 183498 418102
rect 183554 418046 183622 418102
rect 183678 418046 183774 418102
rect 183154 417978 183774 418046
rect 183154 417922 183250 417978
rect 183306 417922 183374 417978
rect 183430 417922 183498 417978
rect 183554 417922 183622 417978
rect 183678 417922 183774 417978
rect 183154 400350 183774 417922
rect 183154 400294 183250 400350
rect 183306 400294 183374 400350
rect 183430 400294 183498 400350
rect 183554 400294 183622 400350
rect 183678 400294 183774 400350
rect 183154 400226 183774 400294
rect 183154 400170 183250 400226
rect 183306 400170 183374 400226
rect 183430 400170 183498 400226
rect 183554 400170 183622 400226
rect 183678 400170 183774 400226
rect 183154 400102 183774 400170
rect 183154 400046 183250 400102
rect 183306 400046 183374 400102
rect 183430 400046 183498 400102
rect 183554 400046 183622 400102
rect 183678 400046 183774 400102
rect 183154 399978 183774 400046
rect 183154 399922 183250 399978
rect 183306 399922 183374 399978
rect 183430 399922 183498 399978
rect 183554 399922 183622 399978
rect 183678 399922 183774 399978
rect 183154 382350 183774 399922
rect 183154 382294 183250 382350
rect 183306 382294 183374 382350
rect 183430 382294 183498 382350
rect 183554 382294 183622 382350
rect 183678 382294 183774 382350
rect 183154 382226 183774 382294
rect 183154 382170 183250 382226
rect 183306 382170 183374 382226
rect 183430 382170 183498 382226
rect 183554 382170 183622 382226
rect 183678 382170 183774 382226
rect 183154 382102 183774 382170
rect 183154 382046 183250 382102
rect 183306 382046 183374 382102
rect 183430 382046 183498 382102
rect 183554 382046 183622 382102
rect 183678 382046 183774 382102
rect 183154 381978 183774 382046
rect 183154 381922 183250 381978
rect 183306 381922 183374 381978
rect 183430 381922 183498 381978
rect 183554 381922 183622 381978
rect 183678 381922 183774 381978
rect 183154 364350 183774 381922
rect 183154 364294 183250 364350
rect 183306 364294 183374 364350
rect 183430 364294 183498 364350
rect 183554 364294 183622 364350
rect 183678 364294 183774 364350
rect 183154 364226 183774 364294
rect 183154 364170 183250 364226
rect 183306 364170 183374 364226
rect 183430 364170 183498 364226
rect 183554 364170 183622 364226
rect 183678 364170 183774 364226
rect 183154 364102 183774 364170
rect 183154 364046 183250 364102
rect 183306 364046 183374 364102
rect 183430 364046 183498 364102
rect 183554 364046 183622 364102
rect 183678 364046 183774 364102
rect 183154 363978 183774 364046
rect 183154 363922 183250 363978
rect 183306 363922 183374 363978
rect 183430 363922 183498 363978
rect 183554 363922 183622 363978
rect 183678 363922 183774 363978
rect 183154 346350 183774 363922
rect 183154 346294 183250 346350
rect 183306 346294 183374 346350
rect 183430 346294 183498 346350
rect 183554 346294 183622 346350
rect 183678 346294 183774 346350
rect 183154 346226 183774 346294
rect 183154 346170 183250 346226
rect 183306 346170 183374 346226
rect 183430 346170 183498 346226
rect 183554 346170 183622 346226
rect 183678 346170 183774 346226
rect 183154 346102 183774 346170
rect 183154 346046 183250 346102
rect 183306 346046 183374 346102
rect 183430 346046 183498 346102
rect 183554 346046 183622 346102
rect 183678 346046 183774 346102
rect 183154 345978 183774 346046
rect 183154 345922 183250 345978
rect 183306 345922 183374 345978
rect 183430 345922 183498 345978
rect 183554 345922 183622 345978
rect 183678 345922 183774 345978
rect 183154 328350 183774 345922
rect 183154 328294 183250 328350
rect 183306 328294 183374 328350
rect 183430 328294 183498 328350
rect 183554 328294 183622 328350
rect 183678 328294 183774 328350
rect 183154 328226 183774 328294
rect 183154 328170 183250 328226
rect 183306 328170 183374 328226
rect 183430 328170 183498 328226
rect 183554 328170 183622 328226
rect 183678 328170 183774 328226
rect 183154 328102 183774 328170
rect 183154 328046 183250 328102
rect 183306 328046 183374 328102
rect 183430 328046 183498 328102
rect 183554 328046 183622 328102
rect 183678 328046 183774 328102
rect 183154 327978 183774 328046
rect 183154 327922 183250 327978
rect 183306 327922 183374 327978
rect 183430 327922 183498 327978
rect 183554 327922 183622 327978
rect 183678 327922 183774 327978
rect 183154 310350 183774 327922
rect 183154 310294 183250 310350
rect 183306 310294 183374 310350
rect 183430 310294 183498 310350
rect 183554 310294 183622 310350
rect 183678 310294 183774 310350
rect 183154 310226 183774 310294
rect 183154 310170 183250 310226
rect 183306 310170 183374 310226
rect 183430 310170 183498 310226
rect 183554 310170 183622 310226
rect 183678 310170 183774 310226
rect 183154 310102 183774 310170
rect 183154 310046 183250 310102
rect 183306 310046 183374 310102
rect 183430 310046 183498 310102
rect 183554 310046 183622 310102
rect 183678 310046 183774 310102
rect 183154 309978 183774 310046
rect 183154 309922 183250 309978
rect 183306 309922 183374 309978
rect 183430 309922 183498 309978
rect 183554 309922 183622 309978
rect 183678 309922 183774 309978
rect 183154 292350 183774 309922
rect 183154 292294 183250 292350
rect 183306 292294 183374 292350
rect 183430 292294 183498 292350
rect 183554 292294 183622 292350
rect 183678 292294 183774 292350
rect 183154 292226 183774 292294
rect 183154 292170 183250 292226
rect 183306 292170 183374 292226
rect 183430 292170 183498 292226
rect 183554 292170 183622 292226
rect 183678 292170 183774 292226
rect 183154 292102 183774 292170
rect 183154 292046 183250 292102
rect 183306 292046 183374 292102
rect 183430 292046 183498 292102
rect 183554 292046 183622 292102
rect 183678 292046 183774 292102
rect 183154 291978 183774 292046
rect 183154 291922 183250 291978
rect 183306 291922 183374 291978
rect 183430 291922 183498 291978
rect 183554 291922 183622 291978
rect 183678 291922 183774 291978
rect 183154 274350 183774 291922
rect 183154 274294 183250 274350
rect 183306 274294 183374 274350
rect 183430 274294 183498 274350
rect 183554 274294 183622 274350
rect 183678 274294 183774 274350
rect 183154 274226 183774 274294
rect 183154 274170 183250 274226
rect 183306 274170 183374 274226
rect 183430 274170 183498 274226
rect 183554 274170 183622 274226
rect 183678 274170 183774 274226
rect 183154 274102 183774 274170
rect 183154 274046 183250 274102
rect 183306 274046 183374 274102
rect 183430 274046 183498 274102
rect 183554 274046 183622 274102
rect 183678 274046 183774 274102
rect 183154 273978 183774 274046
rect 183154 273922 183250 273978
rect 183306 273922 183374 273978
rect 183430 273922 183498 273978
rect 183554 273922 183622 273978
rect 183678 273922 183774 273978
rect 183154 256350 183774 273922
rect 183154 256294 183250 256350
rect 183306 256294 183374 256350
rect 183430 256294 183498 256350
rect 183554 256294 183622 256350
rect 183678 256294 183774 256350
rect 183154 256226 183774 256294
rect 183154 256170 183250 256226
rect 183306 256170 183374 256226
rect 183430 256170 183498 256226
rect 183554 256170 183622 256226
rect 183678 256170 183774 256226
rect 183154 256102 183774 256170
rect 183154 256046 183250 256102
rect 183306 256046 183374 256102
rect 183430 256046 183498 256102
rect 183554 256046 183622 256102
rect 183678 256046 183774 256102
rect 183154 255978 183774 256046
rect 183154 255922 183250 255978
rect 183306 255922 183374 255978
rect 183430 255922 183498 255978
rect 183554 255922 183622 255978
rect 183678 255922 183774 255978
rect 183154 238350 183774 255922
rect 183154 238294 183250 238350
rect 183306 238294 183374 238350
rect 183430 238294 183498 238350
rect 183554 238294 183622 238350
rect 183678 238294 183774 238350
rect 183154 238226 183774 238294
rect 183154 238170 183250 238226
rect 183306 238170 183374 238226
rect 183430 238170 183498 238226
rect 183554 238170 183622 238226
rect 183678 238170 183774 238226
rect 183154 238102 183774 238170
rect 183154 238046 183250 238102
rect 183306 238046 183374 238102
rect 183430 238046 183498 238102
rect 183554 238046 183622 238102
rect 183678 238046 183774 238102
rect 183154 237978 183774 238046
rect 183154 237922 183250 237978
rect 183306 237922 183374 237978
rect 183430 237922 183498 237978
rect 183554 237922 183622 237978
rect 183678 237922 183774 237978
rect 168874 226294 168970 226350
rect 169026 226294 169094 226350
rect 169150 226294 169218 226350
rect 169274 226294 169342 226350
rect 169398 226294 169494 226350
rect 168874 226226 169494 226294
rect 168874 226170 168970 226226
rect 169026 226170 169094 226226
rect 169150 226170 169218 226226
rect 169274 226170 169342 226226
rect 169398 226170 169494 226226
rect 168874 226102 169494 226170
rect 168874 226046 168970 226102
rect 169026 226046 169094 226102
rect 169150 226046 169218 226102
rect 169274 226046 169342 226102
rect 169398 226046 169494 226102
rect 168874 225978 169494 226046
rect 168874 225922 168970 225978
rect 169026 225922 169094 225978
rect 169150 225922 169218 225978
rect 169274 225922 169342 225978
rect 169398 225922 169494 225978
rect 168874 219134 169494 225922
rect 171968 226350 172288 226384
rect 171968 226294 172038 226350
rect 172094 226294 172162 226350
rect 172218 226294 172288 226350
rect 171968 226226 172288 226294
rect 171968 226170 172038 226226
rect 172094 226170 172162 226226
rect 172218 226170 172288 226226
rect 171968 226102 172288 226170
rect 171968 226046 172038 226102
rect 172094 226046 172162 226102
rect 172218 226046 172288 226102
rect 171968 225978 172288 226046
rect 171968 225922 172038 225978
rect 172094 225922 172162 225978
rect 172218 225922 172288 225978
rect 171968 225888 172288 225922
rect 183154 220350 183774 237922
rect 186874 598172 187494 598268
rect 186874 598116 186970 598172
rect 187026 598116 187094 598172
rect 187150 598116 187218 598172
rect 187274 598116 187342 598172
rect 187398 598116 187494 598172
rect 186874 598048 187494 598116
rect 186874 597992 186970 598048
rect 187026 597992 187094 598048
rect 187150 597992 187218 598048
rect 187274 597992 187342 598048
rect 187398 597992 187494 598048
rect 186874 597924 187494 597992
rect 186874 597868 186970 597924
rect 187026 597868 187094 597924
rect 187150 597868 187218 597924
rect 187274 597868 187342 597924
rect 187398 597868 187494 597924
rect 186874 597800 187494 597868
rect 186874 597744 186970 597800
rect 187026 597744 187094 597800
rect 187150 597744 187218 597800
rect 187274 597744 187342 597800
rect 187398 597744 187494 597800
rect 186874 586350 187494 597744
rect 186874 586294 186970 586350
rect 187026 586294 187094 586350
rect 187150 586294 187218 586350
rect 187274 586294 187342 586350
rect 187398 586294 187494 586350
rect 186874 586226 187494 586294
rect 186874 586170 186970 586226
rect 187026 586170 187094 586226
rect 187150 586170 187218 586226
rect 187274 586170 187342 586226
rect 187398 586170 187494 586226
rect 186874 586102 187494 586170
rect 186874 586046 186970 586102
rect 187026 586046 187094 586102
rect 187150 586046 187218 586102
rect 187274 586046 187342 586102
rect 187398 586046 187494 586102
rect 186874 585978 187494 586046
rect 186874 585922 186970 585978
rect 187026 585922 187094 585978
rect 187150 585922 187218 585978
rect 187274 585922 187342 585978
rect 187398 585922 187494 585978
rect 186874 568350 187494 585922
rect 186874 568294 186970 568350
rect 187026 568294 187094 568350
rect 187150 568294 187218 568350
rect 187274 568294 187342 568350
rect 187398 568294 187494 568350
rect 186874 568226 187494 568294
rect 186874 568170 186970 568226
rect 187026 568170 187094 568226
rect 187150 568170 187218 568226
rect 187274 568170 187342 568226
rect 187398 568170 187494 568226
rect 186874 568102 187494 568170
rect 186874 568046 186970 568102
rect 187026 568046 187094 568102
rect 187150 568046 187218 568102
rect 187274 568046 187342 568102
rect 187398 568046 187494 568102
rect 186874 567978 187494 568046
rect 186874 567922 186970 567978
rect 187026 567922 187094 567978
rect 187150 567922 187218 567978
rect 187274 567922 187342 567978
rect 187398 567922 187494 567978
rect 186874 550350 187494 567922
rect 186874 550294 186970 550350
rect 187026 550294 187094 550350
rect 187150 550294 187218 550350
rect 187274 550294 187342 550350
rect 187398 550294 187494 550350
rect 186874 550226 187494 550294
rect 186874 550170 186970 550226
rect 187026 550170 187094 550226
rect 187150 550170 187218 550226
rect 187274 550170 187342 550226
rect 187398 550170 187494 550226
rect 186874 550102 187494 550170
rect 186874 550046 186970 550102
rect 187026 550046 187094 550102
rect 187150 550046 187218 550102
rect 187274 550046 187342 550102
rect 187398 550046 187494 550102
rect 186874 549978 187494 550046
rect 186874 549922 186970 549978
rect 187026 549922 187094 549978
rect 187150 549922 187218 549978
rect 187274 549922 187342 549978
rect 187398 549922 187494 549978
rect 186874 532350 187494 549922
rect 186874 532294 186970 532350
rect 187026 532294 187094 532350
rect 187150 532294 187218 532350
rect 187274 532294 187342 532350
rect 187398 532294 187494 532350
rect 186874 532226 187494 532294
rect 186874 532170 186970 532226
rect 187026 532170 187094 532226
rect 187150 532170 187218 532226
rect 187274 532170 187342 532226
rect 187398 532170 187494 532226
rect 186874 532102 187494 532170
rect 186874 532046 186970 532102
rect 187026 532046 187094 532102
rect 187150 532046 187218 532102
rect 187274 532046 187342 532102
rect 187398 532046 187494 532102
rect 186874 531978 187494 532046
rect 186874 531922 186970 531978
rect 187026 531922 187094 531978
rect 187150 531922 187218 531978
rect 187274 531922 187342 531978
rect 187398 531922 187494 531978
rect 186874 514350 187494 531922
rect 186874 514294 186970 514350
rect 187026 514294 187094 514350
rect 187150 514294 187218 514350
rect 187274 514294 187342 514350
rect 187398 514294 187494 514350
rect 186874 514226 187494 514294
rect 186874 514170 186970 514226
rect 187026 514170 187094 514226
rect 187150 514170 187218 514226
rect 187274 514170 187342 514226
rect 187398 514170 187494 514226
rect 186874 514102 187494 514170
rect 186874 514046 186970 514102
rect 187026 514046 187094 514102
rect 187150 514046 187218 514102
rect 187274 514046 187342 514102
rect 187398 514046 187494 514102
rect 186874 513978 187494 514046
rect 186874 513922 186970 513978
rect 187026 513922 187094 513978
rect 187150 513922 187218 513978
rect 187274 513922 187342 513978
rect 187398 513922 187494 513978
rect 186874 496350 187494 513922
rect 186874 496294 186970 496350
rect 187026 496294 187094 496350
rect 187150 496294 187218 496350
rect 187274 496294 187342 496350
rect 187398 496294 187494 496350
rect 186874 496226 187494 496294
rect 186874 496170 186970 496226
rect 187026 496170 187094 496226
rect 187150 496170 187218 496226
rect 187274 496170 187342 496226
rect 187398 496170 187494 496226
rect 186874 496102 187494 496170
rect 186874 496046 186970 496102
rect 187026 496046 187094 496102
rect 187150 496046 187218 496102
rect 187274 496046 187342 496102
rect 187398 496046 187494 496102
rect 186874 495978 187494 496046
rect 186874 495922 186970 495978
rect 187026 495922 187094 495978
rect 187150 495922 187218 495978
rect 187274 495922 187342 495978
rect 187398 495922 187494 495978
rect 186874 478350 187494 495922
rect 186874 478294 186970 478350
rect 187026 478294 187094 478350
rect 187150 478294 187218 478350
rect 187274 478294 187342 478350
rect 187398 478294 187494 478350
rect 186874 478226 187494 478294
rect 186874 478170 186970 478226
rect 187026 478170 187094 478226
rect 187150 478170 187218 478226
rect 187274 478170 187342 478226
rect 187398 478170 187494 478226
rect 186874 478102 187494 478170
rect 186874 478046 186970 478102
rect 187026 478046 187094 478102
rect 187150 478046 187218 478102
rect 187274 478046 187342 478102
rect 187398 478046 187494 478102
rect 186874 477978 187494 478046
rect 186874 477922 186970 477978
rect 187026 477922 187094 477978
rect 187150 477922 187218 477978
rect 187274 477922 187342 477978
rect 187398 477922 187494 477978
rect 186874 460350 187494 477922
rect 186874 460294 186970 460350
rect 187026 460294 187094 460350
rect 187150 460294 187218 460350
rect 187274 460294 187342 460350
rect 187398 460294 187494 460350
rect 186874 460226 187494 460294
rect 186874 460170 186970 460226
rect 187026 460170 187094 460226
rect 187150 460170 187218 460226
rect 187274 460170 187342 460226
rect 187398 460170 187494 460226
rect 186874 460102 187494 460170
rect 186874 460046 186970 460102
rect 187026 460046 187094 460102
rect 187150 460046 187218 460102
rect 187274 460046 187342 460102
rect 187398 460046 187494 460102
rect 186874 459978 187494 460046
rect 186874 459922 186970 459978
rect 187026 459922 187094 459978
rect 187150 459922 187218 459978
rect 187274 459922 187342 459978
rect 187398 459922 187494 459978
rect 186874 442350 187494 459922
rect 186874 442294 186970 442350
rect 187026 442294 187094 442350
rect 187150 442294 187218 442350
rect 187274 442294 187342 442350
rect 187398 442294 187494 442350
rect 186874 442226 187494 442294
rect 186874 442170 186970 442226
rect 187026 442170 187094 442226
rect 187150 442170 187218 442226
rect 187274 442170 187342 442226
rect 187398 442170 187494 442226
rect 186874 442102 187494 442170
rect 186874 442046 186970 442102
rect 187026 442046 187094 442102
rect 187150 442046 187218 442102
rect 187274 442046 187342 442102
rect 187398 442046 187494 442102
rect 186874 441978 187494 442046
rect 186874 441922 186970 441978
rect 187026 441922 187094 441978
rect 187150 441922 187218 441978
rect 187274 441922 187342 441978
rect 187398 441922 187494 441978
rect 186874 424350 187494 441922
rect 186874 424294 186970 424350
rect 187026 424294 187094 424350
rect 187150 424294 187218 424350
rect 187274 424294 187342 424350
rect 187398 424294 187494 424350
rect 186874 424226 187494 424294
rect 186874 424170 186970 424226
rect 187026 424170 187094 424226
rect 187150 424170 187218 424226
rect 187274 424170 187342 424226
rect 187398 424170 187494 424226
rect 186874 424102 187494 424170
rect 186874 424046 186970 424102
rect 187026 424046 187094 424102
rect 187150 424046 187218 424102
rect 187274 424046 187342 424102
rect 187398 424046 187494 424102
rect 186874 423978 187494 424046
rect 186874 423922 186970 423978
rect 187026 423922 187094 423978
rect 187150 423922 187218 423978
rect 187274 423922 187342 423978
rect 187398 423922 187494 423978
rect 186874 406350 187494 423922
rect 186874 406294 186970 406350
rect 187026 406294 187094 406350
rect 187150 406294 187218 406350
rect 187274 406294 187342 406350
rect 187398 406294 187494 406350
rect 186874 406226 187494 406294
rect 186874 406170 186970 406226
rect 187026 406170 187094 406226
rect 187150 406170 187218 406226
rect 187274 406170 187342 406226
rect 187398 406170 187494 406226
rect 186874 406102 187494 406170
rect 186874 406046 186970 406102
rect 187026 406046 187094 406102
rect 187150 406046 187218 406102
rect 187274 406046 187342 406102
rect 187398 406046 187494 406102
rect 186874 405978 187494 406046
rect 186874 405922 186970 405978
rect 187026 405922 187094 405978
rect 187150 405922 187218 405978
rect 187274 405922 187342 405978
rect 187398 405922 187494 405978
rect 186874 388350 187494 405922
rect 186874 388294 186970 388350
rect 187026 388294 187094 388350
rect 187150 388294 187218 388350
rect 187274 388294 187342 388350
rect 187398 388294 187494 388350
rect 186874 388226 187494 388294
rect 186874 388170 186970 388226
rect 187026 388170 187094 388226
rect 187150 388170 187218 388226
rect 187274 388170 187342 388226
rect 187398 388170 187494 388226
rect 186874 388102 187494 388170
rect 186874 388046 186970 388102
rect 187026 388046 187094 388102
rect 187150 388046 187218 388102
rect 187274 388046 187342 388102
rect 187398 388046 187494 388102
rect 186874 387978 187494 388046
rect 186874 387922 186970 387978
rect 187026 387922 187094 387978
rect 187150 387922 187218 387978
rect 187274 387922 187342 387978
rect 187398 387922 187494 387978
rect 186874 370350 187494 387922
rect 186874 370294 186970 370350
rect 187026 370294 187094 370350
rect 187150 370294 187218 370350
rect 187274 370294 187342 370350
rect 187398 370294 187494 370350
rect 186874 370226 187494 370294
rect 186874 370170 186970 370226
rect 187026 370170 187094 370226
rect 187150 370170 187218 370226
rect 187274 370170 187342 370226
rect 187398 370170 187494 370226
rect 186874 370102 187494 370170
rect 186874 370046 186970 370102
rect 187026 370046 187094 370102
rect 187150 370046 187218 370102
rect 187274 370046 187342 370102
rect 187398 370046 187494 370102
rect 186874 369978 187494 370046
rect 186874 369922 186970 369978
rect 187026 369922 187094 369978
rect 187150 369922 187218 369978
rect 187274 369922 187342 369978
rect 187398 369922 187494 369978
rect 186874 352350 187494 369922
rect 186874 352294 186970 352350
rect 187026 352294 187094 352350
rect 187150 352294 187218 352350
rect 187274 352294 187342 352350
rect 187398 352294 187494 352350
rect 186874 352226 187494 352294
rect 186874 352170 186970 352226
rect 187026 352170 187094 352226
rect 187150 352170 187218 352226
rect 187274 352170 187342 352226
rect 187398 352170 187494 352226
rect 186874 352102 187494 352170
rect 186874 352046 186970 352102
rect 187026 352046 187094 352102
rect 187150 352046 187218 352102
rect 187274 352046 187342 352102
rect 187398 352046 187494 352102
rect 186874 351978 187494 352046
rect 186874 351922 186970 351978
rect 187026 351922 187094 351978
rect 187150 351922 187218 351978
rect 187274 351922 187342 351978
rect 187398 351922 187494 351978
rect 186874 334350 187494 351922
rect 186874 334294 186970 334350
rect 187026 334294 187094 334350
rect 187150 334294 187218 334350
rect 187274 334294 187342 334350
rect 187398 334294 187494 334350
rect 186874 334226 187494 334294
rect 186874 334170 186970 334226
rect 187026 334170 187094 334226
rect 187150 334170 187218 334226
rect 187274 334170 187342 334226
rect 187398 334170 187494 334226
rect 186874 334102 187494 334170
rect 186874 334046 186970 334102
rect 187026 334046 187094 334102
rect 187150 334046 187218 334102
rect 187274 334046 187342 334102
rect 187398 334046 187494 334102
rect 186874 333978 187494 334046
rect 186874 333922 186970 333978
rect 187026 333922 187094 333978
rect 187150 333922 187218 333978
rect 187274 333922 187342 333978
rect 187398 333922 187494 333978
rect 186874 316350 187494 333922
rect 186874 316294 186970 316350
rect 187026 316294 187094 316350
rect 187150 316294 187218 316350
rect 187274 316294 187342 316350
rect 187398 316294 187494 316350
rect 186874 316226 187494 316294
rect 186874 316170 186970 316226
rect 187026 316170 187094 316226
rect 187150 316170 187218 316226
rect 187274 316170 187342 316226
rect 187398 316170 187494 316226
rect 186874 316102 187494 316170
rect 186874 316046 186970 316102
rect 187026 316046 187094 316102
rect 187150 316046 187218 316102
rect 187274 316046 187342 316102
rect 187398 316046 187494 316102
rect 186874 315978 187494 316046
rect 186874 315922 186970 315978
rect 187026 315922 187094 315978
rect 187150 315922 187218 315978
rect 187274 315922 187342 315978
rect 187398 315922 187494 315978
rect 186874 298350 187494 315922
rect 186874 298294 186970 298350
rect 187026 298294 187094 298350
rect 187150 298294 187218 298350
rect 187274 298294 187342 298350
rect 187398 298294 187494 298350
rect 186874 298226 187494 298294
rect 186874 298170 186970 298226
rect 187026 298170 187094 298226
rect 187150 298170 187218 298226
rect 187274 298170 187342 298226
rect 187398 298170 187494 298226
rect 186874 298102 187494 298170
rect 186874 298046 186970 298102
rect 187026 298046 187094 298102
rect 187150 298046 187218 298102
rect 187274 298046 187342 298102
rect 187398 298046 187494 298102
rect 186874 297978 187494 298046
rect 186874 297922 186970 297978
rect 187026 297922 187094 297978
rect 187150 297922 187218 297978
rect 187274 297922 187342 297978
rect 187398 297922 187494 297978
rect 186874 280350 187494 297922
rect 186874 280294 186970 280350
rect 187026 280294 187094 280350
rect 187150 280294 187218 280350
rect 187274 280294 187342 280350
rect 187398 280294 187494 280350
rect 186874 280226 187494 280294
rect 186874 280170 186970 280226
rect 187026 280170 187094 280226
rect 187150 280170 187218 280226
rect 187274 280170 187342 280226
rect 187398 280170 187494 280226
rect 186874 280102 187494 280170
rect 186874 280046 186970 280102
rect 187026 280046 187094 280102
rect 187150 280046 187218 280102
rect 187274 280046 187342 280102
rect 187398 280046 187494 280102
rect 186874 279978 187494 280046
rect 186874 279922 186970 279978
rect 187026 279922 187094 279978
rect 187150 279922 187218 279978
rect 187274 279922 187342 279978
rect 187398 279922 187494 279978
rect 186874 262350 187494 279922
rect 186874 262294 186970 262350
rect 187026 262294 187094 262350
rect 187150 262294 187218 262350
rect 187274 262294 187342 262350
rect 187398 262294 187494 262350
rect 186874 262226 187494 262294
rect 186874 262170 186970 262226
rect 187026 262170 187094 262226
rect 187150 262170 187218 262226
rect 187274 262170 187342 262226
rect 187398 262170 187494 262226
rect 186874 262102 187494 262170
rect 186874 262046 186970 262102
rect 187026 262046 187094 262102
rect 187150 262046 187218 262102
rect 187274 262046 187342 262102
rect 187398 262046 187494 262102
rect 186874 261978 187494 262046
rect 186874 261922 186970 261978
rect 187026 261922 187094 261978
rect 187150 261922 187218 261978
rect 187274 261922 187342 261978
rect 187398 261922 187494 261978
rect 186874 244350 187494 261922
rect 186874 244294 186970 244350
rect 187026 244294 187094 244350
rect 187150 244294 187218 244350
rect 187274 244294 187342 244350
rect 187398 244294 187494 244350
rect 186874 244226 187494 244294
rect 186874 244170 186970 244226
rect 187026 244170 187094 244226
rect 187150 244170 187218 244226
rect 187274 244170 187342 244226
rect 187398 244170 187494 244226
rect 186874 244102 187494 244170
rect 186874 244046 186970 244102
rect 187026 244046 187094 244102
rect 187150 244046 187218 244102
rect 187274 244046 187342 244102
rect 187398 244046 187494 244102
rect 186874 243978 187494 244046
rect 186874 243922 186970 243978
rect 187026 243922 187094 243978
rect 187150 243922 187218 243978
rect 187274 243922 187342 243978
rect 187398 243922 187494 243978
rect 186874 228956 187494 243922
rect 201154 597212 201774 598268
rect 201154 597156 201250 597212
rect 201306 597156 201374 597212
rect 201430 597156 201498 597212
rect 201554 597156 201622 597212
rect 201678 597156 201774 597212
rect 201154 597088 201774 597156
rect 201154 597032 201250 597088
rect 201306 597032 201374 597088
rect 201430 597032 201498 597088
rect 201554 597032 201622 597088
rect 201678 597032 201774 597088
rect 201154 596964 201774 597032
rect 201154 596908 201250 596964
rect 201306 596908 201374 596964
rect 201430 596908 201498 596964
rect 201554 596908 201622 596964
rect 201678 596908 201774 596964
rect 201154 596840 201774 596908
rect 201154 596784 201250 596840
rect 201306 596784 201374 596840
rect 201430 596784 201498 596840
rect 201554 596784 201622 596840
rect 201678 596784 201774 596840
rect 201154 580350 201774 596784
rect 201154 580294 201250 580350
rect 201306 580294 201374 580350
rect 201430 580294 201498 580350
rect 201554 580294 201622 580350
rect 201678 580294 201774 580350
rect 201154 580226 201774 580294
rect 201154 580170 201250 580226
rect 201306 580170 201374 580226
rect 201430 580170 201498 580226
rect 201554 580170 201622 580226
rect 201678 580170 201774 580226
rect 201154 580102 201774 580170
rect 201154 580046 201250 580102
rect 201306 580046 201374 580102
rect 201430 580046 201498 580102
rect 201554 580046 201622 580102
rect 201678 580046 201774 580102
rect 201154 579978 201774 580046
rect 201154 579922 201250 579978
rect 201306 579922 201374 579978
rect 201430 579922 201498 579978
rect 201554 579922 201622 579978
rect 201678 579922 201774 579978
rect 201154 562350 201774 579922
rect 201154 562294 201250 562350
rect 201306 562294 201374 562350
rect 201430 562294 201498 562350
rect 201554 562294 201622 562350
rect 201678 562294 201774 562350
rect 201154 562226 201774 562294
rect 201154 562170 201250 562226
rect 201306 562170 201374 562226
rect 201430 562170 201498 562226
rect 201554 562170 201622 562226
rect 201678 562170 201774 562226
rect 201154 562102 201774 562170
rect 201154 562046 201250 562102
rect 201306 562046 201374 562102
rect 201430 562046 201498 562102
rect 201554 562046 201622 562102
rect 201678 562046 201774 562102
rect 201154 561978 201774 562046
rect 201154 561922 201250 561978
rect 201306 561922 201374 561978
rect 201430 561922 201498 561978
rect 201554 561922 201622 561978
rect 201678 561922 201774 561978
rect 201154 544350 201774 561922
rect 201154 544294 201250 544350
rect 201306 544294 201374 544350
rect 201430 544294 201498 544350
rect 201554 544294 201622 544350
rect 201678 544294 201774 544350
rect 201154 544226 201774 544294
rect 201154 544170 201250 544226
rect 201306 544170 201374 544226
rect 201430 544170 201498 544226
rect 201554 544170 201622 544226
rect 201678 544170 201774 544226
rect 201154 544102 201774 544170
rect 201154 544046 201250 544102
rect 201306 544046 201374 544102
rect 201430 544046 201498 544102
rect 201554 544046 201622 544102
rect 201678 544046 201774 544102
rect 201154 543978 201774 544046
rect 201154 543922 201250 543978
rect 201306 543922 201374 543978
rect 201430 543922 201498 543978
rect 201554 543922 201622 543978
rect 201678 543922 201774 543978
rect 201154 526350 201774 543922
rect 201154 526294 201250 526350
rect 201306 526294 201374 526350
rect 201430 526294 201498 526350
rect 201554 526294 201622 526350
rect 201678 526294 201774 526350
rect 201154 526226 201774 526294
rect 201154 526170 201250 526226
rect 201306 526170 201374 526226
rect 201430 526170 201498 526226
rect 201554 526170 201622 526226
rect 201678 526170 201774 526226
rect 201154 526102 201774 526170
rect 201154 526046 201250 526102
rect 201306 526046 201374 526102
rect 201430 526046 201498 526102
rect 201554 526046 201622 526102
rect 201678 526046 201774 526102
rect 201154 525978 201774 526046
rect 201154 525922 201250 525978
rect 201306 525922 201374 525978
rect 201430 525922 201498 525978
rect 201554 525922 201622 525978
rect 201678 525922 201774 525978
rect 201154 508350 201774 525922
rect 201154 508294 201250 508350
rect 201306 508294 201374 508350
rect 201430 508294 201498 508350
rect 201554 508294 201622 508350
rect 201678 508294 201774 508350
rect 201154 508226 201774 508294
rect 201154 508170 201250 508226
rect 201306 508170 201374 508226
rect 201430 508170 201498 508226
rect 201554 508170 201622 508226
rect 201678 508170 201774 508226
rect 201154 508102 201774 508170
rect 201154 508046 201250 508102
rect 201306 508046 201374 508102
rect 201430 508046 201498 508102
rect 201554 508046 201622 508102
rect 201678 508046 201774 508102
rect 201154 507978 201774 508046
rect 201154 507922 201250 507978
rect 201306 507922 201374 507978
rect 201430 507922 201498 507978
rect 201554 507922 201622 507978
rect 201678 507922 201774 507978
rect 201154 490350 201774 507922
rect 201154 490294 201250 490350
rect 201306 490294 201374 490350
rect 201430 490294 201498 490350
rect 201554 490294 201622 490350
rect 201678 490294 201774 490350
rect 201154 490226 201774 490294
rect 201154 490170 201250 490226
rect 201306 490170 201374 490226
rect 201430 490170 201498 490226
rect 201554 490170 201622 490226
rect 201678 490170 201774 490226
rect 201154 490102 201774 490170
rect 201154 490046 201250 490102
rect 201306 490046 201374 490102
rect 201430 490046 201498 490102
rect 201554 490046 201622 490102
rect 201678 490046 201774 490102
rect 201154 489978 201774 490046
rect 201154 489922 201250 489978
rect 201306 489922 201374 489978
rect 201430 489922 201498 489978
rect 201554 489922 201622 489978
rect 201678 489922 201774 489978
rect 201154 472350 201774 489922
rect 201154 472294 201250 472350
rect 201306 472294 201374 472350
rect 201430 472294 201498 472350
rect 201554 472294 201622 472350
rect 201678 472294 201774 472350
rect 201154 472226 201774 472294
rect 201154 472170 201250 472226
rect 201306 472170 201374 472226
rect 201430 472170 201498 472226
rect 201554 472170 201622 472226
rect 201678 472170 201774 472226
rect 201154 472102 201774 472170
rect 201154 472046 201250 472102
rect 201306 472046 201374 472102
rect 201430 472046 201498 472102
rect 201554 472046 201622 472102
rect 201678 472046 201774 472102
rect 201154 471978 201774 472046
rect 201154 471922 201250 471978
rect 201306 471922 201374 471978
rect 201430 471922 201498 471978
rect 201554 471922 201622 471978
rect 201678 471922 201774 471978
rect 201154 454350 201774 471922
rect 201154 454294 201250 454350
rect 201306 454294 201374 454350
rect 201430 454294 201498 454350
rect 201554 454294 201622 454350
rect 201678 454294 201774 454350
rect 201154 454226 201774 454294
rect 201154 454170 201250 454226
rect 201306 454170 201374 454226
rect 201430 454170 201498 454226
rect 201554 454170 201622 454226
rect 201678 454170 201774 454226
rect 201154 454102 201774 454170
rect 201154 454046 201250 454102
rect 201306 454046 201374 454102
rect 201430 454046 201498 454102
rect 201554 454046 201622 454102
rect 201678 454046 201774 454102
rect 201154 453978 201774 454046
rect 201154 453922 201250 453978
rect 201306 453922 201374 453978
rect 201430 453922 201498 453978
rect 201554 453922 201622 453978
rect 201678 453922 201774 453978
rect 201154 436350 201774 453922
rect 201154 436294 201250 436350
rect 201306 436294 201374 436350
rect 201430 436294 201498 436350
rect 201554 436294 201622 436350
rect 201678 436294 201774 436350
rect 201154 436226 201774 436294
rect 201154 436170 201250 436226
rect 201306 436170 201374 436226
rect 201430 436170 201498 436226
rect 201554 436170 201622 436226
rect 201678 436170 201774 436226
rect 201154 436102 201774 436170
rect 201154 436046 201250 436102
rect 201306 436046 201374 436102
rect 201430 436046 201498 436102
rect 201554 436046 201622 436102
rect 201678 436046 201774 436102
rect 201154 435978 201774 436046
rect 201154 435922 201250 435978
rect 201306 435922 201374 435978
rect 201430 435922 201498 435978
rect 201554 435922 201622 435978
rect 201678 435922 201774 435978
rect 201154 418350 201774 435922
rect 201154 418294 201250 418350
rect 201306 418294 201374 418350
rect 201430 418294 201498 418350
rect 201554 418294 201622 418350
rect 201678 418294 201774 418350
rect 201154 418226 201774 418294
rect 201154 418170 201250 418226
rect 201306 418170 201374 418226
rect 201430 418170 201498 418226
rect 201554 418170 201622 418226
rect 201678 418170 201774 418226
rect 201154 418102 201774 418170
rect 201154 418046 201250 418102
rect 201306 418046 201374 418102
rect 201430 418046 201498 418102
rect 201554 418046 201622 418102
rect 201678 418046 201774 418102
rect 201154 417978 201774 418046
rect 201154 417922 201250 417978
rect 201306 417922 201374 417978
rect 201430 417922 201498 417978
rect 201554 417922 201622 417978
rect 201678 417922 201774 417978
rect 201154 400350 201774 417922
rect 201154 400294 201250 400350
rect 201306 400294 201374 400350
rect 201430 400294 201498 400350
rect 201554 400294 201622 400350
rect 201678 400294 201774 400350
rect 201154 400226 201774 400294
rect 201154 400170 201250 400226
rect 201306 400170 201374 400226
rect 201430 400170 201498 400226
rect 201554 400170 201622 400226
rect 201678 400170 201774 400226
rect 201154 400102 201774 400170
rect 201154 400046 201250 400102
rect 201306 400046 201374 400102
rect 201430 400046 201498 400102
rect 201554 400046 201622 400102
rect 201678 400046 201774 400102
rect 201154 399978 201774 400046
rect 201154 399922 201250 399978
rect 201306 399922 201374 399978
rect 201430 399922 201498 399978
rect 201554 399922 201622 399978
rect 201678 399922 201774 399978
rect 201154 382350 201774 399922
rect 201154 382294 201250 382350
rect 201306 382294 201374 382350
rect 201430 382294 201498 382350
rect 201554 382294 201622 382350
rect 201678 382294 201774 382350
rect 201154 382226 201774 382294
rect 201154 382170 201250 382226
rect 201306 382170 201374 382226
rect 201430 382170 201498 382226
rect 201554 382170 201622 382226
rect 201678 382170 201774 382226
rect 201154 382102 201774 382170
rect 201154 382046 201250 382102
rect 201306 382046 201374 382102
rect 201430 382046 201498 382102
rect 201554 382046 201622 382102
rect 201678 382046 201774 382102
rect 201154 381978 201774 382046
rect 201154 381922 201250 381978
rect 201306 381922 201374 381978
rect 201430 381922 201498 381978
rect 201554 381922 201622 381978
rect 201678 381922 201774 381978
rect 201154 364350 201774 381922
rect 201154 364294 201250 364350
rect 201306 364294 201374 364350
rect 201430 364294 201498 364350
rect 201554 364294 201622 364350
rect 201678 364294 201774 364350
rect 201154 364226 201774 364294
rect 201154 364170 201250 364226
rect 201306 364170 201374 364226
rect 201430 364170 201498 364226
rect 201554 364170 201622 364226
rect 201678 364170 201774 364226
rect 201154 364102 201774 364170
rect 201154 364046 201250 364102
rect 201306 364046 201374 364102
rect 201430 364046 201498 364102
rect 201554 364046 201622 364102
rect 201678 364046 201774 364102
rect 201154 363978 201774 364046
rect 201154 363922 201250 363978
rect 201306 363922 201374 363978
rect 201430 363922 201498 363978
rect 201554 363922 201622 363978
rect 201678 363922 201774 363978
rect 201154 346350 201774 363922
rect 201154 346294 201250 346350
rect 201306 346294 201374 346350
rect 201430 346294 201498 346350
rect 201554 346294 201622 346350
rect 201678 346294 201774 346350
rect 201154 346226 201774 346294
rect 201154 346170 201250 346226
rect 201306 346170 201374 346226
rect 201430 346170 201498 346226
rect 201554 346170 201622 346226
rect 201678 346170 201774 346226
rect 201154 346102 201774 346170
rect 201154 346046 201250 346102
rect 201306 346046 201374 346102
rect 201430 346046 201498 346102
rect 201554 346046 201622 346102
rect 201678 346046 201774 346102
rect 201154 345978 201774 346046
rect 201154 345922 201250 345978
rect 201306 345922 201374 345978
rect 201430 345922 201498 345978
rect 201554 345922 201622 345978
rect 201678 345922 201774 345978
rect 201154 328350 201774 345922
rect 201154 328294 201250 328350
rect 201306 328294 201374 328350
rect 201430 328294 201498 328350
rect 201554 328294 201622 328350
rect 201678 328294 201774 328350
rect 201154 328226 201774 328294
rect 201154 328170 201250 328226
rect 201306 328170 201374 328226
rect 201430 328170 201498 328226
rect 201554 328170 201622 328226
rect 201678 328170 201774 328226
rect 201154 328102 201774 328170
rect 201154 328046 201250 328102
rect 201306 328046 201374 328102
rect 201430 328046 201498 328102
rect 201554 328046 201622 328102
rect 201678 328046 201774 328102
rect 201154 327978 201774 328046
rect 201154 327922 201250 327978
rect 201306 327922 201374 327978
rect 201430 327922 201498 327978
rect 201554 327922 201622 327978
rect 201678 327922 201774 327978
rect 201154 310350 201774 327922
rect 201154 310294 201250 310350
rect 201306 310294 201374 310350
rect 201430 310294 201498 310350
rect 201554 310294 201622 310350
rect 201678 310294 201774 310350
rect 201154 310226 201774 310294
rect 201154 310170 201250 310226
rect 201306 310170 201374 310226
rect 201430 310170 201498 310226
rect 201554 310170 201622 310226
rect 201678 310170 201774 310226
rect 201154 310102 201774 310170
rect 201154 310046 201250 310102
rect 201306 310046 201374 310102
rect 201430 310046 201498 310102
rect 201554 310046 201622 310102
rect 201678 310046 201774 310102
rect 201154 309978 201774 310046
rect 201154 309922 201250 309978
rect 201306 309922 201374 309978
rect 201430 309922 201498 309978
rect 201554 309922 201622 309978
rect 201678 309922 201774 309978
rect 201154 292350 201774 309922
rect 201154 292294 201250 292350
rect 201306 292294 201374 292350
rect 201430 292294 201498 292350
rect 201554 292294 201622 292350
rect 201678 292294 201774 292350
rect 201154 292226 201774 292294
rect 201154 292170 201250 292226
rect 201306 292170 201374 292226
rect 201430 292170 201498 292226
rect 201554 292170 201622 292226
rect 201678 292170 201774 292226
rect 201154 292102 201774 292170
rect 201154 292046 201250 292102
rect 201306 292046 201374 292102
rect 201430 292046 201498 292102
rect 201554 292046 201622 292102
rect 201678 292046 201774 292102
rect 201154 291978 201774 292046
rect 201154 291922 201250 291978
rect 201306 291922 201374 291978
rect 201430 291922 201498 291978
rect 201554 291922 201622 291978
rect 201678 291922 201774 291978
rect 201154 274350 201774 291922
rect 201154 274294 201250 274350
rect 201306 274294 201374 274350
rect 201430 274294 201498 274350
rect 201554 274294 201622 274350
rect 201678 274294 201774 274350
rect 201154 274226 201774 274294
rect 201154 274170 201250 274226
rect 201306 274170 201374 274226
rect 201430 274170 201498 274226
rect 201554 274170 201622 274226
rect 201678 274170 201774 274226
rect 201154 274102 201774 274170
rect 201154 274046 201250 274102
rect 201306 274046 201374 274102
rect 201430 274046 201498 274102
rect 201554 274046 201622 274102
rect 201678 274046 201774 274102
rect 201154 273978 201774 274046
rect 201154 273922 201250 273978
rect 201306 273922 201374 273978
rect 201430 273922 201498 273978
rect 201554 273922 201622 273978
rect 201678 273922 201774 273978
rect 201154 256350 201774 273922
rect 201154 256294 201250 256350
rect 201306 256294 201374 256350
rect 201430 256294 201498 256350
rect 201554 256294 201622 256350
rect 201678 256294 201774 256350
rect 201154 256226 201774 256294
rect 201154 256170 201250 256226
rect 201306 256170 201374 256226
rect 201430 256170 201498 256226
rect 201554 256170 201622 256226
rect 201678 256170 201774 256226
rect 201154 256102 201774 256170
rect 201154 256046 201250 256102
rect 201306 256046 201374 256102
rect 201430 256046 201498 256102
rect 201554 256046 201622 256102
rect 201678 256046 201774 256102
rect 201154 255978 201774 256046
rect 201154 255922 201250 255978
rect 201306 255922 201374 255978
rect 201430 255922 201498 255978
rect 201554 255922 201622 255978
rect 201678 255922 201774 255978
rect 201154 238350 201774 255922
rect 219154 597212 219774 598268
rect 219154 597156 219250 597212
rect 219306 597156 219374 597212
rect 219430 597156 219498 597212
rect 219554 597156 219622 597212
rect 219678 597156 219774 597212
rect 219154 597088 219774 597156
rect 219154 597032 219250 597088
rect 219306 597032 219374 597088
rect 219430 597032 219498 597088
rect 219554 597032 219622 597088
rect 219678 597032 219774 597088
rect 219154 596964 219774 597032
rect 219154 596908 219250 596964
rect 219306 596908 219374 596964
rect 219430 596908 219498 596964
rect 219554 596908 219622 596964
rect 219678 596908 219774 596964
rect 219154 596840 219774 596908
rect 219154 596784 219250 596840
rect 219306 596784 219374 596840
rect 219430 596784 219498 596840
rect 219554 596784 219622 596840
rect 219678 596784 219774 596840
rect 219154 580350 219774 596784
rect 219154 580294 219250 580350
rect 219306 580294 219374 580350
rect 219430 580294 219498 580350
rect 219554 580294 219622 580350
rect 219678 580294 219774 580350
rect 219154 580226 219774 580294
rect 219154 580170 219250 580226
rect 219306 580170 219374 580226
rect 219430 580170 219498 580226
rect 219554 580170 219622 580226
rect 219678 580170 219774 580226
rect 219154 580102 219774 580170
rect 219154 580046 219250 580102
rect 219306 580046 219374 580102
rect 219430 580046 219498 580102
rect 219554 580046 219622 580102
rect 219678 580046 219774 580102
rect 219154 579978 219774 580046
rect 219154 579922 219250 579978
rect 219306 579922 219374 579978
rect 219430 579922 219498 579978
rect 219554 579922 219622 579978
rect 219678 579922 219774 579978
rect 219154 562350 219774 579922
rect 219154 562294 219250 562350
rect 219306 562294 219374 562350
rect 219430 562294 219498 562350
rect 219554 562294 219622 562350
rect 219678 562294 219774 562350
rect 219154 562226 219774 562294
rect 219154 562170 219250 562226
rect 219306 562170 219374 562226
rect 219430 562170 219498 562226
rect 219554 562170 219622 562226
rect 219678 562170 219774 562226
rect 219154 562102 219774 562170
rect 219154 562046 219250 562102
rect 219306 562046 219374 562102
rect 219430 562046 219498 562102
rect 219554 562046 219622 562102
rect 219678 562046 219774 562102
rect 219154 561978 219774 562046
rect 219154 561922 219250 561978
rect 219306 561922 219374 561978
rect 219430 561922 219498 561978
rect 219554 561922 219622 561978
rect 219678 561922 219774 561978
rect 219154 544350 219774 561922
rect 219154 544294 219250 544350
rect 219306 544294 219374 544350
rect 219430 544294 219498 544350
rect 219554 544294 219622 544350
rect 219678 544294 219774 544350
rect 219154 544226 219774 544294
rect 219154 544170 219250 544226
rect 219306 544170 219374 544226
rect 219430 544170 219498 544226
rect 219554 544170 219622 544226
rect 219678 544170 219774 544226
rect 219154 544102 219774 544170
rect 219154 544046 219250 544102
rect 219306 544046 219374 544102
rect 219430 544046 219498 544102
rect 219554 544046 219622 544102
rect 219678 544046 219774 544102
rect 219154 543978 219774 544046
rect 219154 543922 219250 543978
rect 219306 543922 219374 543978
rect 219430 543922 219498 543978
rect 219554 543922 219622 543978
rect 219678 543922 219774 543978
rect 219154 526350 219774 543922
rect 219154 526294 219250 526350
rect 219306 526294 219374 526350
rect 219430 526294 219498 526350
rect 219554 526294 219622 526350
rect 219678 526294 219774 526350
rect 219154 526226 219774 526294
rect 219154 526170 219250 526226
rect 219306 526170 219374 526226
rect 219430 526170 219498 526226
rect 219554 526170 219622 526226
rect 219678 526170 219774 526226
rect 219154 526102 219774 526170
rect 219154 526046 219250 526102
rect 219306 526046 219374 526102
rect 219430 526046 219498 526102
rect 219554 526046 219622 526102
rect 219678 526046 219774 526102
rect 219154 525978 219774 526046
rect 219154 525922 219250 525978
rect 219306 525922 219374 525978
rect 219430 525922 219498 525978
rect 219554 525922 219622 525978
rect 219678 525922 219774 525978
rect 219154 508350 219774 525922
rect 219154 508294 219250 508350
rect 219306 508294 219374 508350
rect 219430 508294 219498 508350
rect 219554 508294 219622 508350
rect 219678 508294 219774 508350
rect 219154 508226 219774 508294
rect 219154 508170 219250 508226
rect 219306 508170 219374 508226
rect 219430 508170 219498 508226
rect 219554 508170 219622 508226
rect 219678 508170 219774 508226
rect 219154 508102 219774 508170
rect 219154 508046 219250 508102
rect 219306 508046 219374 508102
rect 219430 508046 219498 508102
rect 219554 508046 219622 508102
rect 219678 508046 219774 508102
rect 219154 507978 219774 508046
rect 219154 507922 219250 507978
rect 219306 507922 219374 507978
rect 219430 507922 219498 507978
rect 219554 507922 219622 507978
rect 219678 507922 219774 507978
rect 219154 490350 219774 507922
rect 219154 490294 219250 490350
rect 219306 490294 219374 490350
rect 219430 490294 219498 490350
rect 219554 490294 219622 490350
rect 219678 490294 219774 490350
rect 219154 490226 219774 490294
rect 219154 490170 219250 490226
rect 219306 490170 219374 490226
rect 219430 490170 219498 490226
rect 219554 490170 219622 490226
rect 219678 490170 219774 490226
rect 219154 490102 219774 490170
rect 219154 490046 219250 490102
rect 219306 490046 219374 490102
rect 219430 490046 219498 490102
rect 219554 490046 219622 490102
rect 219678 490046 219774 490102
rect 219154 489978 219774 490046
rect 219154 489922 219250 489978
rect 219306 489922 219374 489978
rect 219430 489922 219498 489978
rect 219554 489922 219622 489978
rect 219678 489922 219774 489978
rect 219154 472350 219774 489922
rect 219154 472294 219250 472350
rect 219306 472294 219374 472350
rect 219430 472294 219498 472350
rect 219554 472294 219622 472350
rect 219678 472294 219774 472350
rect 219154 472226 219774 472294
rect 219154 472170 219250 472226
rect 219306 472170 219374 472226
rect 219430 472170 219498 472226
rect 219554 472170 219622 472226
rect 219678 472170 219774 472226
rect 219154 472102 219774 472170
rect 219154 472046 219250 472102
rect 219306 472046 219374 472102
rect 219430 472046 219498 472102
rect 219554 472046 219622 472102
rect 219678 472046 219774 472102
rect 219154 471978 219774 472046
rect 219154 471922 219250 471978
rect 219306 471922 219374 471978
rect 219430 471922 219498 471978
rect 219554 471922 219622 471978
rect 219678 471922 219774 471978
rect 219154 454350 219774 471922
rect 219154 454294 219250 454350
rect 219306 454294 219374 454350
rect 219430 454294 219498 454350
rect 219554 454294 219622 454350
rect 219678 454294 219774 454350
rect 219154 454226 219774 454294
rect 219154 454170 219250 454226
rect 219306 454170 219374 454226
rect 219430 454170 219498 454226
rect 219554 454170 219622 454226
rect 219678 454170 219774 454226
rect 219154 454102 219774 454170
rect 219154 454046 219250 454102
rect 219306 454046 219374 454102
rect 219430 454046 219498 454102
rect 219554 454046 219622 454102
rect 219678 454046 219774 454102
rect 219154 453978 219774 454046
rect 219154 453922 219250 453978
rect 219306 453922 219374 453978
rect 219430 453922 219498 453978
rect 219554 453922 219622 453978
rect 219678 453922 219774 453978
rect 219154 436350 219774 453922
rect 219154 436294 219250 436350
rect 219306 436294 219374 436350
rect 219430 436294 219498 436350
rect 219554 436294 219622 436350
rect 219678 436294 219774 436350
rect 219154 436226 219774 436294
rect 219154 436170 219250 436226
rect 219306 436170 219374 436226
rect 219430 436170 219498 436226
rect 219554 436170 219622 436226
rect 219678 436170 219774 436226
rect 219154 436102 219774 436170
rect 219154 436046 219250 436102
rect 219306 436046 219374 436102
rect 219430 436046 219498 436102
rect 219554 436046 219622 436102
rect 219678 436046 219774 436102
rect 219154 435978 219774 436046
rect 219154 435922 219250 435978
rect 219306 435922 219374 435978
rect 219430 435922 219498 435978
rect 219554 435922 219622 435978
rect 219678 435922 219774 435978
rect 219154 418350 219774 435922
rect 219154 418294 219250 418350
rect 219306 418294 219374 418350
rect 219430 418294 219498 418350
rect 219554 418294 219622 418350
rect 219678 418294 219774 418350
rect 219154 418226 219774 418294
rect 219154 418170 219250 418226
rect 219306 418170 219374 418226
rect 219430 418170 219498 418226
rect 219554 418170 219622 418226
rect 219678 418170 219774 418226
rect 219154 418102 219774 418170
rect 219154 418046 219250 418102
rect 219306 418046 219374 418102
rect 219430 418046 219498 418102
rect 219554 418046 219622 418102
rect 219678 418046 219774 418102
rect 219154 417978 219774 418046
rect 219154 417922 219250 417978
rect 219306 417922 219374 417978
rect 219430 417922 219498 417978
rect 219554 417922 219622 417978
rect 219678 417922 219774 417978
rect 219154 400350 219774 417922
rect 219154 400294 219250 400350
rect 219306 400294 219374 400350
rect 219430 400294 219498 400350
rect 219554 400294 219622 400350
rect 219678 400294 219774 400350
rect 219154 400226 219774 400294
rect 219154 400170 219250 400226
rect 219306 400170 219374 400226
rect 219430 400170 219498 400226
rect 219554 400170 219622 400226
rect 219678 400170 219774 400226
rect 219154 400102 219774 400170
rect 219154 400046 219250 400102
rect 219306 400046 219374 400102
rect 219430 400046 219498 400102
rect 219554 400046 219622 400102
rect 219678 400046 219774 400102
rect 219154 399978 219774 400046
rect 219154 399922 219250 399978
rect 219306 399922 219374 399978
rect 219430 399922 219498 399978
rect 219554 399922 219622 399978
rect 219678 399922 219774 399978
rect 219154 382350 219774 399922
rect 219154 382294 219250 382350
rect 219306 382294 219374 382350
rect 219430 382294 219498 382350
rect 219554 382294 219622 382350
rect 219678 382294 219774 382350
rect 219154 382226 219774 382294
rect 219154 382170 219250 382226
rect 219306 382170 219374 382226
rect 219430 382170 219498 382226
rect 219554 382170 219622 382226
rect 219678 382170 219774 382226
rect 219154 382102 219774 382170
rect 219154 382046 219250 382102
rect 219306 382046 219374 382102
rect 219430 382046 219498 382102
rect 219554 382046 219622 382102
rect 219678 382046 219774 382102
rect 219154 381978 219774 382046
rect 219154 381922 219250 381978
rect 219306 381922 219374 381978
rect 219430 381922 219498 381978
rect 219554 381922 219622 381978
rect 219678 381922 219774 381978
rect 219154 364350 219774 381922
rect 219154 364294 219250 364350
rect 219306 364294 219374 364350
rect 219430 364294 219498 364350
rect 219554 364294 219622 364350
rect 219678 364294 219774 364350
rect 219154 364226 219774 364294
rect 219154 364170 219250 364226
rect 219306 364170 219374 364226
rect 219430 364170 219498 364226
rect 219554 364170 219622 364226
rect 219678 364170 219774 364226
rect 219154 364102 219774 364170
rect 219154 364046 219250 364102
rect 219306 364046 219374 364102
rect 219430 364046 219498 364102
rect 219554 364046 219622 364102
rect 219678 364046 219774 364102
rect 219154 363978 219774 364046
rect 219154 363922 219250 363978
rect 219306 363922 219374 363978
rect 219430 363922 219498 363978
rect 219554 363922 219622 363978
rect 219678 363922 219774 363978
rect 219154 346350 219774 363922
rect 219154 346294 219250 346350
rect 219306 346294 219374 346350
rect 219430 346294 219498 346350
rect 219554 346294 219622 346350
rect 219678 346294 219774 346350
rect 219154 346226 219774 346294
rect 219154 346170 219250 346226
rect 219306 346170 219374 346226
rect 219430 346170 219498 346226
rect 219554 346170 219622 346226
rect 219678 346170 219774 346226
rect 219154 346102 219774 346170
rect 219154 346046 219250 346102
rect 219306 346046 219374 346102
rect 219430 346046 219498 346102
rect 219554 346046 219622 346102
rect 219678 346046 219774 346102
rect 219154 345978 219774 346046
rect 219154 345922 219250 345978
rect 219306 345922 219374 345978
rect 219430 345922 219498 345978
rect 219554 345922 219622 345978
rect 219678 345922 219774 345978
rect 219154 328350 219774 345922
rect 219154 328294 219250 328350
rect 219306 328294 219374 328350
rect 219430 328294 219498 328350
rect 219554 328294 219622 328350
rect 219678 328294 219774 328350
rect 219154 328226 219774 328294
rect 219154 328170 219250 328226
rect 219306 328170 219374 328226
rect 219430 328170 219498 328226
rect 219554 328170 219622 328226
rect 219678 328170 219774 328226
rect 219154 328102 219774 328170
rect 219154 328046 219250 328102
rect 219306 328046 219374 328102
rect 219430 328046 219498 328102
rect 219554 328046 219622 328102
rect 219678 328046 219774 328102
rect 219154 327978 219774 328046
rect 219154 327922 219250 327978
rect 219306 327922 219374 327978
rect 219430 327922 219498 327978
rect 219554 327922 219622 327978
rect 219678 327922 219774 327978
rect 219154 310350 219774 327922
rect 219154 310294 219250 310350
rect 219306 310294 219374 310350
rect 219430 310294 219498 310350
rect 219554 310294 219622 310350
rect 219678 310294 219774 310350
rect 219154 310226 219774 310294
rect 219154 310170 219250 310226
rect 219306 310170 219374 310226
rect 219430 310170 219498 310226
rect 219554 310170 219622 310226
rect 219678 310170 219774 310226
rect 219154 310102 219774 310170
rect 219154 310046 219250 310102
rect 219306 310046 219374 310102
rect 219430 310046 219498 310102
rect 219554 310046 219622 310102
rect 219678 310046 219774 310102
rect 219154 309978 219774 310046
rect 219154 309922 219250 309978
rect 219306 309922 219374 309978
rect 219430 309922 219498 309978
rect 219554 309922 219622 309978
rect 219678 309922 219774 309978
rect 219154 292350 219774 309922
rect 219154 292294 219250 292350
rect 219306 292294 219374 292350
rect 219430 292294 219498 292350
rect 219554 292294 219622 292350
rect 219678 292294 219774 292350
rect 219154 292226 219774 292294
rect 219154 292170 219250 292226
rect 219306 292170 219374 292226
rect 219430 292170 219498 292226
rect 219554 292170 219622 292226
rect 219678 292170 219774 292226
rect 219154 292102 219774 292170
rect 219154 292046 219250 292102
rect 219306 292046 219374 292102
rect 219430 292046 219498 292102
rect 219554 292046 219622 292102
rect 219678 292046 219774 292102
rect 219154 291978 219774 292046
rect 219154 291922 219250 291978
rect 219306 291922 219374 291978
rect 219430 291922 219498 291978
rect 219554 291922 219622 291978
rect 219678 291922 219774 291978
rect 219154 274350 219774 291922
rect 219154 274294 219250 274350
rect 219306 274294 219374 274350
rect 219430 274294 219498 274350
rect 219554 274294 219622 274350
rect 219678 274294 219774 274350
rect 219154 274226 219774 274294
rect 219154 274170 219250 274226
rect 219306 274170 219374 274226
rect 219430 274170 219498 274226
rect 219554 274170 219622 274226
rect 219678 274170 219774 274226
rect 219154 274102 219774 274170
rect 219154 274046 219250 274102
rect 219306 274046 219374 274102
rect 219430 274046 219498 274102
rect 219554 274046 219622 274102
rect 219678 274046 219774 274102
rect 219154 273978 219774 274046
rect 219154 273922 219250 273978
rect 219306 273922 219374 273978
rect 219430 273922 219498 273978
rect 219554 273922 219622 273978
rect 219678 273922 219774 273978
rect 219154 256350 219774 273922
rect 219154 256294 219250 256350
rect 219306 256294 219374 256350
rect 219430 256294 219498 256350
rect 219554 256294 219622 256350
rect 219678 256294 219774 256350
rect 219154 256226 219774 256294
rect 219154 256170 219250 256226
rect 219306 256170 219374 256226
rect 219430 256170 219498 256226
rect 219554 256170 219622 256226
rect 219678 256170 219774 256226
rect 219154 256102 219774 256170
rect 219154 256046 219250 256102
rect 219306 256046 219374 256102
rect 219430 256046 219498 256102
rect 219554 256046 219622 256102
rect 219678 256046 219774 256102
rect 219154 255978 219774 256046
rect 219154 255922 219250 255978
rect 219306 255922 219374 255978
rect 219430 255922 219498 255978
rect 219554 255922 219622 255978
rect 219678 255922 219774 255978
rect 201154 238294 201250 238350
rect 201306 238294 201374 238350
rect 201430 238294 201498 238350
rect 201554 238294 201622 238350
rect 201678 238294 201774 238350
rect 201154 238226 201774 238294
rect 201154 238170 201250 238226
rect 201306 238170 201374 238226
rect 201430 238170 201498 238226
rect 201554 238170 201622 238226
rect 201678 238170 201774 238226
rect 201154 238102 201774 238170
rect 201154 238046 201250 238102
rect 201306 238046 201374 238102
rect 201430 238046 201498 238102
rect 201554 238046 201622 238102
rect 201678 238046 201774 238102
rect 201154 237978 201774 238046
rect 201154 237922 201250 237978
rect 201306 237922 201374 237978
rect 201430 237922 201498 237978
rect 201554 237922 201622 237978
rect 201678 237922 201774 237978
rect 193228 229348 193284 229358
rect 193228 227780 193284 229292
rect 193228 227714 193284 227724
rect 183154 220294 183250 220350
rect 183306 220294 183374 220350
rect 183430 220294 183498 220350
rect 183554 220294 183622 220350
rect 183678 220294 183774 220350
rect 183154 220226 183774 220294
rect 183154 220170 183250 220226
rect 183306 220170 183374 220226
rect 183430 220170 183498 220226
rect 183554 220170 183622 220226
rect 183678 220170 183774 220226
rect 183154 220102 183774 220170
rect 183154 220046 183250 220102
rect 183306 220046 183374 220102
rect 183430 220046 183498 220102
rect 183554 220046 183622 220102
rect 183678 220046 183774 220102
rect 183154 219978 183774 220046
rect 183154 219922 183250 219978
rect 183306 219922 183374 219978
rect 183430 219922 183498 219978
rect 183554 219922 183622 219978
rect 183678 219922 183774 219978
rect 183154 219134 183774 219922
rect 187328 220350 187648 220384
rect 187328 220294 187398 220350
rect 187454 220294 187522 220350
rect 187578 220294 187648 220350
rect 187328 220226 187648 220294
rect 187328 220170 187398 220226
rect 187454 220170 187522 220226
rect 187578 220170 187648 220226
rect 187328 220102 187648 220170
rect 187328 220046 187398 220102
rect 187454 220046 187522 220102
rect 187578 220046 187648 220102
rect 187328 219978 187648 220046
rect 187328 219922 187398 219978
rect 187454 219922 187522 219978
rect 187578 219922 187648 219978
rect 187328 219888 187648 219922
rect 201154 220350 201774 237922
rect 202688 226350 203008 226384
rect 202688 226294 202758 226350
rect 202814 226294 202882 226350
rect 202938 226294 203008 226350
rect 202688 226226 203008 226294
rect 202688 226170 202758 226226
rect 202814 226170 202882 226226
rect 202938 226170 203008 226226
rect 202688 226102 203008 226170
rect 202688 226046 202758 226102
rect 202814 226046 202882 226102
rect 202938 226046 203008 226102
rect 202688 225978 203008 226046
rect 202688 225922 202758 225978
rect 202814 225922 202882 225978
rect 202938 225922 203008 225978
rect 202688 225888 203008 225922
rect 204874 226350 205494 242964
rect 204874 226294 204970 226350
rect 205026 226294 205094 226350
rect 205150 226294 205218 226350
rect 205274 226294 205342 226350
rect 205398 226294 205494 226350
rect 204874 226226 205494 226294
rect 204874 226170 204970 226226
rect 205026 226170 205094 226226
rect 205150 226170 205218 226226
rect 205274 226170 205342 226226
rect 205398 226170 205494 226226
rect 204874 226102 205494 226170
rect 204874 226046 204970 226102
rect 205026 226046 205094 226102
rect 205150 226046 205218 226102
rect 205274 226046 205342 226102
rect 205398 226046 205494 226102
rect 204874 225978 205494 226046
rect 204874 225922 204970 225978
rect 205026 225922 205094 225978
rect 205150 225922 205218 225978
rect 205274 225922 205342 225978
rect 205398 225922 205494 225978
rect 201154 220294 201250 220350
rect 201306 220294 201374 220350
rect 201430 220294 201498 220350
rect 201554 220294 201622 220350
rect 201678 220294 201774 220350
rect 201154 220226 201774 220294
rect 201154 220170 201250 220226
rect 201306 220170 201374 220226
rect 201430 220170 201498 220226
rect 201554 220170 201622 220226
rect 201678 220170 201774 220226
rect 201154 220102 201774 220170
rect 201154 220046 201250 220102
rect 201306 220046 201374 220102
rect 201430 220046 201498 220102
rect 201554 220046 201622 220102
rect 201678 220046 201774 220102
rect 201154 219978 201774 220046
rect 201154 219922 201250 219978
rect 201306 219922 201374 219978
rect 201430 219922 201498 219978
rect 201554 219922 201622 219978
rect 201678 219922 201774 219978
rect 201154 219134 201774 219922
rect 204874 219134 205494 225922
rect 219154 238350 219774 255922
rect 219154 238294 219250 238350
rect 219306 238294 219374 238350
rect 219430 238294 219498 238350
rect 219554 238294 219622 238350
rect 219678 238294 219774 238350
rect 219154 238226 219774 238294
rect 219154 238170 219250 238226
rect 219306 238170 219374 238226
rect 219430 238170 219498 238226
rect 219554 238170 219622 238226
rect 219678 238170 219774 238226
rect 219154 238102 219774 238170
rect 219154 238046 219250 238102
rect 219306 238046 219374 238102
rect 219430 238046 219498 238102
rect 219554 238046 219622 238102
rect 219678 238046 219774 238102
rect 219154 237978 219774 238046
rect 219154 237922 219250 237978
rect 219306 237922 219374 237978
rect 219430 237922 219498 237978
rect 219554 237922 219622 237978
rect 219678 237922 219774 237978
rect 218048 220350 218368 220384
rect 218048 220294 218118 220350
rect 218174 220294 218242 220350
rect 218298 220294 218368 220350
rect 218048 220226 218368 220294
rect 218048 220170 218118 220226
rect 218174 220170 218242 220226
rect 218298 220170 218368 220226
rect 218048 220102 218368 220170
rect 218048 220046 218118 220102
rect 218174 220046 218242 220102
rect 218298 220046 218368 220102
rect 218048 219978 218368 220046
rect 218048 219922 218118 219978
rect 218174 219922 218242 219978
rect 218298 219922 218368 219978
rect 218048 219888 218368 219922
rect 219154 220350 219774 237922
rect 219154 220294 219250 220350
rect 219306 220294 219374 220350
rect 219430 220294 219498 220350
rect 219554 220294 219622 220350
rect 219678 220294 219774 220350
rect 219154 220226 219774 220294
rect 219154 220170 219250 220226
rect 219306 220170 219374 220226
rect 219430 220170 219498 220226
rect 219554 220170 219622 220226
rect 219678 220170 219774 220226
rect 219154 220102 219774 220170
rect 219154 220046 219250 220102
rect 219306 220046 219374 220102
rect 219430 220046 219498 220102
rect 219554 220046 219622 220102
rect 219678 220046 219774 220102
rect 219154 219978 219774 220046
rect 219154 219922 219250 219978
rect 219306 219922 219374 219978
rect 219430 219922 219498 219978
rect 219554 219922 219622 219978
rect 219678 219922 219774 219978
rect 219154 219134 219774 219922
rect 222874 598172 223494 598268
rect 222874 598116 222970 598172
rect 223026 598116 223094 598172
rect 223150 598116 223218 598172
rect 223274 598116 223342 598172
rect 223398 598116 223494 598172
rect 222874 598048 223494 598116
rect 222874 597992 222970 598048
rect 223026 597992 223094 598048
rect 223150 597992 223218 598048
rect 223274 597992 223342 598048
rect 223398 597992 223494 598048
rect 222874 597924 223494 597992
rect 222874 597868 222970 597924
rect 223026 597868 223094 597924
rect 223150 597868 223218 597924
rect 223274 597868 223342 597924
rect 223398 597868 223494 597924
rect 222874 597800 223494 597868
rect 222874 597744 222970 597800
rect 223026 597744 223094 597800
rect 223150 597744 223218 597800
rect 223274 597744 223342 597800
rect 223398 597744 223494 597800
rect 222874 586350 223494 597744
rect 222874 586294 222970 586350
rect 223026 586294 223094 586350
rect 223150 586294 223218 586350
rect 223274 586294 223342 586350
rect 223398 586294 223494 586350
rect 222874 586226 223494 586294
rect 222874 586170 222970 586226
rect 223026 586170 223094 586226
rect 223150 586170 223218 586226
rect 223274 586170 223342 586226
rect 223398 586170 223494 586226
rect 222874 586102 223494 586170
rect 222874 586046 222970 586102
rect 223026 586046 223094 586102
rect 223150 586046 223218 586102
rect 223274 586046 223342 586102
rect 223398 586046 223494 586102
rect 222874 585978 223494 586046
rect 222874 585922 222970 585978
rect 223026 585922 223094 585978
rect 223150 585922 223218 585978
rect 223274 585922 223342 585978
rect 223398 585922 223494 585978
rect 222874 568350 223494 585922
rect 222874 568294 222970 568350
rect 223026 568294 223094 568350
rect 223150 568294 223218 568350
rect 223274 568294 223342 568350
rect 223398 568294 223494 568350
rect 222874 568226 223494 568294
rect 222874 568170 222970 568226
rect 223026 568170 223094 568226
rect 223150 568170 223218 568226
rect 223274 568170 223342 568226
rect 223398 568170 223494 568226
rect 222874 568102 223494 568170
rect 222874 568046 222970 568102
rect 223026 568046 223094 568102
rect 223150 568046 223218 568102
rect 223274 568046 223342 568102
rect 223398 568046 223494 568102
rect 222874 567978 223494 568046
rect 222874 567922 222970 567978
rect 223026 567922 223094 567978
rect 223150 567922 223218 567978
rect 223274 567922 223342 567978
rect 223398 567922 223494 567978
rect 222874 550350 223494 567922
rect 222874 550294 222970 550350
rect 223026 550294 223094 550350
rect 223150 550294 223218 550350
rect 223274 550294 223342 550350
rect 223398 550294 223494 550350
rect 222874 550226 223494 550294
rect 222874 550170 222970 550226
rect 223026 550170 223094 550226
rect 223150 550170 223218 550226
rect 223274 550170 223342 550226
rect 223398 550170 223494 550226
rect 222874 550102 223494 550170
rect 222874 550046 222970 550102
rect 223026 550046 223094 550102
rect 223150 550046 223218 550102
rect 223274 550046 223342 550102
rect 223398 550046 223494 550102
rect 222874 549978 223494 550046
rect 222874 549922 222970 549978
rect 223026 549922 223094 549978
rect 223150 549922 223218 549978
rect 223274 549922 223342 549978
rect 223398 549922 223494 549978
rect 222874 532350 223494 549922
rect 222874 532294 222970 532350
rect 223026 532294 223094 532350
rect 223150 532294 223218 532350
rect 223274 532294 223342 532350
rect 223398 532294 223494 532350
rect 222874 532226 223494 532294
rect 222874 532170 222970 532226
rect 223026 532170 223094 532226
rect 223150 532170 223218 532226
rect 223274 532170 223342 532226
rect 223398 532170 223494 532226
rect 222874 532102 223494 532170
rect 222874 532046 222970 532102
rect 223026 532046 223094 532102
rect 223150 532046 223218 532102
rect 223274 532046 223342 532102
rect 223398 532046 223494 532102
rect 222874 531978 223494 532046
rect 222874 531922 222970 531978
rect 223026 531922 223094 531978
rect 223150 531922 223218 531978
rect 223274 531922 223342 531978
rect 223398 531922 223494 531978
rect 222874 514350 223494 531922
rect 222874 514294 222970 514350
rect 223026 514294 223094 514350
rect 223150 514294 223218 514350
rect 223274 514294 223342 514350
rect 223398 514294 223494 514350
rect 222874 514226 223494 514294
rect 222874 514170 222970 514226
rect 223026 514170 223094 514226
rect 223150 514170 223218 514226
rect 223274 514170 223342 514226
rect 223398 514170 223494 514226
rect 222874 514102 223494 514170
rect 222874 514046 222970 514102
rect 223026 514046 223094 514102
rect 223150 514046 223218 514102
rect 223274 514046 223342 514102
rect 223398 514046 223494 514102
rect 222874 513978 223494 514046
rect 222874 513922 222970 513978
rect 223026 513922 223094 513978
rect 223150 513922 223218 513978
rect 223274 513922 223342 513978
rect 223398 513922 223494 513978
rect 222874 496350 223494 513922
rect 222874 496294 222970 496350
rect 223026 496294 223094 496350
rect 223150 496294 223218 496350
rect 223274 496294 223342 496350
rect 223398 496294 223494 496350
rect 222874 496226 223494 496294
rect 222874 496170 222970 496226
rect 223026 496170 223094 496226
rect 223150 496170 223218 496226
rect 223274 496170 223342 496226
rect 223398 496170 223494 496226
rect 222874 496102 223494 496170
rect 222874 496046 222970 496102
rect 223026 496046 223094 496102
rect 223150 496046 223218 496102
rect 223274 496046 223342 496102
rect 223398 496046 223494 496102
rect 222874 495978 223494 496046
rect 222874 495922 222970 495978
rect 223026 495922 223094 495978
rect 223150 495922 223218 495978
rect 223274 495922 223342 495978
rect 223398 495922 223494 495978
rect 222874 478350 223494 495922
rect 222874 478294 222970 478350
rect 223026 478294 223094 478350
rect 223150 478294 223218 478350
rect 223274 478294 223342 478350
rect 223398 478294 223494 478350
rect 222874 478226 223494 478294
rect 222874 478170 222970 478226
rect 223026 478170 223094 478226
rect 223150 478170 223218 478226
rect 223274 478170 223342 478226
rect 223398 478170 223494 478226
rect 222874 478102 223494 478170
rect 222874 478046 222970 478102
rect 223026 478046 223094 478102
rect 223150 478046 223218 478102
rect 223274 478046 223342 478102
rect 223398 478046 223494 478102
rect 222874 477978 223494 478046
rect 222874 477922 222970 477978
rect 223026 477922 223094 477978
rect 223150 477922 223218 477978
rect 223274 477922 223342 477978
rect 223398 477922 223494 477978
rect 222874 460350 223494 477922
rect 222874 460294 222970 460350
rect 223026 460294 223094 460350
rect 223150 460294 223218 460350
rect 223274 460294 223342 460350
rect 223398 460294 223494 460350
rect 222874 460226 223494 460294
rect 222874 460170 222970 460226
rect 223026 460170 223094 460226
rect 223150 460170 223218 460226
rect 223274 460170 223342 460226
rect 223398 460170 223494 460226
rect 222874 460102 223494 460170
rect 222874 460046 222970 460102
rect 223026 460046 223094 460102
rect 223150 460046 223218 460102
rect 223274 460046 223342 460102
rect 223398 460046 223494 460102
rect 222874 459978 223494 460046
rect 222874 459922 222970 459978
rect 223026 459922 223094 459978
rect 223150 459922 223218 459978
rect 223274 459922 223342 459978
rect 223398 459922 223494 459978
rect 222874 442350 223494 459922
rect 222874 442294 222970 442350
rect 223026 442294 223094 442350
rect 223150 442294 223218 442350
rect 223274 442294 223342 442350
rect 223398 442294 223494 442350
rect 222874 442226 223494 442294
rect 222874 442170 222970 442226
rect 223026 442170 223094 442226
rect 223150 442170 223218 442226
rect 223274 442170 223342 442226
rect 223398 442170 223494 442226
rect 222874 442102 223494 442170
rect 222874 442046 222970 442102
rect 223026 442046 223094 442102
rect 223150 442046 223218 442102
rect 223274 442046 223342 442102
rect 223398 442046 223494 442102
rect 222874 441978 223494 442046
rect 222874 441922 222970 441978
rect 223026 441922 223094 441978
rect 223150 441922 223218 441978
rect 223274 441922 223342 441978
rect 223398 441922 223494 441978
rect 222874 424350 223494 441922
rect 222874 424294 222970 424350
rect 223026 424294 223094 424350
rect 223150 424294 223218 424350
rect 223274 424294 223342 424350
rect 223398 424294 223494 424350
rect 222874 424226 223494 424294
rect 222874 424170 222970 424226
rect 223026 424170 223094 424226
rect 223150 424170 223218 424226
rect 223274 424170 223342 424226
rect 223398 424170 223494 424226
rect 222874 424102 223494 424170
rect 222874 424046 222970 424102
rect 223026 424046 223094 424102
rect 223150 424046 223218 424102
rect 223274 424046 223342 424102
rect 223398 424046 223494 424102
rect 222874 423978 223494 424046
rect 222874 423922 222970 423978
rect 223026 423922 223094 423978
rect 223150 423922 223218 423978
rect 223274 423922 223342 423978
rect 223398 423922 223494 423978
rect 222874 406350 223494 423922
rect 222874 406294 222970 406350
rect 223026 406294 223094 406350
rect 223150 406294 223218 406350
rect 223274 406294 223342 406350
rect 223398 406294 223494 406350
rect 222874 406226 223494 406294
rect 222874 406170 222970 406226
rect 223026 406170 223094 406226
rect 223150 406170 223218 406226
rect 223274 406170 223342 406226
rect 223398 406170 223494 406226
rect 222874 406102 223494 406170
rect 222874 406046 222970 406102
rect 223026 406046 223094 406102
rect 223150 406046 223218 406102
rect 223274 406046 223342 406102
rect 223398 406046 223494 406102
rect 222874 405978 223494 406046
rect 222874 405922 222970 405978
rect 223026 405922 223094 405978
rect 223150 405922 223218 405978
rect 223274 405922 223342 405978
rect 223398 405922 223494 405978
rect 222874 388350 223494 405922
rect 222874 388294 222970 388350
rect 223026 388294 223094 388350
rect 223150 388294 223218 388350
rect 223274 388294 223342 388350
rect 223398 388294 223494 388350
rect 222874 388226 223494 388294
rect 222874 388170 222970 388226
rect 223026 388170 223094 388226
rect 223150 388170 223218 388226
rect 223274 388170 223342 388226
rect 223398 388170 223494 388226
rect 222874 388102 223494 388170
rect 222874 388046 222970 388102
rect 223026 388046 223094 388102
rect 223150 388046 223218 388102
rect 223274 388046 223342 388102
rect 223398 388046 223494 388102
rect 222874 387978 223494 388046
rect 222874 387922 222970 387978
rect 223026 387922 223094 387978
rect 223150 387922 223218 387978
rect 223274 387922 223342 387978
rect 223398 387922 223494 387978
rect 222874 370350 223494 387922
rect 222874 370294 222970 370350
rect 223026 370294 223094 370350
rect 223150 370294 223218 370350
rect 223274 370294 223342 370350
rect 223398 370294 223494 370350
rect 222874 370226 223494 370294
rect 222874 370170 222970 370226
rect 223026 370170 223094 370226
rect 223150 370170 223218 370226
rect 223274 370170 223342 370226
rect 223398 370170 223494 370226
rect 222874 370102 223494 370170
rect 222874 370046 222970 370102
rect 223026 370046 223094 370102
rect 223150 370046 223218 370102
rect 223274 370046 223342 370102
rect 223398 370046 223494 370102
rect 222874 369978 223494 370046
rect 222874 369922 222970 369978
rect 223026 369922 223094 369978
rect 223150 369922 223218 369978
rect 223274 369922 223342 369978
rect 223398 369922 223494 369978
rect 222874 352350 223494 369922
rect 222874 352294 222970 352350
rect 223026 352294 223094 352350
rect 223150 352294 223218 352350
rect 223274 352294 223342 352350
rect 223398 352294 223494 352350
rect 222874 352226 223494 352294
rect 222874 352170 222970 352226
rect 223026 352170 223094 352226
rect 223150 352170 223218 352226
rect 223274 352170 223342 352226
rect 223398 352170 223494 352226
rect 222874 352102 223494 352170
rect 222874 352046 222970 352102
rect 223026 352046 223094 352102
rect 223150 352046 223218 352102
rect 223274 352046 223342 352102
rect 223398 352046 223494 352102
rect 222874 351978 223494 352046
rect 222874 351922 222970 351978
rect 223026 351922 223094 351978
rect 223150 351922 223218 351978
rect 223274 351922 223342 351978
rect 223398 351922 223494 351978
rect 222874 334350 223494 351922
rect 222874 334294 222970 334350
rect 223026 334294 223094 334350
rect 223150 334294 223218 334350
rect 223274 334294 223342 334350
rect 223398 334294 223494 334350
rect 222874 334226 223494 334294
rect 222874 334170 222970 334226
rect 223026 334170 223094 334226
rect 223150 334170 223218 334226
rect 223274 334170 223342 334226
rect 223398 334170 223494 334226
rect 222874 334102 223494 334170
rect 222874 334046 222970 334102
rect 223026 334046 223094 334102
rect 223150 334046 223218 334102
rect 223274 334046 223342 334102
rect 223398 334046 223494 334102
rect 222874 333978 223494 334046
rect 222874 333922 222970 333978
rect 223026 333922 223094 333978
rect 223150 333922 223218 333978
rect 223274 333922 223342 333978
rect 223398 333922 223494 333978
rect 222874 316350 223494 333922
rect 222874 316294 222970 316350
rect 223026 316294 223094 316350
rect 223150 316294 223218 316350
rect 223274 316294 223342 316350
rect 223398 316294 223494 316350
rect 222874 316226 223494 316294
rect 222874 316170 222970 316226
rect 223026 316170 223094 316226
rect 223150 316170 223218 316226
rect 223274 316170 223342 316226
rect 223398 316170 223494 316226
rect 222874 316102 223494 316170
rect 222874 316046 222970 316102
rect 223026 316046 223094 316102
rect 223150 316046 223218 316102
rect 223274 316046 223342 316102
rect 223398 316046 223494 316102
rect 222874 315978 223494 316046
rect 222874 315922 222970 315978
rect 223026 315922 223094 315978
rect 223150 315922 223218 315978
rect 223274 315922 223342 315978
rect 223398 315922 223494 315978
rect 222874 298350 223494 315922
rect 222874 298294 222970 298350
rect 223026 298294 223094 298350
rect 223150 298294 223218 298350
rect 223274 298294 223342 298350
rect 223398 298294 223494 298350
rect 222874 298226 223494 298294
rect 222874 298170 222970 298226
rect 223026 298170 223094 298226
rect 223150 298170 223218 298226
rect 223274 298170 223342 298226
rect 223398 298170 223494 298226
rect 222874 298102 223494 298170
rect 222874 298046 222970 298102
rect 223026 298046 223094 298102
rect 223150 298046 223218 298102
rect 223274 298046 223342 298102
rect 223398 298046 223494 298102
rect 222874 297978 223494 298046
rect 222874 297922 222970 297978
rect 223026 297922 223094 297978
rect 223150 297922 223218 297978
rect 223274 297922 223342 297978
rect 223398 297922 223494 297978
rect 222874 280350 223494 297922
rect 222874 280294 222970 280350
rect 223026 280294 223094 280350
rect 223150 280294 223218 280350
rect 223274 280294 223342 280350
rect 223398 280294 223494 280350
rect 222874 280226 223494 280294
rect 222874 280170 222970 280226
rect 223026 280170 223094 280226
rect 223150 280170 223218 280226
rect 223274 280170 223342 280226
rect 223398 280170 223494 280226
rect 222874 280102 223494 280170
rect 222874 280046 222970 280102
rect 223026 280046 223094 280102
rect 223150 280046 223218 280102
rect 223274 280046 223342 280102
rect 223398 280046 223494 280102
rect 222874 279978 223494 280046
rect 222874 279922 222970 279978
rect 223026 279922 223094 279978
rect 223150 279922 223218 279978
rect 223274 279922 223342 279978
rect 223398 279922 223494 279978
rect 222874 262350 223494 279922
rect 222874 262294 222970 262350
rect 223026 262294 223094 262350
rect 223150 262294 223218 262350
rect 223274 262294 223342 262350
rect 223398 262294 223494 262350
rect 222874 262226 223494 262294
rect 222874 262170 222970 262226
rect 223026 262170 223094 262226
rect 223150 262170 223218 262226
rect 223274 262170 223342 262226
rect 223398 262170 223494 262226
rect 222874 262102 223494 262170
rect 222874 262046 222970 262102
rect 223026 262046 223094 262102
rect 223150 262046 223218 262102
rect 223274 262046 223342 262102
rect 223398 262046 223494 262102
rect 222874 261978 223494 262046
rect 222874 261922 222970 261978
rect 223026 261922 223094 261978
rect 223150 261922 223218 261978
rect 223274 261922 223342 261978
rect 223398 261922 223494 261978
rect 222874 244350 223494 261922
rect 222874 244294 222970 244350
rect 223026 244294 223094 244350
rect 223150 244294 223218 244350
rect 223274 244294 223342 244350
rect 223398 244294 223494 244350
rect 222874 244226 223494 244294
rect 222874 244170 222970 244226
rect 223026 244170 223094 244226
rect 223150 244170 223218 244226
rect 223274 244170 223342 244226
rect 223398 244170 223494 244226
rect 222874 244102 223494 244170
rect 222874 244046 222970 244102
rect 223026 244046 223094 244102
rect 223150 244046 223218 244102
rect 223274 244046 223342 244102
rect 223398 244046 223494 244102
rect 222874 243978 223494 244046
rect 222874 243922 222970 243978
rect 223026 243922 223094 243978
rect 223150 243922 223218 243978
rect 223274 243922 223342 243978
rect 223398 243922 223494 243978
rect 222874 226350 223494 243922
rect 237154 597212 237774 598268
rect 237154 597156 237250 597212
rect 237306 597156 237374 597212
rect 237430 597156 237498 597212
rect 237554 597156 237622 597212
rect 237678 597156 237774 597212
rect 237154 597088 237774 597156
rect 237154 597032 237250 597088
rect 237306 597032 237374 597088
rect 237430 597032 237498 597088
rect 237554 597032 237622 597088
rect 237678 597032 237774 597088
rect 237154 596964 237774 597032
rect 237154 596908 237250 596964
rect 237306 596908 237374 596964
rect 237430 596908 237498 596964
rect 237554 596908 237622 596964
rect 237678 596908 237774 596964
rect 237154 596840 237774 596908
rect 237154 596784 237250 596840
rect 237306 596784 237374 596840
rect 237430 596784 237498 596840
rect 237554 596784 237622 596840
rect 237678 596784 237774 596840
rect 237154 580350 237774 596784
rect 237154 580294 237250 580350
rect 237306 580294 237374 580350
rect 237430 580294 237498 580350
rect 237554 580294 237622 580350
rect 237678 580294 237774 580350
rect 237154 580226 237774 580294
rect 237154 580170 237250 580226
rect 237306 580170 237374 580226
rect 237430 580170 237498 580226
rect 237554 580170 237622 580226
rect 237678 580170 237774 580226
rect 237154 580102 237774 580170
rect 237154 580046 237250 580102
rect 237306 580046 237374 580102
rect 237430 580046 237498 580102
rect 237554 580046 237622 580102
rect 237678 580046 237774 580102
rect 237154 579978 237774 580046
rect 237154 579922 237250 579978
rect 237306 579922 237374 579978
rect 237430 579922 237498 579978
rect 237554 579922 237622 579978
rect 237678 579922 237774 579978
rect 237154 562350 237774 579922
rect 237154 562294 237250 562350
rect 237306 562294 237374 562350
rect 237430 562294 237498 562350
rect 237554 562294 237622 562350
rect 237678 562294 237774 562350
rect 237154 562226 237774 562294
rect 237154 562170 237250 562226
rect 237306 562170 237374 562226
rect 237430 562170 237498 562226
rect 237554 562170 237622 562226
rect 237678 562170 237774 562226
rect 237154 562102 237774 562170
rect 237154 562046 237250 562102
rect 237306 562046 237374 562102
rect 237430 562046 237498 562102
rect 237554 562046 237622 562102
rect 237678 562046 237774 562102
rect 237154 561978 237774 562046
rect 237154 561922 237250 561978
rect 237306 561922 237374 561978
rect 237430 561922 237498 561978
rect 237554 561922 237622 561978
rect 237678 561922 237774 561978
rect 237154 544350 237774 561922
rect 237154 544294 237250 544350
rect 237306 544294 237374 544350
rect 237430 544294 237498 544350
rect 237554 544294 237622 544350
rect 237678 544294 237774 544350
rect 237154 544226 237774 544294
rect 237154 544170 237250 544226
rect 237306 544170 237374 544226
rect 237430 544170 237498 544226
rect 237554 544170 237622 544226
rect 237678 544170 237774 544226
rect 237154 544102 237774 544170
rect 237154 544046 237250 544102
rect 237306 544046 237374 544102
rect 237430 544046 237498 544102
rect 237554 544046 237622 544102
rect 237678 544046 237774 544102
rect 237154 543978 237774 544046
rect 237154 543922 237250 543978
rect 237306 543922 237374 543978
rect 237430 543922 237498 543978
rect 237554 543922 237622 543978
rect 237678 543922 237774 543978
rect 237154 526350 237774 543922
rect 237154 526294 237250 526350
rect 237306 526294 237374 526350
rect 237430 526294 237498 526350
rect 237554 526294 237622 526350
rect 237678 526294 237774 526350
rect 237154 526226 237774 526294
rect 237154 526170 237250 526226
rect 237306 526170 237374 526226
rect 237430 526170 237498 526226
rect 237554 526170 237622 526226
rect 237678 526170 237774 526226
rect 237154 526102 237774 526170
rect 237154 526046 237250 526102
rect 237306 526046 237374 526102
rect 237430 526046 237498 526102
rect 237554 526046 237622 526102
rect 237678 526046 237774 526102
rect 237154 525978 237774 526046
rect 237154 525922 237250 525978
rect 237306 525922 237374 525978
rect 237430 525922 237498 525978
rect 237554 525922 237622 525978
rect 237678 525922 237774 525978
rect 237154 508350 237774 525922
rect 237154 508294 237250 508350
rect 237306 508294 237374 508350
rect 237430 508294 237498 508350
rect 237554 508294 237622 508350
rect 237678 508294 237774 508350
rect 237154 508226 237774 508294
rect 237154 508170 237250 508226
rect 237306 508170 237374 508226
rect 237430 508170 237498 508226
rect 237554 508170 237622 508226
rect 237678 508170 237774 508226
rect 237154 508102 237774 508170
rect 237154 508046 237250 508102
rect 237306 508046 237374 508102
rect 237430 508046 237498 508102
rect 237554 508046 237622 508102
rect 237678 508046 237774 508102
rect 237154 507978 237774 508046
rect 237154 507922 237250 507978
rect 237306 507922 237374 507978
rect 237430 507922 237498 507978
rect 237554 507922 237622 507978
rect 237678 507922 237774 507978
rect 237154 490350 237774 507922
rect 237154 490294 237250 490350
rect 237306 490294 237374 490350
rect 237430 490294 237498 490350
rect 237554 490294 237622 490350
rect 237678 490294 237774 490350
rect 237154 490226 237774 490294
rect 237154 490170 237250 490226
rect 237306 490170 237374 490226
rect 237430 490170 237498 490226
rect 237554 490170 237622 490226
rect 237678 490170 237774 490226
rect 237154 490102 237774 490170
rect 237154 490046 237250 490102
rect 237306 490046 237374 490102
rect 237430 490046 237498 490102
rect 237554 490046 237622 490102
rect 237678 490046 237774 490102
rect 237154 489978 237774 490046
rect 237154 489922 237250 489978
rect 237306 489922 237374 489978
rect 237430 489922 237498 489978
rect 237554 489922 237622 489978
rect 237678 489922 237774 489978
rect 237154 472350 237774 489922
rect 237154 472294 237250 472350
rect 237306 472294 237374 472350
rect 237430 472294 237498 472350
rect 237554 472294 237622 472350
rect 237678 472294 237774 472350
rect 237154 472226 237774 472294
rect 237154 472170 237250 472226
rect 237306 472170 237374 472226
rect 237430 472170 237498 472226
rect 237554 472170 237622 472226
rect 237678 472170 237774 472226
rect 237154 472102 237774 472170
rect 237154 472046 237250 472102
rect 237306 472046 237374 472102
rect 237430 472046 237498 472102
rect 237554 472046 237622 472102
rect 237678 472046 237774 472102
rect 237154 471978 237774 472046
rect 237154 471922 237250 471978
rect 237306 471922 237374 471978
rect 237430 471922 237498 471978
rect 237554 471922 237622 471978
rect 237678 471922 237774 471978
rect 237154 454350 237774 471922
rect 237154 454294 237250 454350
rect 237306 454294 237374 454350
rect 237430 454294 237498 454350
rect 237554 454294 237622 454350
rect 237678 454294 237774 454350
rect 237154 454226 237774 454294
rect 237154 454170 237250 454226
rect 237306 454170 237374 454226
rect 237430 454170 237498 454226
rect 237554 454170 237622 454226
rect 237678 454170 237774 454226
rect 237154 454102 237774 454170
rect 237154 454046 237250 454102
rect 237306 454046 237374 454102
rect 237430 454046 237498 454102
rect 237554 454046 237622 454102
rect 237678 454046 237774 454102
rect 237154 453978 237774 454046
rect 237154 453922 237250 453978
rect 237306 453922 237374 453978
rect 237430 453922 237498 453978
rect 237554 453922 237622 453978
rect 237678 453922 237774 453978
rect 237154 436350 237774 453922
rect 237154 436294 237250 436350
rect 237306 436294 237374 436350
rect 237430 436294 237498 436350
rect 237554 436294 237622 436350
rect 237678 436294 237774 436350
rect 237154 436226 237774 436294
rect 237154 436170 237250 436226
rect 237306 436170 237374 436226
rect 237430 436170 237498 436226
rect 237554 436170 237622 436226
rect 237678 436170 237774 436226
rect 237154 436102 237774 436170
rect 237154 436046 237250 436102
rect 237306 436046 237374 436102
rect 237430 436046 237498 436102
rect 237554 436046 237622 436102
rect 237678 436046 237774 436102
rect 237154 435978 237774 436046
rect 237154 435922 237250 435978
rect 237306 435922 237374 435978
rect 237430 435922 237498 435978
rect 237554 435922 237622 435978
rect 237678 435922 237774 435978
rect 237154 418350 237774 435922
rect 237154 418294 237250 418350
rect 237306 418294 237374 418350
rect 237430 418294 237498 418350
rect 237554 418294 237622 418350
rect 237678 418294 237774 418350
rect 237154 418226 237774 418294
rect 237154 418170 237250 418226
rect 237306 418170 237374 418226
rect 237430 418170 237498 418226
rect 237554 418170 237622 418226
rect 237678 418170 237774 418226
rect 237154 418102 237774 418170
rect 237154 418046 237250 418102
rect 237306 418046 237374 418102
rect 237430 418046 237498 418102
rect 237554 418046 237622 418102
rect 237678 418046 237774 418102
rect 237154 417978 237774 418046
rect 237154 417922 237250 417978
rect 237306 417922 237374 417978
rect 237430 417922 237498 417978
rect 237554 417922 237622 417978
rect 237678 417922 237774 417978
rect 237154 400350 237774 417922
rect 237154 400294 237250 400350
rect 237306 400294 237374 400350
rect 237430 400294 237498 400350
rect 237554 400294 237622 400350
rect 237678 400294 237774 400350
rect 237154 400226 237774 400294
rect 237154 400170 237250 400226
rect 237306 400170 237374 400226
rect 237430 400170 237498 400226
rect 237554 400170 237622 400226
rect 237678 400170 237774 400226
rect 237154 400102 237774 400170
rect 237154 400046 237250 400102
rect 237306 400046 237374 400102
rect 237430 400046 237498 400102
rect 237554 400046 237622 400102
rect 237678 400046 237774 400102
rect 237154 399978 237774 400046
rect 237154 399922 237250 399978
rect 237306 399922 237374 399978
rect 237430 399922 237498 399978
rect 237554 399922 237622 399978
rect 237678 399922 237774 399978
rect 237154 382350 237774 399922
rect 237154 382294 237250 382350
rect 237306 382294 237374 382350
rect 237430 382294 237498 382350
rect 237554 382294 237622 382350
rect 237678 382294 237774 382350
rect 237154 382226 237774 382294
rect 237154 382170 237250 382226
rect 237306 382170 237374 382226
rect 237430 382170 237498 382226
rect 237554 382170 237622 382226
rect 237678 382170 237774 382226
rect 237154 382102 237774 382170
rect 237154 382046 237250 382102
rect 237306 382046 237374 382102
rect 237430 382046 237498 382102
rect 237554 382046 237622 382102
rect 237678 382046 237774 382102
rect 237154 381978 237774 382046
rect 237154 381922 237250 381978
rect 237306 381922 237374 381978
rect 237430 381922 237498 381978
rect 237554 381922 237622 381978
rect 237678 381922 237774 381978
rect 237154 364350 237774 381922
rect 237154 364294 237250 364350
rect 237306 364294 237374 364350
rect 237430 364294 237498 364350
rect 237554 364294 237622 364350
rect 237678 364294 237774 364350
rect 237154 364226 237774 364294
rect 237154 364170 237250 364226
rect 237306 364170 237374 364226
rect 237430 364170 237498 364226
rect 237554 364170 237622 364226
rect 237678 364170 237774 364226
rect 237154 364102 237774 364170
rect 237154 364046 237250 364102
rect 237306 364046 237374 364102
rect 237430 364046 237498 364102
rect 237554 364046 237622 364102
rect 237678 364046 237774 364102
rect 237154 363978 237774 364046
rect 237154 363922 237250 363978
rect 237306 363922 237374 363978
rect 237430 363922 237498 363978
rect 237554 363922 237622 363978
rect 237678 363922 237774 363978
rect 237154 346350 237774 363922
rect 237154 346294 237250 346350
rect 237306 346294 237374 346350
rect 237430 346294 237498 346350
rect 237554 346294 237622 346350
rect 237678 346294 237774 346350
rect 237154 346226 237774 346294
rect 237154 346170 237250 346226
rect 237306 346170 237374 346226
rect 237430 346170 237498 346226
rect 237554 346170 237622 346226
rect 237678 346170 237774 346226
rect 237154 346102 237774 346170
rect 237154 346046 237250 346102
rect 237306 346046 237374 346102
rect 237430 346046 237498 346102
rect 237554 346046 237622 346102
rect 237678 346046 237774 346102
rect 237154 345978 237774 346046
rect 237154 345922 237250 345978
rect 237306 345922 237374 345978
rect 237430 345922 237498 345978
rect 237554 345922 237622 345978
rect 237678 345922 237774 345978
rect 237154 328350 237774 345922
rect 237154 328294 237250 328350
rect 237306 328294 237374 328350
rect 237430 328294 237498 328350
rect 237554 328294 237622 328350
rect 237678 328294 237774 328350
rect 237154 328226 237774 328294
rect 237154 328170 237250 328226
rect 237306 328170 237374 328226
rect 237430 328170 237498 328226
rect 237554 328170 237622 328226
rect 237678 328170 237774 328226
rect 237154 328102 237774 328170
rect 237154 328046 237250 328102
rect 237306 328046 237374 328102
rect 237430 328046 237498 328102
rect 237554 328046 237622 328102
rect 237678 328046 237774 328102
rect 237154 327978 237774 328046
rect 237154 327922 237250 327978
rect 237306 327922 237374 327978
rect 237430 327922 237498 327978
rect 237554 327922 237622 327978
rect 237678 327922 237774 327978
rect 237154 310350 237774 327922
rect 237154 310294 237250 310350
rect 237306 310294 237374 310350
rect 237430 310294 237498 310350
rect 237554 310294 237622 310350
rect 237678 310294 237774 310350
rect 237154 310226 237774 310294
rect 237154 310170 237250 310226
rect 237306 310170 237374 310226
rect 237430 310170 237498 310226
rect 237554 310170 237622 310226
rect 237678 310170 237774 310226
rect 237154 310102 237774 310170
rect 237154 310046 237250 310102
rect 237306 310046 237374 310102
rect 237430 310046 237498 310102
rect 237554 310046 237622 310102
rect 237678 310046 237774 310102
rect 237154 309978 237774 310046
rect 237154 309922 237250 309978
rect 237306 309922 237374 309978
rect 237430 309922 237498 309978
rect 237554 309922 237622 309978
rect 237678 309922 237774 309978
rect 237154 292350 237774 309922
rect 237154 292294 237250 292350
rect 237306 292294 237374 292350
rect 237430 292294 237498 292350
rect 237554 292294 237622 292350
rect 237678 292294 237774 292350
rect 237154 292226 237774 292294
rect 237154 292170 237250 292226
rect 237306 292170 237374 292226
rect 237430 292170 237498 292226
rect 237554 292170 237622 292226
rect 237678 292170 237774 292226
rect 237154 292102 237774 292170
rect 237154 292046 237250 292102
rect 237306 292046 237374 292102
rect 237430 292046 237498 292102
rect 237554 292046 237622 292102
rect 237678 292046 237774 292102
rect 237154 291978 237774 292046
rect 237154 291922 237250 291978
rect 237306 291922 237374 291978
rect 237430 291922 237498 291978
rect 237554 291922 237622 291978
rect 237678 291922 237774 291978
rect 237154 274350 237774 291922
rect 237154 274294 237250 274350
rect 237306 274294 237374 274350
rect 237430 274294 237498 274350
rect 237554 274294 237622 274350
rect 237678 274294 237774 274350
rect 237154 274226 237774 274294
rect 237154 274170 237250 274226
rect 237306 274170 237374 274226
rect 237430 274170 237498 274226
rect 237554 274170 237622 274226
rect 237678 274170 237774 274226
rect 237154 274102 237774 274170
rect 237154 274046 237250 274102
rect 237306 274046 237374 274102
rect 237430 274046 237498 274102
rect 237554 274046 237622 274102
rect 237678 274046 237774 274102
rect 237154 273978 237774 274046
rect 237154 273922 237250 273978
rect 237306 273922 237374 273978
rect 237430 273922 237498 273978
rect 237554 273922 237622 273978
rect 237678 273922 237774 273978
rect 237154 256350 237774 273922
rect 237154 256294 237250 256350
rect 237306 256294 237374 256350
rect 237430 256294 237498 256350
rect 237554 256294 237622 256350
rect 237678 256294 237774 256350
rect 237154 256226 237774 256294
rect 237154 256170 237250 256226
rect 237306 256170 237374 256226
rect 237430 256170 237498 256226
rect 237554 256170 237622 256226
rect 237678 256170 237774 256226
rect 237154 256102 237774 256170
rect 237154 256046 237250 256102
rect 237306 256046 237374 256102
rect 237430 256046 237498 256102
rect 237554 256046 237622 256102
rect 237678 256046 237774 256102
rect 237154 255978 237774 256046
rect 237154 255922 237250 255978
rect 237306 255922 237374 255978
rect 237430 255922 237498 255978
rect 237554 255922 237622 255978
rect 237678 255922 237774 255978
rect 237154 238350 237774 255922
rect 237154 238294 237250 238350
rect 237306 238294 237374 238350
rect 237430 238294 237498 238350
rect 237554 238294 237622 238350
rect 237678 238294 237774 238350
rect 237154 238226 237774 238294
rect 237154 238170 237250 238226
rect 237306 238170 237374 238226
rect 237430 238170 237498 238226
rect 237554 238170 237622 238226
rect 237678 238170 237774 238226
rect 237154 238102 237774 238170
rect 237154 238046 237250 238102
rect 237306 238046 237374 238102
rect 237430 238046 237498 238102
rect 237554 238046 237622 238102
rect 237678 238046 237774 238102
rect 237154 237978 237774 238046
rect 237154 237922 237250 237978
rect 237306 237922 237374 237978
rect 237430 237922 237498 237978
rect 237554 237922 237622 237978
rect 237678 237922 237774 237978
rect 222874 226294 222970 226350
rect 223026 226294 223094 226350
rect 223150 226294 223218 226350
rect 223274 226294 223342 226350
rect 223398 226294 223494 226350
rect 222874 226226 223494 226294
rect 222874 226170 222970 226226
rect 223026 226170 223094 226226
rect 223150 226170 223218 226226
rect 223274 226170 223342 226226
rect 223398 226170 223494 226226
rect 222874 226102 223494 226170
rect 222874 226046 222970 226102
rect 223026 226046 223094 226102
rect 223150 226046 223218 226102
rect 223274 226046 223342 226102
rect 223398 226046 223494 226102
rect 222874 225978 223494 226046
rect 222874 225922 222970 225978
rect 223026 225922 223094 225978
rect 223150 225922 223218 225978
rect 223274 225922 223342 225978
rect 223398 225922 223494 225978
rect 222874 219134 223494 225922
rect 233408 226350 233728 226384
rect 233408 226294 233478 226350
rect 233534 226294 233602 226350
rect 233658 226294 233728 226350
rect 233408 226226 233728 226294
rect 233408 226170 233478 226226
rect 233534 226170 233602 226226
rect 233658 226170 233728 226226
rect 233408 226102 233728 226170
rect 233408 226046 233478 226102
rect 233534 226046 233602 226102
rect 233658 226046 233728 226102
rect 233408 225978 233728 226046
rect 233408 225922 233478 225978
rect 233534 225922 233602 225978
rect 233658 225922 233728 225978
rect 233408 225888 233728 225922
rect 237154 220350 237774 237922
rect 237154 220294 237250 220350
rect 237306 220294 237374 220350
rect 237430 220294 237498 220350
rect 237554 220294 237622 220350
rect 237678 220294 237774 220350
rect 237154 220226 237774 220294
rect 237154 220170 237250 220226
rect 237306 220170 237374 220226
rect 237430 220170 237498 220226
rect 237554 220170 237622 220226
rect 237678 220170 237774 220226
rect 237154 220102 237774 220170
rect 237154 220046 237250 220102
rect 237306 220046 237374 220102
rect 237430 220046 237498 220102
rect 237554 220046 237622 220102
rect 237678 220046 237774 220102
rect 237154 219978 237774 220046
rect 237154 219922 237250 219978
rect 237306 219922 237374 219978
rect 237430 219922 237498 219978
rect 237554 219922 237622 219978
rect 237678 219922 237774 219978
rect 237154 219134 237774 219922
rect 240874 598172 241494 598268
rect 240874 598116 240970 598172
rect 241026 598116 241094 598172
rect 241150 598116 241218 598172
rect 241274 598116 241342 598172
rect 241398 598116 241494 598172
rect 240874 598048 241494 598116
rect 240874 597992 240970 598048
rect 241026 597992 241094 598048
rect 241150 597992 241218 598048
rect 241274 597992 241342 598048
rect 241398 597992 241494 598048
rect 240874 597924 241494 597992
rect 240874 597868 240970 597924
rect 241026 597868 241094 597924
rect 241150 597868 241218 597924
rect 241274 597868 241342 597924
rect 241398 597868 241494 597924
rect 240874 597800 241494 597868
rect 240874 597744 240970 597800
rect 241026 597744 241094 597800
rect 241150 597744 241218 597800
rect 241274 597744 241342 597800
rect 241398 597744 241494 597800
rect 240874 586350 241494 597744
rect 240874 586294 240970 586350
rect 241026 586294 241094 586350
rect 241150 586294 241218 586350
rect 241274 586294 241342 586350
rect 241398 586294 241494 586350
rect 240874 586226 241494 586294
rect 240874 586170 240970 586226
rect 241026 586170 241094 586226
rect 241150 586170 241218 586226
rect 241274 586170 241342 586226
rect 241398 586170 241494 586226
rect 240874 586102 241494 586170
rect 240874 586046 240970 586102
rect 241026 586046 241094 586102
rect 241150 586046 241218 586102
rect 241274 586046 241342 586102
rect 241398 586046 241494 586102
rect 240874 585978 241494 586046
rect 240874 585922 240970 585978
rect 241026 585922 241094 585978
rect 241150 585922 241218 585978
rect 241274 585922 241342 585978
rect 241398 585922 241494 585978
rect 240874 568350 241494 585922
rect 240874 568294 240970 568350
rect 241026 568294 241094 568350
rect 241150 568294 241218 568350
rect 241274 568294 241342 568350
rect 241398 568294 241494 568350
rect 240874 568226 241494 568294
rect 240874 568170 240970 568226
rect 241026 568170 241094 568226
rect 241150 568170 241218 568226
rect 241274 568170 241342 568226
rect 241398 568170 241494 568226
rect 240874 568102 241494 568170
rect 240874 568046 240970 568102
rect 241026 568046 241094 568102
rect 241150 568046 241218 568102
rect 241274 568046 241342 568102
rect 241398 568046 241494 568102
rect 240874 567978 241494 568046
rect 240874 567922 240970 567978
rect 241026 567922 241094 567978
rect 241150 567922 241218 567978
rect 241274 567922 241342 567978
rect 241398 567922 241494 567978
rect 240874 550350 241494 567922
rect 240874 550294 240970 550350
rect 241026 550294 241094 550350
rect 241150 550294 241218 550350
rect 241274 550294 241342 550350
rect 241398 550294 241494 550350
rect 240874 550226 241494 550294
rect 240874 550170 240970 550226
rect 241026 550170 241094 550226
rect 241150 550170 241218 550226
rect 241274 550170 241342 550226
rect 241398 550170 241494 550226
rect 240874 550102 241494 550170
rect 240874 550046 240970 550102
rect 241026 550046 241094 550102
rect 241150 550046 241218 550102
rect 241274 550046 241342 550102
rect 241398 550046 241494 550102
rect 240874 549978 241494 550046
rect 240874 549922 240970 549978
rect 241026 549922 241094 549978
rect 241150 549922 241218 549978
rect 241274 549922 241342 549978
rect 241398 549922 241494 549978
rect 240874 532350 241494 549922
rect 240874 532294 240970 532350
rect 241026 532294 241094 532350
rect 241150 532294 241218 532350
rect 241274 532294 241342 532350
rect 241398 532294 241494 532350
rect 240874 532226 241494 532294
rect 240874 532170 240970 532226
rect 241026 532170 241094 532226
rect 241150 532170 241218 532226
rect 241274 532170 241342 532226
rect 241398 532170 241494 532226
rect 240874 532102 241494 532170
rect 240874 532046 240970 532102
rect 241026 532046 241094 532102
rect 241150 532046 241218 532102
rect 241274 532046 241342 532102
rect 241398 532046 241494 532102
rect 240874 531978 241494 532046
rect 240874 531922 240970 531978
rect 241026 531922 241094 531978
rect 241150 531922 241218 531978
rect 241274 531922 241342 531978
rect 241398 531922 241494 531978
rect 240874 514350 241494 531922
rect 240874 514294 240970 514350
rect 241026 514294 241094 514350
rect 241150 514294 241218 514350
rect 241274 514294 241342 514350
rect 241398 514294 241494 514350
rect 240874 514226 241494 514294
rect 240874 514170 240970 514226
rect 241026 514170 241094 514226
rect 241150 514170 241218 514226
rect 241274 514170 241342 514226
rect 241398 514170 241494 514226
rect 240874 514102 241494 514170
rect 240874 514046 240970 514102
rect 241026 514046 241094 514102
rect 241150 514046 241218 514102
rect 241274 514046 241342 514102
rect 241398 514046 241494 514102
rect 240874 513978 241494 514046
rect 240874 513922 240970 513978
rect 241026 513922 241094 513978
rect 241150 513922 241218 513978
rect 241274 513922 241342 513978
rect 241398 513922 241494 513978
rect 240874 496350 241494 513922
rect 240874 496294 240970 496350
rect 241026 496294 241094 496350
rect 241150 496294 241218 496350
rect 241274 496294 241342 496350
rect 241398 496294 241494 496350
rect 240874 496226 241494 496294
rect 240874 496170 240970 496226
rect 241026 496170 241094 496226
rect 241150 496170 241218 496226
rect 241274 496170 241342 496226
rect 241398 496170 241494 496226
rect 240874 496102 241494 496170
rect 240874 496046 240970 496102
rect 241026 496046 241094 496102
rect 241150 496046 241218 496102
rect 241274 496046 241342 496102
rect 241398 496046 241494 496102
rect 240874 495978 241494 496046
rect 240874 495922 240970 495978
rect 241026 495922 241094 495978
rect 241150 495922 241218 495978
rect 241274 495922 241342 495978
rect 241398 495922 241494 495978
rect 240874 478350 241494 495922
rect 240874 478294 240970 478350
rect 241026 478294 241094 478350
rect 241150 478294 241218 478350
rect 241274 478294 241342 478350
rect 241398 478294 241494 478350
rect 240874 478226 241494 478294
rect 240874 478170 240970 478226
rect 241026 478170 241094 478226
rect 241150 478170 241218 478226
rect 241274 478170 241342 478226
rect 241398 478170 241494 478226
rect 240874 478102 241494 478170
rect 240874 478046 240970 478102
rect 241026 478046 241094 478102
rect 241150 478046 241218 478102
rect 241274 478046 241342 478102
rect 241398 478046 241494 478102
rect 240874 477978 241494 478046
rect 240874 477922 240970 477978
rect 241026 477922 241094 477978
rect 241150 477922 241218 477978
rect 241274 477922 241342 477978
rect 241398 477922 241494 477978
rect 240874 460350 241494 477922
rect 240874 460294 240970 460350
rect 241026 460294 241094 460350
rect 241150 460294 241218 460350
rect 241274 460294 241342 460350
rect 241398 460294 241494 460350
rect 240874 460226 241494 460294
rect 240874 460170 240970 460226
rect 241026 460170 241094 460226
rect 241150 460170 241218 460226
rect 241274 460170 241342 460226
rect 241398 460170 241494 460226
rect 240874 460102 241494 460170
rect 240874 460046 240970 460102
rect 241026 460046 241094 460102
rect 241150 460046 241218 460102
rect 241274 460046 241342 460102
rect 241398 460046 241494 460102
rect 240874 459978 241494 460046
rect 240874 459922 240970 459978
rect 241026 459922 241094 459978
rect 241150 459922 241218 459978
rect 241274 459922 241342 459978
rect 241398 459922 241494 459978
rect 240874 442350 241494 459922
rect 240874 442294 240970 442350
rect 241026 442294 241094 442350
rect 241150 442294 241218 442350
rect 241274 442294 241342 442350
rect 241398 442294 241494 442350
rect 240874 442226 241494 442294
rect 240874 442170 240970 442226
rect 241026 442170 241094 442226
rect 241150 442170 241218 442226
rect 241274 442170 241342 442226
rect 241398 442170 241494 442226
rect 240874 442102 241494 442170
rect 240874 442046 240970 442102
rect 241026 442046 241094 442102
rect 241150 442046 241218 442102
rect 241274 442046 241342 442102
rect 241398 442046 241494 442102
rect 240874 441978 241494 442046
rect 240874 441922 240970 441978
rect 241026 441922 241094 441978
rect 241150 441922 241218 441978
rect 241274 441922 241342 441978
rect 241398 441922 241494 441978
rect 240874 424350 241494 441922
rect 240874 424294 240970 424350
rect 241026 424294 241094 424350
rect 241150 424294 241218 424350
rect 241274 424294 241342 424350
rect 241398 424294 241494 424350
rect 240874 424226 241494 424294
rect 240874 424170 240970 424226
rect 241026 424170 241094 424226
rect 241150 424170 241218 424226
rect 241274 424170 241342 424226
rect 241398 424170 241494 424226
rect 240874 424102 241494 424170
rect 240874 424046 240970 424102
rect 241026 424046 241094 424102
rect 241150 424046 241218 424102
rect 241274 424046 241342 424102
rect 241398 424046 241494 424102
rect 240874 423978 241494 424046
rect 240874 423922 240970 423978
rect 241026 423922 241094 423978
rect 241150 423922 241218 423978
rect 241274 423922 241342 423978
rect 241398 423922 241494 423978
rect 240874 406350 241494 423922
rect 240874 406294 240970 406350
rect 241026 406294 241094 406350
rect 241150 406294 241218 406350
rect 241274 406294 241342 406350
rect 241398 406294 241494 406350
rect 240874 406226 241494 406294
rect 240874 406170 240970 406226
rect 241026 406170 241094 406226
rect 241150 406170 241218 406226
rect 241274 406170 241342 406226
rect 241398 406170 241494 406226
rect 240874 406102 241494 406170
rect 240874 406046 240970 406102
rect 241026 406046 241094 406102
rect 241150 406046 241218 406102
rect 241274 406046 241342 406102
rect 241398 406046 241494 406102
rect 240874 405978 241494 406046
rect 240874 405922 240970 405978
rect 241026 405922 241094 405978
rect 241150 405922 241218 405978
rect 241274 405922 241342 405978
rect 241398 405922 241494 405978
rect 240874 388350 241494 405922
rect 240874 388294 240970 388350
rect 241026 388294 241094 388350
rect 241150 388294 241218 388350
rect 241274 388294 241342 388350
rect 241398 388294 241494 388350
rect 240874 388226 241494 388294
rect 240874 388170 240970 388226
rect 241026 388170 241094 388226
rect 241150 388170 241218 388226
rect 241274 388170 241342 388226
rect 241398 388170 241494 388226
rect 240874 388102 241494 388170
rect 240874 388046 240970 388102
rect 241026 388046 241094 388102
rect 241150 388046 241218 388102
rect 241274 388046 241342 388102
rect 241398 388046 241494 388102
rect 240874 387978 241494 388046
rect 240874 387922 240970 387978
rect 241026 387922 241094 387978
rect 241150 387922 241218 387978
rect 241274 387922 241342 387978
rect 241398 387922 241494 387978
rect 240874 370350 241494 387922
rect 240874 370294 240970 370350
rect 241026 370294 241094 370350
rect 241150 370294 241218 370350
rect 241274 370294 241342 370350
rect 241398 370294 241494 370350
rect 240874 370226 241494 370294
rect 240874 370170 240970 370226
rect 241026 370170 241094 370226
rect 241150 370170 241218 370226
rect 241274 370170 241342 370226
rect 241398 370170 241494 370226
rect 240874 370102 241494 370170
rect 240874 370046 240970 370102
rect 241026 370046 241094 370102
rect 241150 370046 241218 370102
rect 241274 370046 241342 370102
rect 241398 370046 241494 370102
rect 240874 369978 241494 370046
rect 240874 369922 240970 369978
rect 241026 369922 241094 369978
rect 241150 369922 241218 369978
rect 241274 369922 241342 369978
rect 241398 369922 241494 369978
rect 240874 352350 241494 369922
rect 240874 352294 240970 352350
rect 241026 352294 241094 352350
rect 241150 352294 241218 352350
rect 241274 352294 241342 352350
rect 241398 352294 241494 352350
rect 240874 352226 241494 352294
rect 240874 352170 240970 352226
rect 241026 352170 241094 352226
rect 241150 352170 241218 352226
rect 241274 352170 241342 352226
rect 241398 352170 241494 352226
rect 240874 352102 241494 352170
rect 240874 352046 240970 352102
rect 241026 352046 241094 352102
rect 241150 352046 241218 352102
rect 241274 352046 241342 352102
rect 241398 352046 241494 352102
rect 240874 351978 241494 352046
rect 240874 351922 240970 351978
rect 241026 351922 241094 351978
rect 241150 351922 241218 351978
rect 241274 351922 241342 351978
rect 241398 351922 241494 351978
rect 240874 334350 241494 351922
rect 240874 334294 240970 334350
rect 241026 334294 241094 334350
rect 241150 334294 241218 334350
rect 241274 334294 241342 334350
rect 241398 334294 241494 334350
rect 240874 334226 241494 334294
rect 240874 334170 240970 334226
rect 241026 334170 241094 334226
rect 241150 334170 241218 334226
rect 241274 334170 241342 334226
rect 241398 334170 241494 334226
rect 240874 334102 241494 334170
rect 240874 334046 240970 334102
rect 241026 334046 241094 334102
rect 241150 334046 241218 334102
rect 241274 334046 241342 334102
rect 241398 334046 241494 334102
rect 240874 333978 241494 334046
rect 240874 333922 240970 333978
rect 241026 333922 241094 333978
rect 241150 333922 241218 333978
rect 241274 333922 241342 333978
rect 241398 333922 241494 333978
rect 240874 316350 241494 333922
rect 240874 316294 240970 316350
rect 241026 316294 241094 316350
rect 241150 316294 241218 316350
rect 241274 316294 241342 316350
rect 241398 316294 241494 316350
rect 240874 316226 241494 316294
rect 240874 316170 240970 316226
rect 241026 316170 241094 316226
rect 241150 316170 241218 316226
rect 241274 316170 241342 316226
rect 241398 316170 241494 316226
rect 240874 316102 241494 316170
rect 240874 316046 240970 316102
rect 241026 316046 241094 316102
rect 241150 316046 241218 316102
rect 241274 316046 241342 316102
rect 241398 316046 241494 316102
rect 240874 315978 241494 316046
rect 240874 315922 240970 315978
rect 241026 315922 241094 315978
rect 241150 315922 241218 315978
rect 241274 315922 241342 315978
rect 241398 315922 241494 315978
rect 240874 298350 241494 315922
rect 240874 298294 240970 298350
rect 241026 298294 241094 298350
rect 241150 298294 241218 298350
rect 241274 298294 241342 298350
rect 241398 298294 241494 298350
rect 240874 298226 241494 298294
rect 240874 298170 240970 298226
rect 241026 298170 241094 298226
rect 241150 298170 241218 298226
rect 241274 298170 241342 298226
rect 241398 298170 241494 298226
rect 240874 298102 241494 298170
rect 240874 298046 240970 298102
rect 241026 298046 241094 298102
rect 241150 298046 241218 298102
rect 241274 298046 241342 298102
rect 241398 298046 241494 298102
rect 240874 297978 241494 298046
rect 240874 297922 240970 297978
rect 241026 297922 241094 297978
rect 241150 297922 241218 297978
rect 241274 297922 241342 297978
rect 241398 297922 241494 297978
rect 240874 280350 241494 297922
rect 240874 280294 240970 280350
rect 241026 280294 241094 280350
rect 241150 280294 241218 280350
rect 241274 280294 241342 280350
rect 241398 280294 241494 280350
rect 240874 280226 241494 280294
rect 240874 280170 240970 280226
rect 241026 280170 241094 280226
rect 241150 280170 241218 280226
rect 241274 280170 241342 280226
rect 241398 280170 241494 280226
rect 240874 280102 241494 280170
rect 240874 280046 240970 280102
rect 241026 280046 241094 280102
rect 241150 280046 241218 280102
rect 241274 280046 241342 280102
rect 241398 280046 241494 280102
rect 240874 279978 241494 280046
rect 240874 279922 240970 279978
rect 241026 279922 241094 279978
rect 241150 279922 241218 279978
rect 241274 279922 241342 279978
rect 241398 279922 241494 279978
rect 240874 262350 241494 279922
rect 240874 262294 240970 262350
rect 241026 262294 241094 262350
rect 241150 262294 241218 262350
rect 241274 262294 241342 262350
rect 241398 262294 241494 262350
rect 240874 262226 241494 262294
rect 240874 262170 240970 262226
rect 241026 262170 241094 262226
rect 241150 262170 241218 262226
rect 241274 262170 241342 262226
rect 241398 262170 241494 262226
rect 240874 262102 241494 262170
rect 240874 262046 240970 262102
rect 241026 262046 241094 262102
rect 241150 262046 241218 262102
rect 241274 262046 241342 262102
rect 241398 262046 241494 262102
rect 240874 261978 241494 262046
rect 240874 261922 240970 261978
rect 241026 261922 241094 261978
rect 241150 261922 241218 261978
rect 241274 261922 241342 261978
rect 241398 261922 241494 261978
rect 240874 244350 241494 261922
rect 240874 244294 240970 244350
rect 241026 244294 241094 244350
rect 241150 244294 241218 244350
rect 241274 244294 241342 244350
rect 241398 244294 241494 244350
rect 240874 244226 241494 244294
rect 240874 244170 240970 244226
rect 241026 244170 241094 244226
rect 241150 244170 241218 244226
rect 241274 244170 241342 244226
rect 241398 244170 241494 244226
rect 240874 244102 241494 244170
rect 240874 244046 240970 244102
rect 241026 244046 241094 244102
rect 241150 244046 241218 244102
rect 241274 244046 241342 244102
rect 241398 244046 241494 244102
rect 240874 243978 241494 244046
rect 240874 243922 240970 243978
rect 241026 243922 241094 243978
rect 241150 243922 241218 243978
rect 241274 243922 241342 243978
rect 241398 243922 241494 243978
rect 240874 226350 241494 243922
rect 258874 598172 259494 598268
rect 258874 598116 258970 598172
rect 259026 598116 259094 598172
rect 259150 598116 259218 598172
rect 259274 598116 259342 598172
rect 259398 598116 259494 598172
rect 258874 598048 259494 598116
rect 258874 597992 258970 598048
rect 259026 597992 259094 598048
rect 259150 597992 259218 598048
rect 259274 597992 259342 598048
rect 259398 597992 259494 598048
rect 258874 597924 259494 597992
rect 258874 597868 258970 597924
rect 259026 597868 259094 597924
rect 259150 597868 259218 597924
rect 259274 597868 259342 597924
rect 259398 597868 259494 597924
rect 258874 597800 259494 597868
rect 258874 597744 258970 597800
rect 259026 597744 259094 597800
rect 259150 597744 259218 597800
rect 259274 597744 259342 597800
rect 259398 597744 259494 597800
rect 258874 586350 259494 597744
rect 258874 586294 258970 586350
rect 259026 586294 259094 586350
rect 259150 586294 259218 586350
rect 259274 586294 259342 586350
rect 259398 586294 259494 586350
rect 258874 586226 259494 586294
rect 258874 586170 258970 586226
rect 259026 586170 259094 586226
rect 259150 586170 259218 586226
rect 259274 586170 259342 586226
rect 259398 586170 259494 586226
rect 258874 586102 259494 586170
rect 258874 586046 258970 586102
rect 259026 586046 259094 586102
rect 259150 586046 259218 586102
rect 259274 586046 259342 586102
rect 259398 586046 259494 586102
rect 258874 585978 259494 586046
rect 258874 585922 258970 585978
rect 259026 585922 259094 585978
rect 259150 585922 259218 585978
rect 259274 585922 259342 585978
rect 259398 585922 259494 585978
rect 258874 568350 259494 585922
rect 258874 568294 258970 568350
rect 259026 568294 259094 568350
rect 259150 568294 259218 568350
rect 259274 568294 259342 568350
rect 259398 568294 259494 568350
rect 258874 568226 259494 568294
rect 258874 568170 258970 568226
rect 259026 568170 259094 568226
rect 259150 568170 259218 568226
rect 259274 568170 259342 568226
rect 259398 568170 259494 568226
rect 258874 568102 259494 568170
rect 258874 568046 258970 568102
rect 259026 568046 259094 568102
rect 259150 568046 259218 568102
rect 259274 568046 259342 568102
rect 259398 568046 259494 568102
rect 258874 567978 259494 568046
rect 258874 567922 258970 567978
rect 259026 567922 259094 567978
rect 259150 567922 259218 567978
rect 259274 567922 259342 567978
rect 259398 567922 259494 567978
rect 258874 550350 259494 567922
rect 258874 550294 258970 550350
rect 259026 550294 259094 550350
rect 259150 550294 259218 550350
rect 259274 550294 259342 550350
rect 259398 550294 259494 550350
rect 258874 550226 259494 550294
rect 258874 550170 258970 550226
rect 259026 550170 259094 550226
rect 259150 550170 259218 550226
rect 259274 550170 259342 550226
rect 259398 550170 259494 550226
rect 258874 550102 259494 550170
rect 258874 550046 258970 550102
rect 259026 550046 259094 550102
rect 259150 550046 259218 550102
rect 259274 550046 259342 550102
rect 259398 550046 259494 550102
rect 258874 549978 259494 550046
rect 258874 549922 258970 549978
rect 259026 549922 259094 549978
rect 259150 549922 259218 549978
rect 259274 549922 259342 549978
rect 259398 549922 259494 549978
rect 258874 532350 259494 549922
rect 258874 532294 258970 532350
rect 259026 532294 259094 532350
rect 259150 532294 259218 532350
rect 259274 532294 259342 532350
rect 259398 532294 259494 532350
rect 258874 532226 259494 532294
rect 258874 532170 258970 532226
rect 259026 532170 259094 532226
rect 259150 532170 259218 532226
rect 259274 532170 259342 532226
rect 259398 532170 259494 532226
rect 258874 532102 259494 532170
rect 258874 532046 258970 532102
rect 259026 532046 259094 532102
rect 259150 532046 259218 532102
rect 259274 532046 259342 532102
rect 259398 532046 259494 532102
rect 258874 531978 259494 532046
rect 258874 531922 258970 531978
rect 259026 531922 259094 531978
rect 259150 531922 259218 531978
rect 259274 531922 259342 531978
rect 259398 531922 259494 531978
rect 258874 514350 259494 531922
rect 258874 514294 258970 514350
rect 259026 514294 259094 514350
rect 259150 514294 259218 514350
rect 259274 514294 259342 514350
rect 259398 514294 259494 514350
rect 258874 514226 259494 514294
rect 258874 514170 258970 514226
rect 259026 514170 259094 514226
rect 259150 514170 259218 514226
rect 259274 514170 259342 514226
rect 259398 514170 259494 514226
rect 258874 514102 259494 514170
rect 258874 514046 258970 514102
rect 259026 514046 259094 514102
rect 259150 514046 259218 514102
rect 259274 514046 259342 514102
rect 259398 514046 259494 514102
rect 258874 513978 259494 514046
rect 258874 513922 258970 513978
rect 259026 513922 259094 513978
rect 259150 513922 259218 513978
rect 259274 513922 259342 513978
rect 259398 513922 259494 513978
rect 258874 496350 259494 513922
rect 258874 496294 258970 496350
rect 259026 496294 259094 496350
rect 259150 496294 259218 496350
rect 259274 496294 259342 496350
rect 259398 496294 259494 496350
rect 258874 496226 259494 496294
rect 258874 496170 258970 496226
rect 259026 496170 259094 496226
rect 259150 496170 259218 496226
rect 259274 496170 259342 496226
rect 259398 496170 259494 496226
rect 258874 496102 259494 496170
rect 258874 496046 258970 496102
rect 259026 496046 259094 496102
rect 259150 496046 259218 496102
rect 259274 496046 259342 496102
rect 259398 496046 259494 496102
rect 258874 495978 259494 496046
rect 258874 495922 258970 495978
rect 259026 495922 259094 495978
rect 259150 495922 259218 495978
rect 259274 495922 259342 495978
rect 259398 495922 259494 495978
rect 258874 478350 259494 495922
rect 258874 478294 258970 478350
rect 259026 478294 259094 478350
rect 259150 478294 259218 478350
rect 259274 478294 259342 478350
rect 259398 478294 259494 478350
rect 258874 478226 259494 478294
rect 258874 478170 258970 478226
rect 259026 478170 259094 478226
rect 259150 478170 259218 478226
rect 259274 478170 259342 478226
rect 259398 478170 259494 478226
rect 258874 478102 259494 478170
rect 258874 478046 258970 478102
rect 259026 478046 259094 478102
rect 259150 478046 259218 478102
rect 259274 478046 259342 478102
rect 259398 478046 259494 478102
rect 258874 477978 259494 478046
rect 258874 477922 258970 477978
rect 259026 477922 259094 477978
rect 259150 477922 259218 477978
rect 259274 477922 259342 477978
rect 259398 477922 259494 477978
rect 258874 460350 259494 477922
rect 258874 460294 258970 460350
rect 259026 460294 259094 460350
rect 259150 460294 259218 460350
rect 259274 460294 259342 460350
rect 259398 460294 259494 460350
rect 258874 460226 259494 460294
rect 258874 460170 258970 460226
rect 259026 460170 259094 460226
rect 259150 460170 259218 460226
rect 259274 460170 259342 460226
rect 259398 460170 259494 460226
rect 258874 460102 259494 460170
rect 258874 460046 258970 460102
rect 259026 460046 259094 460102
rect 259150 460046 259218 460102
rect 259274 460046 259342 460102
rect 259398 460046 259494 460102
rect 258874 459978 259494 460046
rect 258874 459922 258970 459978
rect 259026 459922 259094 459978
rect 259150 459922 259218 459978
rect 259274 459922 259342 459978
rect 259398 459922 259494 459978
rect 258874 442350 259494 459922
rect 258874 442294 258970 442350
rect 259026 442294 259094 442350
rect 259150 442294 259218 442350
rect 259274 442294 259342 442350
rect 259398 442294 259494 442350
rect 258874 442226 259494 442294
rect 258874 442170 258970 442226
rect 259026 442170 259094 442226
rect 259150 442170 259218 442226
rect 259274 442170 259342 442226
rect 259398 442170 259494 442226
rect 258874 442102 259494 442170
rect 258874 442046 258970 442102
rect 259026 442046 259094 442102
rect 259150 442046 259218 442102
rect 259274 442046 259342 442102
rect 259398 442046 259494 442102
rect 258874 441978 259494 442046
rect 258874 441922 258970 441978
rect 259026 441922 259094 441978
rect 259150 441922 259218 441978
rect 259274 441922 259342 441978
rect 259398 441922 259494 441978
rect 258874 424350 259494 441922
rect 258874 424294 258970 424350
rect 259026 424294 259094 424350
rect 259150 424294 259218 424350
rect 259274 424294 259342 424350
rect 259398 424294 259494 424350
rect 258874 424226 259494 424294
rect 258874 424170 258970 424226
rect 259026 424170 259094 424226
rect 259150 424170 259218 424226
rect 259274 424170 259342 424226
rect 259398 424170 259494 424226
rect 258874 424102 259494 424170
rect 258874 424046 258970 424102
rect 259026 424046 259094 424102
rect 259150 424046 259218 424102
rect 259274 424046 259342 424102
rect 259398 424046 259494 424102
rect 258874 423978 259494 424046
rect 258874 423922 258970 423978
rect 259026 423922 259094 423978
rect 259150 423922 259218 423978
rect 259274 423922 259342 423978
rect 259398 423922 259494 423978
rect 258874 406350 259494 423922
rect 258874 406294 258970 406350
rect 259026 406294 259094 406350
rect 259150 406294 259218 406350
rect 259274 406294 259342 406350
rect 259398 406294 259494 406350
rect 258874 406226 259494 406294
rect 258874 406170 258970 406226
rect 259026 406170 259094 406226
rect 259150 406170 259218 406226
rect 259274 406170 259342 406226
rect 259398 406170 259494 406226
rect 258874 406102 259494 406170
rect 258874 406046 258970 406102
rect 259026 406046 259094 406102
rect 259150 406046 259218 406102
rect 259274 406046 259342 406102
rect 259398 406046 259494 406102
rect 258874 405978 259494 406046
rect 258874 405922 258970 405978
rect 259026 405922 259094 405978
rect 259150 405922 259218 405978
rect 259274 405922 259342 405978
rect 259398 405922 259494 405978
rect 258874 388350 259494 405922
rect 258874 388294 258970 388350
rect 259026 388294 259094 388350
rect 259150 388294 259218 388350
rect 259274 388294 259342 388350
rect 259398 388294 259494 388350
rect 258874 388226 259494 388294
rect 258874 388170 258970 388226
rect 259026 388170 259094 388226
rect 259150 388170 259218 388226
rect 259274 388170 259342 388226
rect 259398 388170 259494 388226
rect 258874 388102 259494 388170
rect 258874 388046 258970 388102
rect 259026 388046 259094 388102
rect 259150 388046 259218 388102
rect 259274 388046 259342 388102
rect 259398 388046 259494 388102
rect 258874 387978 259494 388046
rect 258874 387922 258970 387978
rect 259026 387922 259094 387978
rect 259150 387922 259218 387978
rect 259274 387922 259342 387978
rect 259398 387922 259494 387978
rect 258874 370350 259494 387922
rect 258874 370294 258970 370350
rect 259026 370294 259094 370350
rect 259150 370294 259218 370350
rect 259274 370294 259342 370350
rect 259398 370294 259494 370350
rect 258874 370226 259494 370294
rect 258874 370170 258970 370226
rect 259026 370170 259094 370226
rect 259150 370170 259218 370226
rect 259274 370170 259342 370226
rect 259398 370170 259494 370226
rect 258874 370102 259494 370170
rect 258874 370046 258970 370102
rect 259026 370046 259094 370102
rect 259150 370046 259218 370102
rect 259274 370046 259342 370102
rect 259398 370046 259494 370102
rect 258874 369978 259494 370046
rect 258874 369922 258970 369978
rect 259026 369922 259094 369978
rect 259150 369922 259218 369978
rect 259274 369922 259342 369978
rect 259398 369922 259494 369978
rect 258874 352350 259494 369922
rect 258874 352294 258970 352350
rect 259026 352294 259094 352350
rect 259150 352294 259218 352350
rect 259274 352294 259342 352350
rect 259398 352294 259494 352350
rect 258874 352226 259494 352294
rect 258874 352170 258970 352226
rect 259026 352170 259094 352226
rect 259150 352170 259218 352226
rect 259274 352170 259342 352226
rect 259398 352170 259494 352226
rect 258874 352102 259494 352170
rect 258874 352046 258970 352102
rect 259026 352046 259094 352102
rect 259150 352046 259218 352102
rect 259274 352046 259342 352102
rect 259398 352046 259494 352102
rect 258874 351978 259494 352046
rect 258874 351922 258970 351978
rect 259026 351922 259094 351978
rect 259150 351922 259218 351978
rect 259274 351922 259342 351978
rect 259398 351922 259494 351978
rect 258874 334350 259494 351922
rect 258874 334294 258970 334350
rect 259026 334294 259094 334350
rect 259150 334294 259218 334350
rect 259274 334294 259342 334350
rect 259398 334294 259494 334350
rect 258874 334226 259494 334294
rect 258874 334170 258970 334226
rect 259026 334170 259094 334226
rect 259150 334170 259218 334226
rect 259274 334170 259342 334226
rect 259398 334170 259494 334226
rect 258874 334102 259494 334170
rect 258874 334046 258970 334102
rect 259026 334046 259094 334102
rect 259150 334046 259218 334102
rect 259274 334046 259342 334102
rect 259398 334046 259494 334102
rect 258874 333978 259494 334046
rect 258874 333922 258970 333978
rect 259026 333922 259094 333978
rect 259150 333922 259218 333978
rect 259274 333922 259342 333978
rect 259398 333922 259494 333978
rect 258874 316350 259494 333922
rect 258874 316294 258970 316350
rect 259026 316294 259094 316350
rect 259150 316294 259218 316350
rect 259274 316294 259342 316350
rect 259398 316294 259494 316350
rect 258874 316226 259494 316294
rect 258874 316170 258970 316226
rect 259026 316170 259094 316226
rect 259150 316170 259218 316226
rect 259274 316170 259342 316226
rect 259398 316170 259494 316226
rect 258874 316102 259494 316170
rect 258874 316046 258970 316102
rect 259026 316046 259094 316102
rect 259150 316046 259218 316102
rect 259274 316046 259342 316102
rect 259398 316046 259494 316102
rect 258874 315978 259494 316046
rect 258874 315922 258970 315978
rect 259026 315922 259094 315978
rect 259150 315922 259218 315978
rect 259274 315922 259342 315978
rect 259398 315922 259494 315978
rect 258874 298350 259494 315922
rect 258874 298294 258970 298350
rect 259026 298294 259094 298350
rect 259150 298294 259218 298350
rect 259274 298294 259342 298350
rect 259398 298294 259494 298350
rect 258874 298226 259494 298294
rect 258874 298170 258970 298226
rect 259026 298170 259094 298226
rect 259150 298170 259218 298226
rect 259274 298170 259342 298226
rect 259398 298170 259494 298226
rect 258874 298102 259494 298170
rect 258874 298046 258970 298102
rect 259026 298046 259094 298102
rect 259150 298046 259218 298102
rect 259274 298046 259342 298102
rect 259398 298046 259494 298102
rect 258874 297978 259494 298046
rect 258874 297922 258970 297978
rect 259026 297922 259094 297978
rect 259150 297922 259218 297978
rect 259274 297922 259342 297978
rect 259398 297922 259494 297978
rect 258874 280350 259494 297922
rect 258874 280294 258970 280350
rect 259026 280294 259094 280350
rect 259150 280294 259218 280350
rect 259274 280294 259342 280350
rect 259398 280294 259494 280350
rect 258874 280226 259494 280294
rect 258874 280170 258970 280226
rect 259026 280170 259094 280226
rect 259150 280170 259218 280226
rect 259274 280170 259342 280226
rect 259398 280170 259494 280226
rect 258874 280102 259494 280170
rect 258874 280046 258970 280102
rect 259026 280046 259094 280102
rect 259150 280046 259218 280102
rect 259274 280046 259342 280102
rect 259398 280046 259494 280102
rect 258874 279978 259494 280046
rect 258874 279922 258970 279978
rect 259026 279922 259094 279978
rect 259150 279922 259218 279978
rect 259274 279922 259342 279978
rect 259398 279922 259494 279978
rect 258874 262350 259494 279922
rect 258874 262294 258970 262350
rect 259026 262294 259094 262350
rect 259150 262294 259218 262350
rect 259274 262294 259342 262350
rect 259398 262294 259494 262350
rect 258874 262226 259494 262294
rect 258874 262170 258970 262226
rect 259026 262170 259094 262226
rect 259150 262170 259218 262226
rect 259274 262170 259342 262226
rect 259398 262170 259494 262226
rect 258874 262102 259494 262170
rect 258874 262046 258970 262102
rect 259026 262046 259094 262102
rect 259150 262046 259218 262102
rect 259274 262046 259342 262102
rect 259398 262046 259494 262102
rect 258874 261978 259494 262046
rect 258874 261922 258970 261978
rect 259026 261922 259094 261978
rect 259150 261922 259218 261978
rect 259274 261922 259342 261978
rect 259398 261922 259494 261978
rect 258874 244350 259494 261922
rect 258874 244294 258970 244350
rect 259026 244294 259094 244350
rect 259150 244294 259218 244350
rect 259274 244294 259342 244350
rect 259398 244294 259494 244350
rect 258874 244226 259494 244294
rect 258874 244170 258970 244226
rect 259026 244170 259094 244226
rect 259150 244170 259218 244226
rect 259274 244170 259342 244226
rect 259398 244170 259494 244226
rect 258874 244102 259494 244170
rect 258874 244046 258970 244102
rect 259026 244046 259094 244102
rect 259150 244046 259218 244102
rect 259274 244046 259342 244102
rect 259398 244046 259494 244102
rect 258874 243978 259494 244046
rect 258874 243922 258970 243978
rect 259026 243922 259094 243978
rect 259150 243922 259218 243978
rect 259274 243922 259342 243978
rect 259398 243922 259494 243978
rect 240874 226294 240970 226350
rect 241026 226294 241094 226350
rect 241150 226294 241218 226350
rect 241274 226294 241342 226350
rect 241398 226294 241494 226350
rect 240874 226226 241494 226294
rect 240874 226170 240970 226226
rect 241026 226170 241094 226226
rect 241150 226170 241218 226226
rect 241274 226170 241342 226226
rect 241398 226170 241494 226226
rect 240874 226102 241494 226170
rect 240874 226046 240970 226102
rect 241026 226046 241094 226102
rect 241150 226046 241218 226102
rect 241274 226046 241342 226102
rect 241398 226046 241494 226102
rect 240874 225978 241494 226046
rect 240874 225922 240970 225978
rect 241026 225922 241094 225978
rect 241150 225922 241218 225978
rect 241274 225922 241342 225978
rect 241398 225922 241494 225978
rect 79808 208350 80128 208384
rect 79808 208294 79878 208350
rect 79934 208294 80002 208350
rect 80058 208294 80128 208350
rect 79808 208226 80128 208294
rect 79808 208170 79878 208226
rect 79934 208170 80002 208226
rect 80058 208170 80128 208226
rect 79808 208102 80128 208170
rect 79808 208046 79878 208102
rect 79934 208046 80002 208102
rect 80058 208046 80128 208102
rect 79808 207978 80128 208046
rect 79808 207922 79878 207978
rect 79934 207922 80002 207978
rect 80058 207922 80128 207978
rect 79808 207888 80128 207922
rect 110528 208350 110848 208384
rect 110528 208294 110598 208350
rect 110654 208294 110722 208350
rect 110778 208294 110848 208350
rect 110528 208226 110848 208294
rect 110528 208170 110598 208226
rect 110654 208170 110722 208226
rect 110778 208170 110848 208226
rect 110528 208102 110848 208170
rect 110528 208046 110598 208102
rect 110654 208046 110722 208102
rect 110778 208046 110848 208102
rect 110528 207978 110848 208046
rect 110528 207922 110598 207978
rect 110654 207922 110722 207978
rect 110778 207922 110848 207978
rect 110528 207888 110848 207922
rect 141248 208350 141568 208384
rect 141248 208294 141318 208350
rect 141374 208294 141442 208350
rect 141498 208294 141568 208350
rect 141248 208226 141568 208294
rect 141248 208170 141318 208226
rect 141374 208170 141442 208226
rect 141498 208170 141568 208226
rect 141248 208102 141568 208170
rect 141248 208046 141318 208102
rect 141374 208046 141442 208102
rect 141498 208046 141568 208102
rect 141248 207978 141568 208046
rect 141248 207922 141318 207978
rect 141374 207922 141442 207978
rect 141498 207922 141568 207978
rect 141248 207888 141568 207922
rect 171968 208350 172288 208384
rect 171968 208294 172038 208350
rect 172094 208294 172162 208350
rect 172218 208294 172288 208350
rect 171968 208226 172288 208294
rect 171968 208170 172038 208226
rect 172094 208170 172162 208226
rect 172218 208170 172288 208226
rect 171968 208102 172288 208170
rect 171968 208046 172038 208102
rect 172094 208046 172162 208102
rect 172218 208046 172288 208102
rect 171968 207978 172288 208046
rect 171968 207922 172038 207978
rect 172094 207922 172162 207978
rect 172218 207922 172288 207978
rect 171968 207888 172288 207922
rect 202688 208350 203008 208384
rect 202688 208294 202758 208350
rect 202814 208294 202882 208350
rect 202938 208294 203008 208350
rect 202688 208226 203008 208294
rect 202688 208170 202758 208226
rect 202814 208170 202882 208226
rect 202938 208170 203008 208226
rect 202688 208102 203008 208170
rect 202688 208046 202758 208102
rect 202814 208046 202882 208102
rect 202938 208046 203008 208102
rect 202688 207978 203008 208046
rect 202688 207922 202758 207978
rect 202814 207922 202882 207978
rect 202938 207922 203008 207978
rect 202688 207888 203008 207922
rect 233408 208350 233728 208384
rect 233408 208294 233478 208350
rect 233534 208294 233602 208350
rect 233658 208294 233728 208350
rect 233408 208226 233728 208294
rect 233408 208170 233478 208226
rect 233534 208170 233602 208226
rect 233658 208170 233728 208226
rect 233408 208102 233728 208170
rect 233408 208046 233478 208102
rect 233534 208046 233602 208102
rect 233658 208046 233728 208102
rect 233408 207978 233728 208046
rect 233408 207922 233478 207978
rect 233534 207922 233602 207978
rect 233658 207922 233728 207978
rect 233408 207888 233728 207922
rect 240874 208350 241494 225922
rect 255154 238350 255774 242964
rect 255154 238294 255250 238350
rect 255306 238294 255374 238350
rect 255430 238294 255498 238350
rect 255554 238294 255622 238350
rect 255678 238294 255774 238350
rect 255154 238226 255774 238294
rect 255154 238170 255250 238226
rect 255306 238170 255374 238226
rect 255430 238170 255498 238226
rect 255554 238170 255622 238226
rect 255678 238170 255774 238226
rect 255154 238102 255774 238170
rect 255154 238046 255250 238102
rect 255306 238046 255374 238102
rect 255430 238046 255498 238102
rect 255554 238046 255622 238102
rect 255678 238046 255774 238102
rect 255154 237978 255774 238046
rect 255154 237922 255250 237978
rect 255306 237922 255374 237978
rect 255430 237922 255498 237978
rect 255554 237922 255622 237978
rect 255678 237922 255774 237978
rect 243068 220724 243124 220734
rect 243068 217812 243124 220668
rect 255154 220350 255774 237922
rect 255154 220294 255250 220350
rect 255306 220294 255374 220350
rect 255430 220294 255498 220350
rect 255554 220294 255622 220350
rect 255678 220294 255774 220350
rect 255154 220226 255774 220294
rect 255154 220170 255250 220226
rect 255306 220170 255374 220226
rect 255430 220170 255498 220226
rect 255554 220170 255622 220226
rect 255678 220170 255774 220226
rect 255154 220102 255774 220170
rect 255154 220046 255250 220102
rect 255306 220046 255374 220102
rect 255430 220046 255498 220102
rect 255554 220046 255622 220102
rect 255678 220046 255774 220102
rect 255154 219978 255774 220046
rect 255154 219922 255250 219978
rect 255306 219922 255374 219978
rect 255430 219922 255498 219978
rect 255554 219922 255622 219978
rect 255678 219922 255774 219978
rect 243068 217746 243124 217756
rect 246092 218708 246148 218718
rect 242956 212660 243012 212670
rect 240874 208294 240970 208350
rect 241026 208294 241094 208350
rect 241150 208294 241218 208350
rect 241274 208294 241342 208350
rect 241398 208294 241494 208350
rect 240874 208226 241494 208294
rect 240874 208170 240970 208226
rect 241026 208170 241094 208226
rect 241150 208170 241218 208226
rect 241274 208170 241342 208226
rect 241398 208170 241494 208226
rect 240874 208102 241494 208170
rect 240874 208046 240970 208102
rect 241026 208046 241094 208102
rect 241150 208046 241218 208102
rect 241274 208046 241342 208102
rect 241398 208046 241494 208102
rect 240874 207978 241494 208046
rect 240874 207922 240970 207978
rect 241026 207922 241094 207978
rect 241150 207922 241218 207978
rect 241274 207922 241342 207978
rect 241398 207922 241494 207978
rect 57154 202294 57250 202350
rect 57306 202294 57374 202350
rect 57430 202294 57498 202350
rect 57554 202294 57622 202350
rect 57678 202294 57774 202350
rect 57154 202226 57774 202294
rect 57154 202170 57250 202226
rect 57306 202170 57374 202226
rect 57430 202170 57498 202226
rect 57554 202170 57622 202226
rect 57678 202170 57774 202226
rect 57154 202102 57774 202170
rect 57154 202046 57250 202102
rect 57306 202046 57374 202102
rect 57430 202046 57498 202102
rect 57554 202046 57622 202102
rect 57678 202046 57774 202102
rect 57154 201978 57774 202046
rect 57154 201922 57250 201978
rect 57306 201922 57374 201978
rect 57430 201922 57498 201978
rect 57554 201922 57622 201978
rect 57678 201922 57774 201978
rect 57154 184350 57774 201922
rect 64448 202350 64768 202384
rect 64448 202294 64518 202350
rect 64574 202294 64642 202350
rect 64698 202294 64768 202350
rect 64448 202226 64768 202294
rect 64448 202170 64518 202226
rect 64574 202170 64642 202226
rect 64698 202170 64768 202226
rect 64448 202102 64768 202170
rect 64448 202046 64518 202102
rect 64574 202046 64642 202102
rect 64698 202046 64768 202102
rect 64448 201978 64768 202046
rect 64448 201922 64518 201978
rect 64574 201922 64642 201978
rect 64698 201922 64768 201978
rect 64448 201888 64768 201922
rect 95168 202350 95488 202384
rect 95168 202294 95238 202350
rect 95294 202294 95362 202350
rect 95418 202294 95488 202350
rect 95168 202226 95488 202294
rect 95168 202170 95238 202226
rect 95294 202170 95362 202226
rect 95418 202170 95488 202226
rect 95168 202102 95488 202170
rect 95168 202046 95238 202102
rect 95294 202046 95362 202102
rect 95418 202046 95488 202102
rect 95168 201978 95488 202046
rect 95168 201922 95238 201978
rect 95294 201922 95362 201978
rect 95418 201922 95488 201978
rect 95168 201888 95488 201922
rect 125888 202350 126208 202384
rect 125888 202294 125958 202350
rect 126014 202294 126082 202350
rect 126138 202294 126208 202350
rect 125888 202226 126208 202294
rect 125888 202170 125958 202226
rect 126014 202170 126082 202226
rect 126138 202170 126208 202226
rect 125888 202102 126208 202170
rect 125888 202046 125958 202102
rect 126014 202046 126082 202102
rect 126138 202046 126208 202102
rect 125888 201978 126208 202046
rect 125888 201922 125958 201978
rect 126014 201922 126082 201978
rect 126138 201922 126208 201978
rect 125888 201888 126208 201922
rect 156608 202350 156928 202384
rect 156608 202294 156678 202350
rect 156734 202294 156802 202350
rect 156858 202294 156928 202350
rect 156608 202226 156928 202294
rect 156608 202170 156678 202226
rect 156734 202170 156802 202226
rect 156858 202170 156928 202226
rect 156608 202102 156928 202170
rect 156608 202046 156678 202102
rect 156734 202046 156802 202102
rect 156858 202046 156928 202102
rect 156608 201978 156928 202046
rect 156608 201922 156678 201978
rect 156734 201922 156802 201978
rect 156858 201922 156928 201978
rect 156608 201888 156928 201922
rect 187328 202350 187648 202384
rect 187328 202294 187398 202350
rect 187454 202294 187522 202350
rect 187578 202294 187648 202350
rect 187328 202226 187648 202294
rect 187328 202170 187398 202226
rect 187454 202170 187522 202226
rect 187578 202170 187648 202226
rect 187328 202102 187648 202170
rect 187328 202046 187398 202102
rect 187454 202046 187522 202102
rect 187578 202046 187648 202102
rect 187328 201978 187648 202046
rect 187328 201922 187398 201978
rect 187454 201922 187522 201978
rect 187578 201922 187648 201978
rect 187328 201888 187648 201922
rect 218048 202350 218368 202384
rect 218048 202294 218118 202350
rect 218174 202294 218242 202350
rect 218298 202294 218368 202350
rect 218048 202226 218368 202294
rect 218048 202170 218118 202226
rect 218174 202170 218242 202226
rect 218298 202170 218368 202226
rect 218048 202102 218368 202170
rect 218048 202046 218118 202102
rect 218174 202046 218242 202102
rect 218298 202046 218368 202102
rect 218048 201978 218368 202046
rect 218048 201922 218118 201978
rect 218174 201922 218242 201978
rect 218298 201922 218368 201978
rect 218048 201888 218368 201922
rect 240874 190350 241494 207922
rect 240874 190294 240970 190350
rect 241026 190294 241094 190350
rect 241150 190294 241218 190350
rect 241274 190294 241342 190350
rect 241398 190294 241494 190350
rect 240874 190226 241494 190294
rect 240874 190170 240970 190226
rect 241026 190170 241094 190226
rect 241150 190170 241218 190226
rect 241274 190170 241342 190226
rect 241398 190170 241494 190226
rect 240874 190102 241494 190170
rect 240874 190046 240970 190102
rect 241026 190046 241094 190102
rect 241150 190046 241218 190102
rect 241274 190046 241342 190102
rect 241398 190046 241494 190102
rect 240874 189978 241494 190046
rect 240874 189922 240970 189978
rect 241026 189922 241094 189978
rect 241150 189922 241218 189978
rect 241274 189922 241342 189978
rect 241398 189922 241494 189978
rect 57154 184294 57250 184350
rect 57306 184294 57374 184350
rect 57430 184294 57498 184350
rect 57554 184294 57622 184350
rect 57678 184294 57774 184350
rect 57154 184226 57774 184294
rect 57154 184170 57250 184226
rect 57306 184170 57374 184226
rect 57430 184170 57498 184226
rect 57554 184170 57622 184226
rect 57678 184170 57774 184226
rect 57154 184102 57774 184170
rect 57154 184046 57250 184102
rect 57306 184046 57374 184102
rect 57430 184046 57498 184102
rect 57554 184046 57622 184102
rect 57678 184046 57774 184102
rect 57154 183978 57774 184046
rect 57154 183922 57250 183978
rect 57306 183922 57374 183978
rect 57430 183922 57498 183978
rect 57554 183922 57622 183978
rect 57678 183922 57774 183978
rect 57154 166350 57774 183922
rect 64448 184350 64768 184384
rect 64448 184294 64518 184350
rect 64574 184294 64642 184350
rect 64698 184294 64768 184350
rect 64448 184226 64768 184294
rect 64448 184170 64518 184226
rect 64574 184170 64642 184226
rect 64698 184170 64768 184226
rect 64448 184102 64768 184170
rect 64448 184046 64518 184102
rect 64574 184046 64642 184102
rect 64698 184046 64768 184102
rect 64448 183978 64768 184046
rect 64448 183922 64518 183978
rect 64574 183922 64642 183978
rect 64698 183922 64768 183978
rect 64448 183888 64768 183922
rect 240874 172350 241494 189922
rect 242732 208628 242788 208638
rect 240874 172294 240970 172350
rect 241026 172294 241094 172350
rect 241150 172294 241218 172350
rect 241274 172294 241342 172350
rect 241398 172294 241494 172350
rect 240874 172226 241494 172294
rect 240874 172170 240970 172226
rect 241026 172170 241094 172226
rect 241150 172170 241218 172226
rect 241274 172170 241342 172226
rect 241398 172170 241494 172226
rect 240874 172102 241494 172170
rect 240874 172046 240970 172102
rect 241026 172046 241094 172102
rect 241150 172046 241218 172102
rect 241274 172046 241342 172102
rect 241398 172046 241494 172102
rect 240874 171978 241494 172046
rect 240874 171922 240970 171978
rect 241026 171922 241094 171978
rect 241150 171922 241218 171978
rect 241274 171922 241342 171978
rect 241398 171922 241494 171978
rect 57154 166294 57250 166350
rect 57306 166294 57374 166350
rect 57430 166294 57498 166350
rect 57554 166294 57622 166350
rect 57678 166294 57774 166350
rect 57154 166226 57774 166294
rect 57154 166170 57250 166226
rect 57306 166170 57374 166226
rect 57430 166170 57498 166226
rect 57554 166170 57622 166226
rect 57678 166170 57774 166226
rect 57154 166102 57774 166170
rect 57154 166046 57250 166102
rect 57306 166046 57374 166102
rect 57430 166046 57498 166102
rect 57554 166046 57622 166102
rect 57678 166046 57774 166102
rect 57154 165978 57774 166046
rect 57154 165922 57250 165978
rect 57306 165922 57374 165978
rect 57430 165922 57498 165978
rect 57554 165922 57622 165978
rect 57678 165922 57774 165978
rect 55468 150388 55524 150398
rect 55468 149044 55524 150332
rect 55468 148978 55524 148988
rect 57154 148350 57774 165922
rect 64448 166350 64768 166384
rect 64448 166294 64518 166350
rect 64574 166294 64642 166350
rect 64698 166294 64768 166350
rect 64448 166226 64768 166294
rect 64448 166170 64518 166226
rect 64574 166170 64642 166226
rect 64698 166170 64768 166226
rect 64448 166102 64768 166170
rect 64448 166046 64518 166102
rect 64574 166046 64642 166102
rect 64698 166046 64768 166102
rect 64448 165978 64768 166046
rect 64448 165922 64518 165978
rect 64574 165922 64642 165978
rect 64698 165922 64768 165978
rect 64448 165888 64768 165922
rect 240874 154350 241494 171922
rect 241948 172340 242004 172350
rect 241948 170548 242004 172284
rect 241948 170482 242004 170492
rect 242732 158564 242788 208572
rect 242732 158498 242788 158508
rect 242844 204596 242900 204606
rect 242844 156324 242900 204540
rect 242956 175588 243012 212604
rect 243068 206612 243124 206622
rect 243068 185668 243124 206556
rect 244412 205828 244468 205838
rect 243180 202580 243236 202590
rect 243180 189028 243236 202524
rect 243180 188962 243236 188972
rect 243068 185602 243124 185612
rect 242956 175522 243012 175532
rect 242844 156258 242900 156268
rect 240874 154294 240970 154350
rect 241026 154294 241094 154350
rect 241150 154294 241218 154350
rect 241274 154294 241342 154350
rect 241398 154294 241494 154350
rect 240874 154226 241494 154294
rect 240874 154170 240970 154226
rect 241026 154170 241094 154226
rect 241150 154170 241218 154226
rect 241274 154170 241342 154226
rect 241398 154170 241494 154226
rect 240874 154102 241494 154170
rect 240874 154046 240970 154102
rect 241026 154046 241094 154102
rect 241150 154046 241218 154102
rect 241274 154046 241342 154102
rect 241398 154046 241494 154102
rect 240874 153978 241494 154046
rect 240874 153922 240970 153978
rect 241026 153922 241094 153978
rect 241150 153922 241218 153978
rect 241274 153922 241342 153978
rect 241398 153922 241494 153978
rect 57154 148294 57250 148350
rect 57306 148294 57374 148350
rect 57430 148294 57498 148350
rect 57554 148294 57622 148350
rect 57678 148294 57774 148350
rect 57154 148226 57774 148294
rect 57154 148170 57250 148226
rect 57306 148170 57374 148226
rect 57430 148170 57498 148226
rect 57554 148170 57622 148226
rect 57678 148170 57774 148226
rect 57154 148102 57774 148170
rect 57154 148046 57250 148102
rect 57306 148046 57374 148102
rect 57430 148046 57498 148102
rect 57554 148046 57622 148102
rect 57678 148046 57774 148102
rect 57154 147978 57774 148046
rect 57154 147922 57250 147978
rect 57306 147922 57374 147978
rect 57430 147922 57498 147978
rect 57554 147922 57622 147978
rect 57678 147922 57774 147978
rect 57036 131908 57092 131918
rect 57036 130004 57092 131852
rect 57036 129938 57092 129948
rect 57154 130350 57774 147922
rect 64448 148350 64768 148384
rect 64448 148294 64518 148350
rect 64574 148294 64642 148350
rect 64698 148294 64768 148350
rect 64448 148226 64768 148294
rect 64448 148170 64518 148226
rect 64574 148170 64642 148226
rect 64698 148170 64768 148226
rect 64448 148102 64768 148170
rect 64448 148046 64518 148102
rect 64574 148046 64642 148102
rect 64698 148046 64768 148102
rect 64448 147978 64768 148046
rect 64448 147922 64518 147978
rect 64574 147922 64642 147978
rect 64698 147922 64768 147978
rect 64448 147888 64768 147922
rect 240874 136350 241494 153922
rect 241948 154196 242004 154206
rect 241948 150388 242004 154140
rect 241948 150322 242004 150332
rect 243068 150164 243124 150174
rect 240874 136294 240970 136350
rect 241026 136294 241094 136350
rect 241150 136294 241218 136350
rect 241274 136294 241342 136350
rect 241398 136294 241494 136350
rect 240874 136226 241494 136294
rect 240874 136170 240970 136226
rect 241026 136170 241094 136226
rect 241150 136170 241218 136226
rect 241274 136170 241342 136226
rect 241398 136170 241494 136226
rect 240874 136102 241494 136170
rect 240874 136046 240970 136102
rect 241026 136046 241094 136102
rect 241150 136046 241218 136102
rect 241274 136046 241342 136102
rect 241398 136046 241494 136102
rect 240874 135978 241494 136046
rect 240874 135922 240970 135978
rect 241026 135922 241094 135978
rect 241150 135922 241218 135978
rect 241274 135922 241342 135978
rect 241398 135922 241494 135978
rect 57154 130294 57250 130350
rect 57306 130294 57374 130350
rect 57430 130294 57498 130350
rect 57554 130294 57622 130350
rect 57678 130294 57774 130350
rect 57154 130226 57774 130294
rect 57154 130170 57250 130226
rect 57306 130170 57374 130226
rect 57430 130170 57498 130226
rect 57554 130170 57622 130226
rect 57678 130170 57774 130226
rect 57154 130102 57774 130170
rect 57154 130046 57250 130102
rect 57306 130046 57374 130102
rect 57430 130046 57498 130102
rect 57554 130046 57622 130102
rect 57678 130046 57774 130102
rect 57154 129978 57774 130046
rect 57154 129922 57250 129978
rect 57306 129922 57374 129978
rect 57430 129922 57498 129978
rect 57554 129922 57622 129978
rect 57678 129922 57774 129978
rect 57036 120148 57092 120158
rect 57036 118580 57092 120092
rect 57036 118514 57092 118524
rect 57036 113428 57092 113438
rect 57036 110964 57092 113372
rect 57036 110898 57092 110908
rect 57154 112350 57774 129922
rect 64448 130350 64768 130384
rect 64448 130294 64518 130350
rect 64574 130294 64642 130350
rect 64698 130294 64768 130350
rect 64448 130226 64768 130294
rect 64448 130170 64518 130226
rect 64574 130170 64642 130226
rect 64698 130170 64768 130226
rect 64448 130102 64768 130170
rect 64448 130046 64518 130102
rect 64574 130046 64642 130102
rect 64698 130046 64768 130102
rect 64448 129978 64768 130046
rect 64448 129922 64518 129978
rect 64574 129922 64642 129978
rect 64698 129922 64768 129978
rect 64448 129888 64768 129922
rect 240874 118350 241494 135922
rect 242732 148148 242788 148158
rect 242732 124964 242788 148092
rect 242732 124898 242788 124908
rect 242844 146132 242900 146142
rect 242844 123844 242900 146076
rect 243068 145348 243124 150108
rect 243068 145282 243124 145292
rect 243068 144116 243124 144126
rect 242844 123778 242900 123788
rect 242956 142100 243012 142110
rect 240874 118294 240970 118350
rect 241026 118294 241094 118350
rect 241150 118294 241218 118350
rect 241274 118294 241342 118350
rect 241398 118294 241494 118350
rect 240874 118226 241494 118294
rect 240874 118170 240970 118226
rect 241026 118170 241094 118226
rect 241150 118170 241218 118226
rect 241274 118170 241342 118226
rect 241398 118170 241494 118226
rect 240874 118102 241494 118170
rect 240874 118046 240970 118102
rect 241026 118046 241094 118102
rect 241150 118046 241218 118102
rect 241274 118046 241342 118102
rect 241398 118046 241494 118102
rect 240874 117978 241494 118046
rect 240874 117922 240970 117978
rect 241026 117922 241094 117978
rect 241150 117922 241218 117978
rect 241274 117922 241342 117978
rect 241398 117922 241494 117978
rect 57154 112294 57250 112350
rect 57306 112294 57374 112350
rect 57430 112294 57498 112350
rect 57554 112294 57622 112350
rect 57678 112294 57774 112350
rect 57154 112226 57774 112294
rect 57154 112170 57250 112226
rect 57306 112170 57374 112226
rect 57430 112170 57498 112226
rect 57554 112170 57622 112226
rect 57678 112170 57774 112226
rect 57154 112102 57774 112170
rect 57154 112046 57250 112102
rect 57306 112046 57374 112102
rect 57430 112046 57498 112102
rect 57554 112046 57622 112102
rect 57678 112046 57774 112102
rect 57154 111978 57774 112046
rect 57154 111922 57250 111978
rect 57306 111922 57374 111978
rect 57430 111922 57498 111978
rect 57554 111922 57622 111978
rect 57678 111922 57774 111978
rect 57036 101668 57092 101678
rect 57036 99540 57092 101612
rect 57036 99474 57092 99484
rect 44492 96562 44548 96572
rect 57036 96628 57092 96638
rect 57036 95732 57092 96572
rect 57036 95666 57092 95676
rect 57154 94350 57774 111922
rect 64448 112350 64768 112384
rect 64448 112294 64518 112350
rect 64574 112294 64642 112350
rect 64698 112294 64768 112350
rect 64448 112226 64768 112294
rect 64448 112170 64518 112226
rect 64574 112170 64642 112226
rect 64698 112170 64768 112226
rect 64448 112102 64768 112170
rect 64448 112046 64518 112102
rect 64574 112046 64642 112102
rect 64698 112046 64768 112102
rect 64448 111978 64768 112046
rect 64448 111922 64518 111978
rect 64574 111922 64642 111978
rect 64698 111922 64768 111978
rect 64448 111888 64768 111922
rect 240874 100350 241494 117922
rect 242732 121940 242788 121950
rect 242172 113876 242228 113886
rect 242060 111860 242116 111870
rect 241948 107828 242004 107838
rect 241948 102564 242004 107772
rect 242060 104804 242116 111804
rect 242172 105924 242228 113820
rect 242732 110404 242788 121884
rect 242956 121604 243012 142044
rect 243068 122724 243124 144060
rect 243068 122658 243124 122668
rect 243180 140084 243236 140094
rect 242956 121538 243012 121548
rect 243180 120484 243236 140028
rect 243404 138068 243460 138078
rect 243180 120418 243236 120428
rect 243292 125972 243348 125982
rect 242732 110338 242788 110348
rect 242956 119924 243012 119934
rect 242172 105858 242228 105868
rect 242284 109844 242340 109854
rect 242060 104738 242116 104748
rect 242284 103684 242340 109788
rect 242956 109284 243012 119868
rect 242956 109218 243012 109228
rect 243068 117908 243124 117918
rect 243068 108164 243124 117852
rect 243292 112644 243348 125916
rect 243404 119364 243460 138012
rect 243404 119298 243460 119308
rect 243292 112578 243348 112588
rect 243516 115892 243572 115902
rect 243068 108098 243124 108108
rect 243516 107044 243572 115836
rect 243516 106978 243572 106988
rect 242284 103618 242340 103628
rect 243068 105812 243124 105822
rect 241948 102498 242004 102508
rect 243068 101444 243124 105756
rect 243628 103796 243684 103806
rect 243628 101668 243684 103740
rect 243628 101602 243684 101612
rect 243068 101378 243124 101388
rect 240874 100294 240970 100350
rect 241026 100294 241094 100350
rect 241150 100294 241218 100350
rect 241274 100294 241342 100350
rect 241398 100294 241494 100350
rect 240874 100226 241494 100294
rect 240874 100170 240970 100226
rect 241026 100170 241094 100226
rect 241150 100170 241218 100226
rect 241274 100170 241342 100226
rect 241398 100170 241494 100226
rect 240874 100102 241494 100170
rect 240874 100046 240970 100102
rect 241026 100046 241094 100102
rect 241150 100046 241218 100102
rect 241274 100046 241342 100102
rect 241398 100046 241494 100102
rect 240874 99978 241494 100046
rect 240874 99922 240970 99978
rect 241026 99922 241094 99978
rect 241150 99922 241218 99978
rect 241274 99922 241342 99978
rect 241398 99922 241494 99978
rect 57154 94294 57250 94350
rect 57306 94294 57374 94350
rect 57430 94294 57498 94350
rect 57554 94294 57622 94350
rect 57678 94294 57774 94350
rect 57154 94226 57774 94294
rect 57154 94170 57250 94226
rect 57306 94170 57374 94226
rect 57430 94170 57498 94226
rect 57554 94170 57622 94226
rect 57678 94170 57774 94226
rect 57154 94102 57774 94170
rect 57154 94046 57250 94102
rect 57306 94046 57374 94102
rect 57430 94046 57498 94102
rect 57554 94046 57622 94102
rect 57678 94046 57774 94102
rect 57154 93978 57774 94046
rect 57154 93922 57250 93978
rect 57306 93922 57374 93978
rect 57430 93922 57498 93978
rect 57554 93922 57622 93978
rect 57678 93922 57774 93978
rect 57036 89908 57092 89918
rect 42874 82294 42970 82350
rect 43026 82294 43094 82350
rect 43150 82294 43218 82350
rect 43274 82294 43342 82350
rect 43398 82294 43494 82350
rect 42874 82226 43494 82294
rect 42874 82170 42970 82226
rect 43026 82170 43094 82226
rect 43150 82170 43218 82226
rect 43274 82170 43342 82226
rect 43398 82170 43494 82226
rect 42874 82102 43494 82170
rect 42874 82046 42970 82102
rect 43026 82046 43094 82102
rect 43150 82046 43218 82102
rect 43274 82046 43342 82102
rect 43398 82046 43494 82102
rect 42874 81978 43494 82046
rect 42874 81922 42970 81978
rect 43026 81922 43094 81978
rect 43150 81922 43218 81978
rect 43274 81922 43342 81978
rect 43398 81922 43494 81978
rect 42874 64350 43494 81922
rect 56252 84868 56308 84878
rect 56252 76692 56308 84812
rect 57036 84308 57092 89852
rect 57036 84242 57092 84252
rect 56252 76626 56308 76636
rect 57154 76350 57774 93922
rect 64448 94350 64768 94384
rect 64448 94294 64518 94350
rect 64574 94294 64642 94350
rect 64698 94294 64768 94350
rect 64448 94226 64768 94294
rect 64448 94170 64518 94226
rect 64574 94170 64642 94226
rect 64698 94170 64768 94226
rect 64448 94102 64768 94170
rect 64448 94046 64518 94102
rect 64574 94046 64642 94102
rect 64698 94046 64768 94102
rect 64448 93978 64768 94046
rect 64448 93922 64518 93978
rect 64574 93922 64642 93978
rect 64698 93922 64768 93978
rect 64448 93888 64768 93922
rect 240874 82350 241494 99922
rect 241948 99764 242004 99774
rect 241948 98084 242004 99708
rect 241948 98018 242004 98028
rect 241948 93604 242004 93614
rect 241948 91700 242004 93548
rect 241948 91634 242004 91644
rect 243180 92484 243236 92494
rect 243068 91364 243124 91374
rect 242060 90244 242116 90254
rect 241948 89124 242004 89134
rect 241948 83636 242004 89068
rect 242060 85652 242116 90188
rect 242060 85586 242116 85596
rect 242172 88004 242228 88014
rect 241948 83570 242004 83580
rect 240874 82294 240970 82350
rect 241026 82294 241094 82350
rect 241150 82294 241218 82350
rect 241274 82294 241342 82350
rect 241398 82294 241494 82350
rect 240874 82226 241494 82294
rect 240874 82170 240970 82226
rect 241026 82170 241094 82226
rect 241150 82170 241218 82226
rect 241274 82170 241342 82226
rect 241398 82170 241494 82226
rect 240874 82102 241494 82170
rect 240874 82046 240970 82102
rect 241026 82046 241094 82102
rect 241150 82046 241218 82102
rect 241274 82046 241342 82102
rect 241398 82046 241494 82102
rect 240874 81978 241494 82046
rect 240874 81922 240970 81978
rect 241026 81922 241094 81978
rect 241150 81922 241218 81978
rect 241274 81922 241342 81978
rect 241398 81922 241494 81978
rect 57154 76294 57250 76350
rect 57306 76294 57374 76350
rect 57430 76294 57498 76350
rect 57554 76294 57622 76350
rect 57678 76294 57774 76350
rect 57154 76226 57774 76294
rect 57154 76170 57250 76226
rect 57306 76170 57374 76226
rect 57430 76170 57498 76226
rect 57554 76170 57622 76226
rect 57678 76170 57774 76226
rect 57154 76102 57774 76170
rect 57154 76046 57250 76102
rect 57306 76046 57374 76102
rect 57430 76046 57498 76102
rect 57554 76046 57622 76102
rect 57678 76046 57774 76102
rect 57154 75978 57774 76046
rect 57154 75922 57250 75978
rect 57306 75922 57374 75978
rect 57430 75922 57498 75978
rect 57554 75922 57622 75978
rect 57678 75922 57774 75978
rect 55468 68068 55524 68078
rect 55468 65268 55524 68012
rect 55468 65202 55524 65212
rect 42874 64294 42970 64350
rect 43026 64294 43094 64350
rect 43150 64294 43218 64350
rect 43274 64294 43342 64350
rect 43398 64294 43494 64350
rect 42874 64226 43494 64294
rect 42874 64170 42970 64226
rect 43026 64170 43094 64226
rect 43150 64170 43218 64226
rect 43274 64170 43342 64226
rect 43398 64170 43494 64226
rect 42874 64102 43494 64170
rect 42874 64046 42970 64102
rect 43026 64046 43094 64102
rect 43150 64046 43218 64102
rect 43274 64046 43342 64102
rect 43398 64046 43494 64102
rect 42874 63978 43494 64046
rect 42874 63922 42970 63978
rect 43026 63922 43094 63978
rect 43150 63922 43218 63978
rect 43274 63922 43342 63978
rect 43398 63922 43494 63978
rect 42874 46350 43494 63922
rect 57036 59668 57092 59678
rect 57036 57652 57092 59612
rect 57036 57586 57092 57596
rect 57154 58350 57774 75922
rect 64448 76350 64768 76384
rect 64448 76294 64518 76350
rect 64574 76294 64642 76350
rect 64698 76294 64768 76350
rect 64448 76226 64768 76294
rect 64448 76170 64518 76226
rect 64574 76170 64642 76226
rect 64698 76170 64768 76226
rect 64448 76102 64768 76170
rect 64448 76046 64518 76102
rect 64574 76046 64642 76102
rect 64698 76046 64768 76102
rect 64448 75978 64768 76046
rect 64448 75922 64518 75978
rect 64574 75922 64642 75978
rect 64698 75922 64768 75978
rect 64448 75888 64768 75922
rect 240874 64350 241494 81922
rect 242172 81620 242228 87948
rect 243068 87668 243124 91308
rect 243180 89684 243236 92428
rect 243180 89618 243236 89628
rect 243068 87602 243124 87612
rect 242172 81554 242228 81564
rect 242284 86884 242340 86894
rect 242284 79604 242340 86828
rect 242284 79538 242340 79548
rect 242732 85764 242788 85774
rect 242732 77588 242788 85708
rect 243180 82404 243236 82414
rect 243068 80164 243124 80174
rect 242732 77522 242788 77532
rect 242844 79044 242900 79054
rect 240874 64294 240970 64350
rect 241026 64294 241094 64350
rect 241150 64294 241218 64350
rect 241274 64294 241342 64350
rect 241398 64294 241494 64350
rect 240874 64226 241494 64294
rect 240874 64170 240970 64226
rect 241026 64170 241094 64226
rect 241150 64170 241218 64226
rect 241274 64170 241342 64226
rect 241398 64170 241494 64226
rect 240874 64102 241494 64170
rect 240874 64046 240970 64102
rect 241026 64046 241094 64102
rect 241150 64046 241218 64102
rect 241274 64046 241342 64102
rect 241398 64046 241494 64102
rect 240874 63978 241494 64046
rect 240874 63922 240970 63978
rect 241026 63922 241094 63978
rect 241150 63922 241218 63978
rect 241274 63922 241342 63978
rect 241398 63922 241494 63978
rect 57154 58294 57250 58350
rect 57306 58294 57374 58350
rect 57430 58294 57498 58350
rect 57554 58294 57622 58350
rect 57678 58294 57774 58350
rect 57154 58226 57774 58294
rect 57154 58170 57250 58226
rect 57306 58170 57374 58226
rect 57430 58170 57498 58226
rect 57554 58170 57622 58226
rect 57678 58170 57774 58226
rect 57154 58102 57774 58170
rect 57154 58046 57250 58102
rect 57306 58046 57374 58102
rect 57430 58046 57498 58102
rect 57554 58046 57622 58102
rect 57678 58046 57774 58102
rect 57154 57978 57774 58046
rect 57154 57922 57250 57978
rect 57306 57922 57374 57978
rect 57430 57922 57498 57978
rect 57554 57922 57622 57978
rect 57678 57922 57774 57978
rect 42874 46294 42970 46350
rect 43026 46294 43094 46350
rect 43150 46294 43218 46350
rect 43274 46294 43342 46350
rect 43398 46294 43494 46350
rect 42874 46226 43494 46294
rect 42874 46170 42970 46226
rect 43026 46170 43094 46226
rect 43150 46170 43218 46226
rect 43274 46170 43342 46226
rect 43398 46170 43494 46226
rect 42874 46102 43494 46170
rect 57036 47908 57092 47918
rect 57036 46228 57092 47852
rect 57036 46162 57092 46172
rect 42874 46046 42970 46102
rect 43026 46046 43094 46102
rect 43150 46046 43218 46102
rect 43274 46046 43342 46102
rect 43398 46046 43494 46102
rect 42874 45978 43494 46046
rect 42874 45922 42970 45978
rect 43026 45922 43094 45978
rect 43150 45922 43218 45978
rect 43274 45922 43342 45978
rect 43398 45922 43494 45978
rect 42874 28350 43494 45922
rect 42874 28294 42970 28350
rect 43026 28294 43094 28350
rect 43150 28294 43218 28350
rect 43274 28294 43342 28350
rect 43398 28294 43494 28350
rect 42874 28226 43494 28294
rect 42874 28170 42970 28226
rect 43026 28170 43094 28226
rect 43150 28170 43218 28226
rect 43274 28170 43342 28226
rect 43398 28170 43494 28226
rect 42874 28102 43494 28170
rect 42874 28046 42970 28102
rect 43026 28046 43094 28102
rect 43150 28046 43218 28102
rect 43274 28046 43342 28102
rect 43398 28046 43494 28102
rect 42874 27978 43494 28046
rect 42874 27922 42970 27978
rect 43026 27922 43094 27978
rect 43150 27922 43218 27978
rect 43274 27922 43342 27978
rect 43398 27922 43494 27978
rect 42874 10350 43494 27922
rect 42874 10294 42970 10350
rect 43026 10294 43094 10350
rect 43150 10294 43218 10350
rect 43274 10294 43342 10350
rect 43398 10294 43494 10350
rect 42874 10226 43494 10294
rect 42874 10170 42970 10226
rect 43026 10170 43094 10226
rect 43150 10170 43218 10226
rect 43274 10170 43342 10226
rect 43398 10170 43494 10226
rect 42874 10102 43494 10170
rect 42874 10046 42970 10102
rect 43026 10046 43094 10102
rect 43150 10046 43218 10102
rect 43274 10046 43342 10102
rect 43398 10046 43494 10102
rect 42874 9978 43494 10046
rect 42874 9922 42970 9978
rect 43026 9922 43094 9978
rect 43150 9922 43218 9978
rect 43274 9922 43342 9978
rect 43398 9922 43494 9978
rect 42874 -1120 43494 9922
rect 42874 -1176 42970 -1120
rect 43026 -1176 43094 -1120
rect 43150 -1176 43218 -1120
rect 43274 -1176 43342 -1120
rect 43398 -1176 43494 -1120
rect 42874 -1244 43494 -1176
rect 42874 -1300 42970 -1244
rect 43026 -1300 43094 -1244
rect 43150 -1300 43218 -1244
rect 43274 -1300 43342 -1244
rect 43398 -1300 43494 -1244
rect 42874 -1368 43494 -1300
rect 42874 -1424 42970 -1368
rect 43026 -1424 43094 -1368
rect 43150 -1424 43218 -1368
rect 43274 -1424 43342 -1368
rect 43398 -1424 43494 -1368
rect 42874 -1492 43494 -1424
rect 42874 -1548 42970 -1492
rect 43026 -1548 43094 -1492
rect 43150 -1548 43218 -1492
rect 43274 -1548 43342 -1492
rect 43398 -1548 43494 -1492
rect 42874 -1644 43494 -1548
rect 57154 40350 57774 57922
rect 64448 58350 64768 58384
rect 64448 58294 64518 58350
rect 64574 58294 64642 58350
rect 64698 58294 64768 58350
rect 64448 58226 64768 58294
rect 64448 58170 64518 58226
rect 64574 58170 64642 58226
rect 64698 58170 64768 58226
rect 64448 58102 64768 58170
rect 64448 58046 64518 58102
rect 64574 58046 64642 58102
rect 64698 58046 64768 58102
rect 64448 57978 64768 58046
rect 64448 57922 64518 57978
rect 64574 57922 64642 57978
rect 64698 57922 64768 57978
rect 64448 57888 64768 57922
rect 240874 46350 241494 63922
rect 242732 74564 242788 74574
rect 242732 57428 242788 74508
rect 242844 65492 242900 78988
rect 242844 65426 242900 65436
rect 242956 77924 243012 77934
rect 242956 63476 243012 77868
rect 243068 67508 243124 80108
rect 243180 71540 243236 82348
rect 243180 71474 243236 71484
rect 243292 81284 243348 81294
rect 243292 69524 243348 81228
rect 243292 69458 243348 69468
rect 243068 67442 243124 67452
rect 242956 63410 243012 63420
rect 242732 57362 242788 57372
rect 240874 46294 240970 46350
rect 241026 46294 241094 46350
rect 241150 46294 241218 46350
rect 241274 46294 241342 46350
rect 241398 46294 241494 46350
rect 240874 46226 241494 46294
rect 240874 46170 240970 46226
rect 241026 46170 241094 46226
rect 241150 46170 241218 46226
rect 241274 46170 241342 46226
rect 241398 46170 241494 46226
rect 240874 46102 241494 46170
rect 240874 46046 240970 46102
rect 241026 46046 241094 46102
rect 241150 46046 241218 46102
rect 241274 46046 241342 46102
rect 241398 46046 241494 46102
rect 240874 45978 241494 46046
rect 240874 45922 240970 45978
rect 241026 45922 241094 45978
rect 241150 45922 241218 45978
rect 241274 45922 241342 45978
rect 241398 45922 241494 45978
rect 57154 40294 57250 40350
rect 57306 40294 57374 40350
rect 57430 40294 57498 40350
rect 57554 40294 57622 40350
rect 57678 40294 57774 40350
rect 57154 40226 57774 40294
rect 57154 40170 57250 40226
rect 57306 40170 57374 40226
rect 57430 40170 57498 40226
rect 57554 40170 57622 40226
rect 57678 40170 57774 40226
rect 57154 40102 57774 40170
rect 57154 40046 57250 40102
rect 57306 40046 57374 40102
rect 57430 40046 57498 40102
rect 57554 40046 57622 40102
rect 57678 40046 57774 40102
rect 57154 39978 57774 40046
rect 57154 39922 57250 39978
rect 57306 39922 57374 39978
rect 57430 39922 57498 39978
rect 57554 39922 57622 39978
rect 57678 39922 57774 39978
rect 57154 22350 57774 39922
rect 64448 40350 64768 40384
rect 64448 40294 64518 40350
rect 64574 40294 64642 40350
rect 64698 40294 64768 40350
rect 64448 40226 64768 40294
rect 64448 40170 64518 40226
rect 64574 40170 64642 40226
rect 64698 40170 64768 40226
rect 64448 40102 64768 40170
rect 64448 40046 64518 40102
rect 64574 40046 64642 40102
rect 64698 40046 64768 40102
rect 64448 39978 64768 40046
rect 64448 39922 64518 39978
rect 64574 39922 64642 39978
rect 64698 39922 64768 39978
rect 64448 39888 64768 39922
rect 238476 34498 238532 34508
rect 153468 33238 153524 33248
rect 105084 33012 105140 33022
rect 81788 32900 81844 32910
rect 57154 22294 57250 22350
rect 57306 22294 57374 22350
rect 57430 22294 57498 22350
rect 57554 22294 57622 22350
rect 57678 22294 57774 22350
rect 57154 22226 57774 22294
rect 57154 22170 57250 22226
rect 57306 22170 57374 22226
rect 57430 22170 57498 22226
rect 57554 22170 57622 22226
rect 57678 22170 57774 22226
rect 57154 22102 57774 22170
rect 57154 22046 57250 22102
rect 57306 22046 57374 22102
rect 57430 22046 57498 22102
rect 57554 22046 57622 22102
rect 57678 22046 57774 22102
rect 57154 21978 57774 22046
rect 57154 21922 57250 21978
rect 57306 21922 57374 21978
rect 57430 21922 57498 21978
rect 57554 21922 57622 21978
rect 57678 21922 57774 21978
rect 57154 4350 57774 21922
rect 57154 4294 57250 4350
rect 57306 4294 57374 4350
rect 57430 4294 57498 4350
rect 57554 4294 57622 4350
rect 57678 4294 57774 4350
rect 57154 4226 57774 4294
rect 57154 4170 57250 4226
rect 57306 4170 57374 4226
rect 57430 4170 57498 4226
rect 57554 4170 57622 4226
rect 57678 4170 57774 4226
rect 57154 4102 57774 4170
rect 57154 4046 57250 4102
rect 57306 4046 57374 4102
rect 57430 4046 57498 4102
rect 57554 4046 57622 4102
rect 57678 4046 57774 4102
rect 57154 3978 57774 4046
rect 57154 3922 57250 3978
rect 57306 3922 57374 3978
rect 57430 3922 57498 3978
rect 57554 3922 57622 3978
rect 57678 3922 57774 3978
rect 57154 -160 57774 3922
rect 57154 -216 57250 -160
rect 57306 -216 57374 -160
rect 57430 -216 57498 -160
rect 57554 -216 57622 -160
rect 57678 -216 57774 -160
rect 57154 -284 57774 -216
rect 57154 -340 57250 -284
rect 57306 -340 57374 -284
rect 57430 -340 57498 -284
rect 57554 -340 57622 -284
rect 57678 -340 57774 -284
rect 57154 -408 57774 -340
rect 57154 -464 57250 -408
rect 57306 -464 57374 -408
rect 57430 -464 57498 -408
rect 57554 -464 57622 -408
rect 57678 -464 57774 -408
rect 57154 -532 57774 -464
rect 57154 -588 57250 -532
rect 57306 -588 57374 -532
rect 57430 -588 57498 -532
rect 57554 -588 57622 -532
rect 57678 -588 57774 -532
rect 57154 -1644 57774 -588
rect 60874 28350 61494 31350
rect 60874 28294 60970 28350
rect 61026 28294 61094 28350
rect 61150 28294 61218 28350
rect 61274 28294 61342 28350
rect 61398 28294 61494 28350
rect 60874 28226 61494 28294
rect 60874 28170 60970 28226
rect 61026 28170 61094 28226
rect 61150 28170 61218 28226
rect 61274 28170 61342 28226
rect 61398 28170 61494 28226
rect 60874 28102 61494 28170
rect 60874 28046 60970 28102
rect 61026 28046 61094 28102
rect 61150 28046 61218 28102
rect 61274 28046 61342 28102
rect 61398 28046 61494 28102
rect 60874 27978 61494 28046
rect 60874 27922 60970 27978
rect 61026 27922 61094 27978
rect 61150 27922 61218 27978
rect 61274 27922 61342 27978
rect 61398 27922 61494 27978
rect 60874 10350 61494 27922
rect 73836 26964 73892 26974
rect 73836 20098 73892 26908
rect 73836 20032 73892 20042
rect 75154 22350 75774 31350
rect 75154 22294 75250 22350
rect 75306 22294 75374 22350
rect 75430 22294 75498 22350
rect 75554 22294 75622 22350
rect 75678 22294 75774 22350
rect 75154 22226 75774 22294
rect 75154 22170 75250 22226
rect 75306 22170 75374 22226
rect 75430 22170 75498 22226
rect 75554 22170 75622 22226
rect 75678 22170 75774 22226
rect 75154 22102 75774 22170
rect 75154 22046 75250 22102
rect 75306 22046 75374 22102
rect 75430 22046 75498 22102
rect 75554 22046 75622 22102
rect 75678 22046 75774 22102
rect 75154 21978 75774 22046
rect 75154 21922 75250 21978
rect 75306 21922 75374 21978
rect 75430 21922 75498 21978
rect 75554 21922 75622 21978
rect 75678 21922 75774 21978
rect 60874 10294 60970 10350
rect 61026 10294 61094 10350
rect 61150 10294 61218 10350
rect 61274 10294 61342 10350
rect 61398 10294 61494 10350
rect 60874 10226 61494 10294
rect 60874 10170 60970 10226
rect 61026 10170 61094 10226
rect 61150 10170 61218 10226
rect 61274 10170 61342 10226
rect 61398 10170 61494 10226
rect 60874 10102 61494 10170
rect 60874 10046 60970 10102
rect 61026 10046 61094 10102
rect 61150 10046 61218 10102
rect 61274 10046 61342 10102
rect 61398 10046 61494 10102
rect 60874 9978 61494 10046
rect 60874 9922 60970 9978
rect 61026 9922 61094 9978
rect 61150 9922 61218 9978
rect 61274 9922 61342 9978
rect 61398 9922 61494 9978
rect 60874 -1120 61494 9922
rect 60874 -1176 60970 -1120
rect 61026 -1176 61094 -1120
rect 61150 -1176 61218 -1120
rect 61274 -1176 61342 -1120
rect 61398 -1176 61494 -1120
rect 60874 -1244 61494 -1176
rect 60874 -1300 60970 -1244
rect 61026 -1300 61094 -1244
rect 61150 -1300 61218 -1244
rect 61274 -1300 61342 -1244
rect 61398 -1300 61494 -1244
rect 60874 -1368 61494 -1300
rect 60874 -1424 60970 -1368
rect 61026 -1424 61094 -1368
rect 61150 -1424 61218 -1368
rect 61274 -1424 61342 -1368
rect 61398 -1424 61494 -1368
rect 60874 -1492 61494 -1424
rect 60874 -1548 60970 -1492
rect 61026 -1548 61094 -1492
rect 61150 -1548 61218 -1492
rect 61274 -1548 61342 -1492
rect 61398 -1548 61494 -1492
rect 60874 -1644 61494 -1548
rect 75154 4350 75774 21922
rect 75154 4294 75250 4350
rect 75306 4294 75374 4350
rect 75430 4294 75498 4350
rect 75554 4294 75622 4350
rect 75678 4294 75774 4350
rect 75154 4226 75774 4294
rect 75154 4170 75250 4226
rect 75306 4170 75374 4226
rect 75430 4170 75498 4226
rect 75554 4170 75622 4226
rect 75678 4170 75774 4226
rect 75154 4102 75774 4170
rect 75154 4046 75250 4102
rect 75306 4046 75374 4102
rect 75430 4046 75498 4102
rect 75554 4046 75622 4102
rect 75678 4046 75774 4102
rect 75154 3978 75774 4046
rect 75154 3922 75250 3978
rect 75306 3922 75374 3978
rect 75430 3922 75498 3978
rect 75554 3922 75622 3978
rect 75678 3922 75774 3978
rect 75154 -160 75774 3922
rect 75154 -216 75250 -160
rect 75306 -216 75374 -160
rect 75430 -216 75498 -160
rect 75554 -216 75622 -160
rect 75678 -216 75774 -160
rect 75154 -284 75774 -216
rect 75154 -340 75250 -284
rect 75306 -340 75374 -284
rect 75430 -340 75498 -284
rect 75554 -340 75622 -284
rect 75678 -340 75774 -284
rect 75154 -408 75774 -340
rect 75154 -464 75250 -408
rect 75306 -464 75374 -408
rect 75430 -464 75498 -408
rect 75554 -464 75622 -408
rect 75678 -464 75774 -408
rect 75154 -532 75774 -464
rect 75154 -588 75250 -532
rect 75306 -588 75374 -532
rect 75430 -588 75498 -532
rect 75554 -588 75622 -532
rect 75678 -588 75774 -532
rect 75154 -1644 75774 -588
rect 78874 28350 79494 31350
rect 81788 30100 81844 32844
rect 81788 30034 81844 30044
rect 78874 28294 78970 28350
rect 79026 28294 79094 28350
rect 79150 28294 79218 28350
rect 79274 28294 79342 28350
rect 79398 28294 79494 28350
rect 78874 28226 79494 28294
rect 78874 28170 78970 28226
rect 79026 28170 79094 28226
rect 79150 28170 79218 28226
rect 79274 28170 79342 28226
rect 79398 28170 79494 28226
rect 78874 28102 79494 28170
rect 78874 28046 78970 28102
rect 79026 28046 79094 28102
rect 79150 28046 79218 28102
rect 79274 28046 79342 28102
rect 79398 28046 79494 28102
rect 78874 27978 79494 28046
rect 78874 27922 78970 27978
rect 79026 27922 79094 27978
rect 79150 27922 79218 27978
rect 79274 27922 79342 27978
rect 79398 27922 79494 27978
rect 78874 10350 79494 27922
rect 78874 10294 78970 10350
rect 79026 10294 79094 10350
rect 79150 10294 79218 10350
rect 79274 10294 79342 10350
rect 79398 10294 79494 10350
rect 78874 10226 79494 10294
rect 78874 10170 78970 10226
rect 79026 10170 79094 10226
rect 79150 10170 79218 10226
rect 79274 10170 79342 10226
rect 79398 10170 79494 10226
rect 78874 10102 79494 10170
rect 78874 10046 78970 10102
rect 79026 10046 79094 10102
rect 79150 10046 79218 10102
rect 79274 10046 79342 10102
rect 79398 10046 79494 10102
rect 78874 9978 79494 10046
rect 78874 9922 78970 9978
rect 79026 9922 79094 9978
rect 79150 9922 79218 9978
rect 79274 9922 79342 9978
rect 79398 9922 79494 9978
rect 78874 -1120 79494 9922
rect 80668 27412 80724 27422
rect 80668 7588 80724 27356
rect 80668 7522 80724 7532
rect 93154 22350 93774 31350
rect 93154 22294 93250 22350
rect 93306 22294 93374 22350
rect 93430 22294 93498 22350
rect 93554 22294 93622 22350
rect 93678 22294 93774 22350
rect 93154 22226 93774 22294
rect 93154 22170 93250 22226
rect 93306 22170 93374 22226
rect 93430 22170 93498 22226
rect 93554 22170 93622 22226
rect 93678 22170 93774 22226
rect 93154 22102 93774 22170
rect 93154 22046 93250 22102
rect 93306 22046 93374 22102
rect 93430 22046 93498 22102
rect 93554 22046 93622 22102
rect 93678 22046 93774 22102
rect 93154 21978 93774 22046
rect 93154 21922 93250 21978
rect 93306 21922 93374 21978
rect 93430 21922 93498 21978
rect 93554 21922 93622 21978
rect 93678 21922 93774 21978
rect 78874 -1176 78970 -1120
rect 79026 -1176 79094 -1120
rect 79150 -1176 79218 -1120
rect 79274 -1176 79342 -1120
rect 79398 -1176 79494 -1120
rect 78874 -1244 79494 -1176
rect 78874 -1300 78970 -1244
rect 79026 -1300 79094 -1244
rect 79150 -1300 79218 -1244
rect 79274 -1300 79342 -1244
rect 79398 -1300 79494 -1244
rect 78874 -1368 79494 -1300
rect 78874 -1424 78970 -1368
rect 79026 -1424 79094 -1368
rect 79150 -1424 79218 -1368
rect 79274 -1424 79342 -1368
rect 79398 -1424 79494 -1368
rect 78874 -1492 79494 -1424
rect 78874 -1548 78970 -1492
rect 79026 -1548 79094 -1492
rect 79150 -1548 79218 -1492
rect 79274 -1548 79342 -1492
rect 79398 -1548 79494 -1492
rect 78874 -1644 79494 -1548
rect 93154 4350 93774 21922
rect 93154 4294 93250 4350
rect 93306 4294 93374 4350
rect 93430 4294 93498 4350
rect 93554 4294 93622 4350
rect 93678 4294 93774 4350
rect 93154 4226 93774 4294
rect 93154 4170 93250 4226
rect 93306 4170 93374 4226
rect 93430 4170 93498 4226
rect 93554 4170 93622 4226
rect 93678 4170 93774 4226
rect 93154 4102 93774 4170
rect 93154 4046 93250 4102
rect 93306 4046 93374 4102
rect 93430 4046 93498 4102
rect 93554 4046 93622 4102
rect 93678 4046 93774 4102
rect 93154 3978 93774 4046
rect 93154 3922 93250 3978
rect 93306 3922 93374 3978
rect 93430 3922 93498 3978
rect 93554 3922 93622 3978
rect 93678 3922 93774 3978
rect 93154 -160 93774 3922
rect 93154 -216 93250 -160
rect 93306 -216 93374 -160
rect 93430 -216 93498 -160
rect 93554 -216 93622 -160
rect 93678 -216 93774 -160
rect 93154 -284 93774 -216
rect 93154 -340 93250 -284
rect 93306 -340 93374 -284
rect 93430 -340 93498 -284
rect 93554 -340 93622 -284
rect 93678 -340 93774 -284
rect 93154 -408 93774 -340
rect 93154 -464 93250 -408
rect 93306 -464 93374 -408
rect 93430 -464 93498 -408
rect 93554 -464 93622 -408
rect 93678 -464 93774 -408
rect 93154 -532 93774 -464
rect 93154 -588 93250 -532
rect 93306 -588 93374 -532
rect 93430 -588 93498 -532
rect 93554 -588 93622 -532
rect 93678 -588 93774 -532
rect 93154 -1644 93774 -588
rect 96874 28350 97494 31350
rect 105084 30324 105140 32956
rect 151676 32788 151732 32798
rect 140812 31798 140868 31808
rect 139132 31618 139188 31628
rect 105084 30258 105140 30268
rect 96874 28294 96970 28350
rect 97026 28294 97094 28350
rect 97150 28294 97218 28350
rect 97274 28294 97342 28350
rect 97398 28294 97494 28350
rect 96874 28226 97494 28294
rect 96874 28170 96970 28226
rect 97026 28170 97094 28226
rect 97150 28170 97218 28226
rect 97274 28170 97342 28226
rect 97398 28170 97494 28226
rect 96874 28102 97494 28170
rect 96874 28046 96970 28102
rect 97026 28046 97094 28102
rect 97150 28046 97218 28102
rect 97274 28046 97342 28102
rect 97398 28046 97494 28102
rect 96874 27978 97494 28046
rect 96874 27922 96970 27978
rect 97026 27922 97094 27978
rect 97150 27922 97218 27978
rect 97274 27922 97342 27978
rect 97398 27922 97494 27978
rect 96874 10350 97494 27922
rect 110460 28532 110516 28542
rect 96874 10294 96970 10350
rect 97026 10294 97094 10350
rect 97150 10294 97218 10350
rect 97274 10294 97342 10350
rect 97398 10294 97494 10350
rect 96874 10226 97494 10294
rect 96874 10170 96970 10226
rect 97026 10170 97094 10226
rect 97150 10170 97218 10226
rect 97274 10170 97342 10226
rect 97398 10170 97494 10226
rect 96874 10102 97494 10170
rect 96874 10046 96970 10102
rect 97026 10046 97094 10102
rect 97150 10046 97218 10102
rect 97274 10046 97342 10102
rect 97398 10046 97494 10102
rect 96874 9978 97494 10046
rect 96874 9922 96970 9978
rect 97026 9922 97094 9978
rect 97150 9922 97218 9978
rect 97274 9922 97342 9978
rect 97398 9922 97494 9978
rect 96874 -1120 97494 9922
rect 104188 27412 104244 27422
rect 104188 5908 104244 27356
rect 110460 26938 110516 28476
rect 110460 26872 110516 26882
rect 104188 5842 104244 5852
rect 111154 22350 111774 31350
rect 112252 28532 112308 28542
rect 112252 27658 112308 28476
rect 112252 27592 112308 27602
rect 114874 28350 115494 31350
rect 114874 28294 114970 28350
rect 115026 28294 115094 28350
rect 115150 28294 115218 28350
rect 115274 28294 115342 28350
rect 115398 28294 115494 28350
rect 114874 28226 115494 28294
rect 114874 28170 114970 28226
rect 115026 28170 115094 28226
rect 115150 28170 115218 28226
rect 115274 28170 115342 28226
rect 115398 28170 115494 28226
rect 114874 28102 115494 28170
rect 114874 28046 114970 28102
rect 115026 28046 115094 28102
rect 115150 28046 115218 28102
rect 115274 28046 115342 28102
rect 115398 28046 115494 28102
rect 114874 27978 115494 28046
rect 114874 27922 114970 27978
rect 115026 27922 115094 27978
rect 115150 27922 115218 27978
rect 115274 27922 115342 27978
rect 115398 27922 115494 27978
rect 111154 22294 111250 22350
rect 111306 22294 111374 22350
rect 111430 22294 111498 22350
rect 111554 22294 111622 22350
rect 111678 22294 111774 22350
rect 111154 22226 111774 22294
rect 111154 22170 111250 22226
rect 111306 22170 111374 22226
rect 111430 22170 111498 22226
rect 111554 22170 111622 22226
rect 111678 22170 111774 22226
rect 111154 22102 111774 22170
rect 111154 22046 111250 22102
rect 111306 22046 111374 22102
rect 111430 22046 111498 22102
rect 111554 22046 111622 22102
rect 111678 22046 111774 22102
rect 111154 21978 111774 22046
rect 111154 21922 111250 21978
rect 111306 21922 111374 21978
rect 111430 21922 111498 21978
rect 111554 21922 111622 21978
rect 111678 21922 111774 21978
rect 96874 -1176 96970 -1120
rect 97026 -1176 97094 -1120
rect 97150 -1176 97218 -1120
rect 97274 -1176 97342 -1120
rect 97398 -1176 97494 -1120
rect 96874 -1244 97494 -1176
rect 96874 -1300 96970 -1244
rect 97026 -1300 97094 -1244
rect 97150 -1300 97218 -1244
rect 97274 -1300 97342 -1244
rect 97398 -1300 97494 -1244
rect 96874 -1368 97494 -1300
rect 96874 -1424 96970 -1368
rect 97026 -1424 97094 -1368
rect 97150 -1424 97218 -1368
rect 97274 -1424 97342 -1368
rect 97398 -1424 97494 -1368
rect 96874 -1492 97494 -1424
rect 96874 -1548 96970 -1492
rect 97026 -1548 97094 -1492
rect 97150 -1548 97218 -1492
rect 97274 -1548 97342 -1492
rect 97398 -1548 97494 -1492
rect 96874 -1644 97494 -1548
rect 111154 4350 111774 21922
rect 111154 4294 111250 4350
rect 111306 4294 111374 4350
rect 111430 4294 111498 4350
rect 111554 4294 111622 4350
rect 111678 4294 111774 4350
rect 111154 4226 111774 4294
rect 111154 4170 111250 4226
rect 111306 4170 111374 4226
rect 111430 4170 111498 4226
rect 111554 4170 111622 4226
rect 111678 4170 111774 4226
rect 111154 4102 111774 4170
rect 111154 4046 111250 4102
rect 111306 4046 111374 4102
rect 111430 4046 111498 4102
rect 111554 4046 111622 4102
rect 111678 4046 111774 4102
rect 111154 3978 111774 4046
rect 111154 3922 111250 3978
rect 111306 3922 111374 3978
rect 111430 3922 111498 3978
rect 111554 3922 111622 3978
rect 111678 3922 111774 3978
rect 111154 -160 111774 3922
rect 111154 -216 111250 -160
rect 111306 -216 111374 -160
rect 111430 -216 111498 -160
rect 111554 -216 111622 -160
rect 111678 -216 111774 -160
rect 111154 -284 111774 -216
rect 111154 -340 111250 -284
rect 111306 -340 111374 -284
rect 111430 -340 111498 -284
rect 111554 -340 111622 -284
rect 111678 -340 111774 -284
rect 111154 -408 111774 -340
rect 111154 -464 111250 -408
rect 111306 -464 111374 -408
rect 111430 -464 111498 -408
rect 111554 -464 111622 -408
rect 111678 -464 111774 -408
rect 111154 -532 111774 -464
rect 111154 -588 111250 -532
rect 111306 -588 111374 -532
rect 111430 -588 111498 -532
rect 111554 -588 111622 -532
rect 111678 -588 111774 -532
rect 111154 -1644 111774 -588
rect 114874 10350 115494 27922
rect 114874 10294 114970 10350
rect 115026 10294 115094 10350
rect 115150 10294 115218 10350
rect 115274 10294 115342 10350
rect 115398 10294 115494 10350
rect 114874 10226 115494 10294
rect 114874 10170 114970 10226
rect 115026 10170 115094 10226
rect 115150 10170 115218 10226
rect 115274 10170 115342 10226
rect 115398 10170 115494 10226
rect 114874 10102 115494 10170
rect 114874 10046 114970 10102
rect 115026 10046 115094 10102
rect 115150 10046 115218 10102
rect 115274 10046 115342 10102
rect 115398 10046 115494 10102
rect 114874 9978 115494 10046
rect 114874 9922 114970 9978
rect 115026 9922 115094 9978
rect 115150 9922 115218 9978
rect 115274 9922 115342 9978
rect 115398 9922 115494 9978
rect 114874 -1120 115494 9922
rect 114874 -1176 114970 -1120
rect 115026 -1176 115094 -1120
rect 115150 -1176 115218 -1120
rect 115274 -1176 115342 -1120
rect 115398 -1176 115494 -1120
rect 114874 -1244 115494 -1176
rect 114874 -1300 114970 -1244
rect 115026 -1300 115094 -1244
rect 115150 -1300 115218 -1244
rect 115274 -1300 115342 -1244
rect 115398 -1300 115494 -1244
rect 114874 -1368 115494 -1300
rect 114874 -1424 114970 -1368
rect 115026 -1424 115094 -1368
rect 115150 -1424 115218 -1368
rect 115274 -1424 115342 -1368
rect 115398 -1424 115494 -1368
rect 114874 -1492 115494 -1424
rect 114874 -1548 114970 -1492
rect 115026 -1548 115094 -1492
rect 115150 -1548 115218 -1492
rect 115274 -1548 115342 -1492
rect 115398 -1548 115494 -1492
rect 114874 -1644 115494 -1548
rect 129154 22350 129774 31350
rect 129154 22294 129250 22350
rect 129306 22294 129374 22350
rect 129430 22294 129498 22350
rect 129554 22294 129622 22350
rect 129678 22294 129774 22350
rect 129154 22226 129774 22294
rect 129154 22170 129250 22226
rect 129306 22170 129374 22226
rect 129430 22170 129498 22226
rect 129554 22170 129622 22226
rect 129678 22170 129774 22226
rect 129154 22102 129774 22170
rect 129154 22046 129250 22102
rect 129306 22046 129374 22102
rect 129430 22046 129498 22102
rect 129554 22046 129622 22102
rect 129678 22046 129774 22102
rect 129154 21978 129774 22046
rect 129154 21922 129250 21978
rect 129306 21922 129374 21978
rect 129430 21922 129498 21978
rect 129554 21922 129622 21978
rect 129678 21922 129774 21978
rect 129154 4350 129774 21922
rect 129154 4294 129250 4350
rect 129306 4294 129374 4350
rect 129430 4294 129498 4350
rect 129554 4294 129622 4350
rect 129678 4294 129774 4350
rect 129154 4226 129774 4294
rect 129154 4170 129250 4226
rect 129306 4170 129374 4226
rect 129430 4170 129498 4226
rect 129554 4170 129622 4226
rect 129678 4170 129774 4226
rect 129154 4102 129774 4170
rect 129154 4046 129250 4102
rect 129306 4046 129374 4102
rect 129430 4046 129498 4102
rect 129554 4046 129622 4102
rect 129678 4046 129774 4102
rect 129154 3978 129774 4046
rect 129154 3922 129250 3978
rect 129306 3922 129374 3978
rect 129430 3922 129498 3978
rect 129554 3922 129622 3978
rect 129678 3922 129774 3978
rect 129154 -160 129774 3922
rect 129154 -216 129250 -160
rect 129306 -216 129374 -160
rect 129430 -216 129498 -160
rect 129554 -216 129622 -160
rect 129678 -216 129774 -160
rect 129154 -284 129774 -216
rect 129154 -340 129250 -284
rect 129306 -340 129374 -284
rect 129430 -340 129498 -284
rect 129554 -340 129622 -284
rect 129678 -340 129774 -284
rect 129154 -408 129774 -340
rect 129154 -464 129250 -408
rect 129306 -464 129374 -408
rect 129430 -464 129498 -408
rect 129554 -464 129622 -408
rect 129678 -464 129774 -408
rect 129154 -532 129774 -464
rect 129154 -588 129250 -532
rect 129306 -588 129374 -532
rect 129430 -588 129498 -532
rect 129554 -588 129622 -532
rect 129678 -588 129774 -532
rect 129154 -1644 129774 -588
rect 132874 28350 133494 31350
rect 139132 30772 139188 31562
rect 132874 28294 132970 28350
rect 133026 28294 133094 28350
rect 133150 28294 133218 28350
rect 133274 28294 133342 28350
rect 133398 28294 133494 28350
rect 132874 28226 133494 28294
rect 132874 28170 132970 28226
rect 133026 28170 133094 28226
rect 133150 28170 133218 28226
rect 133274 28170 133342 28226
rect 133398 28170 133494 28226
rect 132874 28102 133494 28170
rect 132874 28046 132970 28102
rect 133026 28046 133094 28102
rect 133150 28046 133218 28102
rect 133274 28046 133342 28102
rect 133398 28046 133494 28102
rect 132874 27978 133494 28046
rect 132874 27922 132970 27978
rect 133026 27922 133094 27978
rect 133150 27922 133218 27978
rect 133274 27922 133342 27978
rect 133398 27922 133494 27978
rect 132874 10350 133494 27922
rect 137788 28532 137844 28542
rect 137788 19796 137844 28476
rect 139132 28532 139188 30716
rect 139132 28466 139188 28476
rect 139580 28532 139636 28542
rect 137788 19730 137844 19740
rect 132874 10294 132970 10350
rect 133026 10294 133094 10350
rect 133150 10294 133218 10350
rect 133274 10294 133342 10350
rect 133398 10294 133494 10350
rect 132874 10226 133494 10294
rect 132874 10170 132970 10226
rect 133026 10170 133094 10226
rect 133150 10170 133218 10226
rect 133274 10170 133342 10226
rect 133398 10170 133494 10226
rect 132874 10102 133494 10170
rect 132874 10046 132970 10102
rect 133026 10046 133094 10102
rect 133150 10046 133218 10102
rect 133274 10046 133342 10102
rect 133398 10046 133494 10102
rect 132874 9978 133494 10046
rect 132874 9922 132970 9978
rect 133026 9922 133094 9978
rect 133150 9922 133218 9978
rect 133274 9922 133342 9978
rect 133398 9922 133494 9978
rect 132874 -1120 133494 9922
rect 139580 6244 139636 28476
rect 140812 28420 140868 31742
rect 140924 31438 140980 31448
rect 140924 30772 140980 31382
rect 140924 28532 140980 30716
rect 142716 31258 142772 31268
rect 142716 30772 142772 31202
rect 140924 28466 140980 28476
rect 141148 28532 141204 28542
rect 140812 28354 140868 28364
rect 141148 16324 141204 28476
rect 142716 28532 142772 30716
rect 142716 28466 142772 28476
rect 144508 26628 144564 26638
rect 144508 26068 144564 26572
rect 144508 26002 144564 26012
rect 141148 16258 141204 16268
rect 147154 22350 147774 31350
rect 149884 31078 149940 31088
rect 149884 30772 149940 31022
rect 147868 29818 147924 29828
rect 147868 29698 147924 29708
rect 147154 22294 147250 22350
rect 147306 22294 147374 22350
rect 147430 22294 147498 22350
rect 147554 22294 147622 22350
rect 147678 22294 147774 22350
rect 147154 22226 147774 22294
rect 147154 22170 147250 22226
rect 147306 22170 147374 22226
rect 147430 22170 147498 22226
rect 147554 22170 147622 22226
rect 147678 22170 147774 22226
rect 147154 22102 147774 22170
rect 147154 22046 147250 22102
rect 147306 22046 147374 22102
rect 147430 22046 147498 22102
rect 147554 22046 147622 22102
rect 147678 22046 147774 22102
rect 147154 21978 147774 22046
rect 147154 21922 147250 21978
rect 147306 21922 147374 21978
rect 147430 21922 147498 21978
rect 147554 21922 147622 21978
rect 147678 21922 147774 21978
rect 139580 6178 139636 6188
rect 132874 -1176 132970 -1120
rect 133026 -1176 133094 -1120
rect 133150 -1176 133218 -1120
rect 133274 -1176 133342 -1120
rect 133398 -1176 133494 -1120
rect 132874 -1244 133494 -1176
rect 132874 -1300 132970 -1244
rect 133026 -1300 133094 -1244
rect 133150 -1300 133218 -1244
rect 133274 -1300 133342 -1244
rect 133398 -1300 133494 -1244
rect 132874 -1368 133494 -1300
rect 132874 -1424 132970 -1368
rect 133026 -1424 133094 -1368
rect 133150 -1424 133218 -1368
rect 133274 -1424 133342 -1368
rect 133398 -1424 133494 -1368
rect 132874 -1492 133494 -1424
rect 132874 -1548 132970 -1492
rect 133026 -1548 133094 -1492
rect 133150 -1548 133218 -1492
rect 133274 -1548 133342 -1492
rect 133398 -1548 133494 -1492
rect 132874 -1644 133494 -1548
rect 147154 4350 147774 21922
rect 147868 26964 147924 26974
rect 147868 12852 147924 26908
rect 149884 19572 149940 30716
rect 149884 19506 149940 19516
rect 150874 28350 151494 31350
rect 151676 30660 151732 32732
rect 151676 30594 151732 30604
rect 153468 30660 153524 33182
rect 153468 30594 153524 30604
rect 158844 33058 158900 33068
rect 158844 30660 158900 33002
rect 158844 30594 158900 30604
rect 160636 32878 160692 32888
rect 160636 30660 160692 32822
rect 160636 30594 160692 30604
rect 162428 32698 162484 32708
rect 162428 30660 162484 32642
rect 223580 32676 223636 32686
rect 191100 32564 191156 32574
rect 162428 30594 162484 30604
rect 157052 30178 157108 30188
rect 150874 28294 150970 28350
rect 151026 28294 151094 28350
rect 151150 28294 151218 28350
rect 151274 28294 151342 28350
rect 151398 28294 151494 28350
rect 150874 28226 151494 28294
rect 150874 28170 150970 28226
rect 151026 28170 151094 28226
rect 151150 28170 151218 28226
rect 151274 28170 151342 28226
rect 151398 28170 151494 28226
rect 150874 28102 151494 28170
rect 150874 28046 150970 28102
rect 151026 28046 151094 28102
rect 151150 28046 151218 28102
rect 151274 28046 151342 28102
rect 151398 28046 151494 28102
rect 150874 27978 151494 28046
rect 150874 27922 150970 27978
rect 151026 27922 151094 27978
rect 151150 27922 151218 27978
rect 151274 27922 151342 27978
rect 151398 27922 151494 27978
rect 147868 12786 147924 12796
rect 147154 4294 147250 4350
rect 147306 4294 147374 4350
rect 147430 4294 147498 4350
rect 147554 4294 147622 4350
rect 147678 4294 147774 4350
rect 147154 4226 147774 4294
rect 147154 4170 147250 4226
rect 147306 4170 147374 4226
rect 147430 4170 147498 4226
rect 147554 4170 147622 4226
rect 147678 4170 147774 4226
rect 147154 4102 147774 4170
rect 147154 4046 147250 4102
rect 147306 4046 147374 4102
rect 147430 4046 147498 4102
rect 147554 4046 147622 4102
rect 147678 4046 147774 4102
rect 147154 3978 147774 4046
rect 147154 3922 147250 3978
rect 147306 3922 147374 3978
rect 147430 3922 147498 3978
rect 147554 3922 147622 3978
rect 147678 3922 147774 3978
rect 147154 -160 147774 3922
rect 147154 -216 147250 -160
rect 147306 -216 147374 -160
rect 147430 -216 147498 -160
rect 147554 -216 147622 -160
rect 147678 -216 147774 -160
rect 147154 -284 147774 -216
rect 147154 -340 147250 -284
rect 147306 -340 147374 -284
rect 147430 -340 147498 -284
rect 147554 -340 147622 -284
rect 147678 -340 147774 -284
rect 147154 -408 147774 -340
rect 147154 -464 147250 -408
rect 147306 -464 147374 -408
rect 147430 -464 147498 -408
rect 147554 -464 147622 -408
rect 147678 -464 147774 -408
rect 147154 -532 147774 -464
rect 147154 -588 147250 -532
rect 147306 -588 147374 -532
rect 147430 -588 147498 -532
rect 147554 -588 147622 -532
rect 147678 -588 147774 -532
rect 147154 -1644 147774 -588
rect 150874 10350 151494 27922
rect 155260 29998 155316 30008
rect 155260 28308 155316 29942
rect 157052 29764 157108 30122
rect 157052 29698 157108 29708
rect 155260 24612 155316 28252
rect 158844 27972 158900 27982
rect 155260 24546 155316 24556
rect 156268 26964 156324 26974
rect 156268 14532 156324 26908
rect 158844 21364 158900 27916
rect 158844 21298 158900 21308
rect 159628 27412 159684 27422
rect 159628 17668 159684 27356
rect 159628 17602 159684 17612
rect 161420 27412 161476 27422
rect 161420 16100 161476 27356
rect 161420 16034 161476 16044
rect 165154 22350 165774 31350
rect 165154 22294 165250 22350
rect 165306 22294 165374 22350
rect 165430 22294 165498 22350
rect 165554 22294 165622 22350
rect 165678 22294 165774 22350
rect 165154 22226 165774 22294
rect 165154 22170 165250 22226
rect 165306 22170 165374 22226
rect 165430 22170 165498 22226
rect 165554 22170 165622 22226
rect 165678 22170 165774 22226
rect 165154 22102 165774 22170
rect 165154 22046 165250 22102
rect 165306 22046 165374 22102
rect 165430 22046 165498 22102
rect 165554 22046 165622 22102
rect 165678 22046 165774 22102
rect 165154 21978 165774 22046
rect 165154 21922 165250 21978
rect 165306 21922 165374 21978
rect 165430 21922 165498 21978
rect 165554 21922 165622 21978
rect 165678 21922 165774 21978
rect 156268 14466 156324 14476
rect 150874 10294 150970 10350
rect 151026 10294 151094 10350
rect 151150 10294 151218 10350
rect 151274 10294 151342 10350
rect 151398 10294 151494 10350
rect 150874 10226 151494 10294
rect 150874 10170 150970 10226
rect 151026 10170 151094 10226
rect 151150 10170 151218 10226
rect 151274 10170 151342 10226
rect 151398 10170 151494 10226
rect 150874 10102 151494 10170
rect 150874 10046 150970 10102
rect 151026 10046 151094 10102
rect 151150 10046 151218 10102
rect 151274 10046 151342 10102
rect 151398 10046 151494 10102
rect 150874 9978 151494 10046
rect 150874 9922 150970 9978
rect 151026 9922 151094 9978
rect 151150 9922 151218 9978
rect 151274 9922 151342 9978
rect 151398 9922 151494 9978
rect 150874 -1120 151494 9922
rect 150874 -1176 150970 -1120
rect 151026 -1176 151094 -1120
rect 151150 -1176 151218 -1120
rect 151274 -1176 151342 -1120
rect 151398 -1176 151494 -1120
rect 150874 -1244 151494 -1176
rect 150874 -1300 150970 -1244
rect 151026 -1300 151094 -1244
rect 151150 -1300 151218 -1244
rect 151274 -1300 151342 -1244
rect 151398 -1300 151494 -1244
rect 150874 -1368 151494 -1300
rect 150874 -1424 150970 -1368
rect 151026 -1424 151094 -1368
rect 151150 -1424 151218 -1368
rect 151274 -1424 151342 -1368
rect 151398 -1424 151494 -1368
rect 150874 -1492 151494 -1424
rect 150874 -1548 150970 -1492
rect 151026 -1548 151094 -1492
rect 151150 -1548 151218 -1492
rect 151274 -1548 151342 -1492
rect 151398 -1548 151494 -1492
rect 150874 -1644 151494 -1548
rect 165154 4350 165774 21922
rect 165154 4294 165250 4350
rect 165306 4294 165374 4350
rect 165430 4294 165498 4350
rect 165554 4294 165622 4350
rect 165678 4294 165774 4350
rect 165154 4226 165774 4294
rect 165154 4170 165250 4226
rect 165306 4170 165374 4226
rect 165430 4170 165498 4226
rect 165554 4170 165622 4226
rect 165678 4170 165774 4226
rect 165154 4102 165774 4170
rect 165154 4046 165250 4102
rect 165306 4046 165374 4102
rect 165430 4046 165498 4102
rect 165554 4046 165622 4102
rect 165678 4046 165774 4102
rect 165154 3978 165774 4046
rect 165154 3922 165250 3978
rect 165306 3922 165374 3978
rect 165430 3922 165498 3978
rect 165554 3922 165622 3978
rect 165678 3922 165774 3978
rect 165154 -160 165774 3922
rect 165154 -216 165250 -160
rect 165306 -216 165374 -160
rect 165430 -216 165498 -160
rect 165554 -216 165622 -160
rect 165678 -216 165774 -160
rect 165154 -284 165774 -216
rect 165154 -340 165250 -284
rect 165306 -340 165374 -284
rect 165430 -340 165498 -284
rect 165554 -340 165622 -284
rect 165678 -340 165774 -284
rect 165154 -408 165774 -340
rect 165154 -464 165250 -408
rect 165306 -464 165374 -408
rect 165430 -464 165498 -408
rect 165554 -464 165622 -408
rect 165678 -464 165774 -408
rect 165154 -532 165774 -464
rect 165154 -588 165250 -532
rect 165306 -588 165374 -532
rect 165430 -588 165498 -532
rect 165554 -588 165622 -532
rect 165678 -588 165774 -532
rect 165154 -1644 165774 -588
rect 168874 28350 169494 31350
rect 168874 28294 168970 28350
rect 169026 28294 169094 28350
rect 169150 28294 169218 28350
rect 169274 28294 169342 28350
rect 169398 28294 169494 28350
rect 168874 28226 169494 28294
rect 168874 28170 168970 28226
rect 169026 28170 169094 28226
rect 169150 28170 169218 28226
rect 169274 28170 169342 28226
rect 169398 28170 169494 28226
rect 168874 28102 169494 28170
rect 168874 28046 168970 28102
rect 169026 28046 169094 28102
rect 169150 28046 169218 28102
rect 169274 28046 169342 28102
rect 169398 28046 169494 28102
rect 168874 27978 169494 28046
rect 168874 27922 168970 27978
rect 169026 27922 169094 27978
rect 169150 27922 169218 27978
rect 169274 27922 169342 27978
rect 169398 27922 169494 27978
rect 168874 10350 169494 27922
rect 168874 10294 168970 10350
rect 169026 10294 169094 10350
rect 169150 10294 169218 10350
rect 169274 10294 169342 10350
rect 169398 10294 169494 10350
rect 168874 10226 169494 10294
rect 168874 10170 168970 10226
rect 169026 10170 169094 10226
rect 169150 10170 169218 10226
rect 169274 10170 169342 10226
rect 169398 10170 169494 10226
rect 168874 10102 169494 10170
rect 168874 10046 168970 10102
rect 169026 10046 169094 10102
rect 169150 10046 169218 10102
rect 169274 10046 169342 10102
rect 169398 10046 169494 10102
rect 168874 9978 169494 10046
rect 168874 9922 168970 9978
rect 169026 9922 169094 9978
rect 169150 9922 169218 9978
rect 169274 9922 169342 9978
rect 169398 9922 169494 9978
rect 168874 -1120 169494 9922
rect 168874 -1176 168970 -1120
rect 169026 -1176 169094 -1120
rect 169150 -1176 169218 -1120
rect 169274 -1176 169342 -1120
rect 169398 -1176 169494 -1120
rect 168874 -1244 169494 -1176
rect 168874 -1300 168970 -1244
rect 169026 -1300 169094 -1244
rect 169150 -1300 169218 -1244
rect 169274 -1300 169342 -1244
rect 169398 -1300 169494 -1244
rect 168874 -1368 169494 -1300
rect 168874 -1424 168970 -1368
rect 169026 -1424 169094 -1368
rect 169150 -1424 169218 -1368
rect 169274 -1424 169342 -1368
rect 169398 -1424 169494 -1368
rect 168874 -1492 169494 -1424
rect 168874 -1548 168970 -1492
rect 169026 -1548 169094 -1492
rect 169150 -1548 169218 -1492
rect 169274 -1548 169342 -1492
rect 169398 -1548 169494 -1492
rect 168874 -1644 169494 -1548
rect 183154 22350 183774 31350
rect 186508 29458 186564 29468
rect 186508 27972 186564 29402
rect 186508 27906 186564 27916
rect 186874 28350 187494 30964
rect 188412 30884 188468 30894
rect 188412 29764 188468 30828
rect 191100 30660 191156 32508
rect 191100 30594 191156 30604
rect 194124 32452 194180 32462
rect 188412 29698 188468 29708
rect 194124 28532 194180 32396
rect 209916 31556 209972 31566
rect 200060 31444 200116 31454
rect 198268 31332 198324 31342
rect 196476 31220 196532 31230
rect 196476 30660 196532 31164
rect 196476 30594 196532 30604
rect 198268 30660 198324 31276
rect 198268 30594 198324 30604
rect 200060 30660 200116 31388
rect 200060 30594 200116 30604
rect 194124 28466 194180 28476
rect 186874 28294 186970 28350
rect 187026 28294 187094 28350
rect 187150 28294 187218 28350
rect 187274 28294 187342 28350
rect 187398 28294 187494 28350
rect 186874 28226 187494 28294
rect 186874 28170 186970 28226
rect 187026 28170 187094 28226
rect 187150 28170 187218 28226
rect 187274 28170 187342 28226
rect 187398 28170 187494 28226
rect 186874 28102 187494 28170
rect 186874 28046 186970 28102
rect 187026 28046 187094 28102
rect 187150 28046 187218 28102
rect 187274 28046 187342 28102
rect 187398 28046 187494 28102
rect 186874 27978 187494 28046
rect 186874 27922 186970 27978
rect 187026 27922 187094 27978
rect 187150 27922 187218 27978
rect 187274 27922 187342 27978
rect 187398 27922 187494 27978
rect 183154 22294 183250 22350
rect 183306 22294 183374 22350
rect 183430 22294 183498 22350
rect 183554 22294 183622 22350
rect 183678 22294 183774 22350
rect 183154 22226 183774 22294
rect 183154 22170 183250 22226
rect 183306 22170 183374 22226
rect 183430 22170 183498 22226
rect 183554 22170 183622 22226
rect 183678 22170 183774 22226
rect 183154 22102 183774 22170
rect 183154 22046 183250 22102
rect 183306 22046 183374 22102
rect 183430 22046 183498 22102
rect 183554 22046 183622 22102
rect 183678 22046 183774 22102
rect 183154 21978 183774 22046
rect 183154 21922 183250 21978
rect 183306 21922 183374 21978
rect 183430 21922 183498 21978
rect 183554 21922 183622 21978
rect 183678 21922 183774 21978
rect 183154 4350 183774 21922
rect 183154 4294 183250 4350
rect 183306 4294 183374 4350
rect 183430 4294 183498 4350
rect 183554 4294 183622 4350
rect 183678 4294 183774 4350
rect 183154 4226 183774 4294
rect 183154 4170 183250 4226
rect 183306 4170 183374 4226
rect 183430 4170 183498 4226
rect 183554 4170 183622 4226
rect 183678 4170 183774 4226
rect 183154 4102 183774 4170
rect 183154 4046 183250 4102
rect 183306 4046 183374 4102
rect 183430 4046 183498 4102
rect 183554 4046 183622 4102
rect 183678 4046 183774 4102
rect 183154 3978 183774 4046
rect 183154 3922 183250 3978
rect 183306 3922 183374 3978
rect 183430 3922 183498 3978
rect 183554 3922 183622 3978
rect 183678 3922 183774 3978
rect 183154 -160 183774 3922
rect 183154 -216 183250 -160
rect 183306 -216 183374 -160
rect 183430 -216 183498 -160
rect 183554 -216 183622 -160
rect 183678 -216 183774 -160
rect 183154 -284 183774 -216
rect 183154 -340 183250 -284
rect 183306 -340 183374 -284
rect 183430 -340 183498 -284
rect 183554 -340 183622 -284
rect 183678 -340 183774 -284
rect 183154 -408 183774 -340
rect 183154 -464 183250 -408
rect 183306 -464 183374 -408
rect 183430 -464 183498 -408
rect 183554 -464 183622 -408
rect 183678 -464 183774 -408
rect 183154 -532 183774 -464
rect 183154 -588 183250 -532
rect 183306 -588 183374 -532
rect 183430 -588 183498 -532
rect 183554 -588 183622 -532
rect 183678 -588 183774 -532
rect 183154 -1644 183774 -588
rect 186874 10350 187494 27922
rect 186874 10294 186970 10350
rect 187026 10294 187094 10350
rect 187150 10294 187218 10350
rect 187274 10294 187342 10350
rect 187398 10294 187494 10350
rect 186874 10226 187494 10294
rect 186874 10170 186970 10226
rect 187026 10170 187094 10226
rect 187150 10170 187218 10226
rect 187274 10170 187342 10226
rect 187398 10170 187494 10226
rect 186874 10102 187494 10170
rect 186874 10046 186970 10102
rect 187026 10046 187094 10102
rect 187150 10046 187218 10102
rect 187274 10046 187342 10102
rect 187398 10046 187494 10102
rect 186874 9978 187494 10046
rect 186874 9922 186970 9978
rect 187026 9922 187094 9978
rect 187150 9922 187218 9978
rect 187274 9922 187342 9978
rect 187398 9922 187494 9978
rect 186874 -1120 187494 9922
rect 186874 -1176 186970 -1120
rect 187026 -1176 187094 -1120
rect 187150 -1176 187218 -1120
rect 187274 -1176 187342 -1120
rect 187398 -1176 187494 -1120
rect 186874 -1244 187494 -1176
rect 186874 -1300 186970 -1244
rect 187026 -1300 187094 -1244
rect 187150 -1300 187218 -1244
rect 187274 -1300 187342 -1244
rect 187398 -1300 187494 -1244
rect 186874 -1368 187494 -1300
rect 186874 -1424 186970 -1368
rect 187026 -1424 187094 -1368
rect 187150 -1424 187218 -1368
rect 187274 -1424 187342 -1368
rect 187398 -1424 187494 -1368
rect 186874 -1492 187494 -1424
rect 186874 -1548 186970 -1492
rect 187026 -1548 187094 -1492
rect 187150 -1548 187218 -1492
rect 187274 -1548 187342 -1492
rect 187398 -1548 187494 -1492
rect 186874 -1644 187494 -1548
rect 201154 22350 201774 31350
rect 204874 28350 205494 31350
rect 209916 28532 209972 31500
rect 223580 31444 223636 32620
rect 223580 31378 223636 31388
rect 209916 28466 209972 28476
rect 215852 28532 215908 28542
rect 204874 28294 204970 28350
rect 205026 28294 205094 28350
rect 205150 28294 205218 28350
rect 205274 28294 205342 28350
rect 205398 28294 205494 28350
rect 204874 28226 205494 28294
rect 204874 28170 204970 28226
rect 205026 28170 205094 28226
rect 205150 28170 205218 28226
rect 205274 28170 205342 28226
rect 205398 28170 205494 28226
rect 204874 28102 205494 28170
rect 204874 28046 204970 28102
rect 205026 28046 205094 28102
rect 205150 28046 205218 28102
rect 205274 28046 205342 28102
rect 205398 28046 205494 28102
rect 204874 27978 205494 28046
rect 204874 27922 204970 27978
rect 205026 27922 205094 27978
rect 205150 27922 205218 27978
rect 205274 27922 205342 27978
rect 205398 27922 205494 27978
rect 203308 27658 203364 27668
rect 203308 27564 203364 27580
rect 201154 22294 201250 22350
rect 201306 22294 201374 22350
rect 201430 22294 201498 22350
rect 201554 22294 201622 22350
rect 201678 22294 201774 22350
rect 201154 22226 201774 22294
rect 201154 22170 201250 22226
rect 201306 22170 201374 22226
rect 201430 22170 201498 22226
rect 201554 22170 201622 22226
rect 201678 22170 201774 22226
rect 201154 22102 201774 22170
rect 201154 22046 201250 22102
rect 201306 22046 201374 22102
rect 201430 22046 201498 22102
rect 201554 22046 201622 22102
rect 201678 22046 201774 22102
rect 201154 21978 201774 22046
rect 201154 21922 201250 21978
rect 201306 21922 201374 21978
rect 201430 21922 201498 21978
rect 201554 21922 201622 21978
rect 201678 21922 201774 21978
rect 201154 4350 201774 21922
rect 201154 4294 201250 4350
rect 201306 4294 201374 4350
rect 201430 4294 201498 4350
rect 201554 4294 201622 4350
rect 201678 4294 201774 4350
rect 201154 4226 201774 4294
rect 201154 4170 201250 4226
rect 201306 4170 201374 4226
rect 201430 4170 201498 4226
rect 201554 4170 201622 4226
rect 201678 4170 201774 4226
rect 201154 4102 201774 4170
rect 201154 4046 201250 4102
rect 201306 4046 201374 4102
rect 201430 4046 201498 4102
rect 201554 4046 201622 4102
rect 201678 4046 201774 4102
rect 201154 3978 201774 4046
rect 201154 3922 201250 3978
rect 201306 3922 201374 3978
rect 201430 3922 201498 3978
rect 201554 3922 201622 3978
rect 201678 3922 201774 3978
rect 201154 -160 201774 3922
rect 201154 -216 201250 -160
rect 201306 -216 201374 -160
rect 201430 -216 201498 -160
rect 201554 -216 201622 -160
rect 201678 -216 201774 -160
rect 201154 -284 201774 -216
rect 201154 -340 201250 -284
rect 201306 -340 201374 -284
rect 201430 -340 201498 -284
rect 201554 -340 201622 -284
rect 201678 -340 201774 -284
rect 201154 -408 201774 -340
rect 201154 -464 201250 -408
rect 201306 -464 201374 -408
rect 201430 -464 201498 -408
rect 201554 -464 201622 -408
rect 201678 -464 201774 -408
rect 201154 -532 201774 -464
rect 201154 -588 201250 -532
rect 201306 -588 201374 -532
rect 201430 -588 201498 -532
rect 201554 -588 201622 -532
rect 201678 -588 201774 -532
rect 201154 -1644 201774 -588
rect 204874 10350 205494 27922
rect 215852 27658 215908 28476
rect 209356 26938 209412 26948
rect 209356 21588 209412 26882
rect 209356 21522 209412 21532
rect 215852 12740 215908 27602
rect 218428 27478 218484 27488
rect 218428 21252 218484 27422
rect 218428 21186 218484 21196
rect 219154 22350 219774 31350
rect 221564 29652 221620 29676
rect 219884 28532 219940 28542
rect 219884 27478 219940 28476
rect 219884 27412 219940 27422
rect 220108 28532 220164 28542
rect 219154 22294 219250 22350
rect 219306 22294 219374 22350
rect 219430 22294 219498 22350
rect 219554 22294 219622 22350
rect 219678 22294 219774 22350
rect 219154 22226 219774 22294
rect 219154 22170 219250 22226
rect 219306 22170 219374 22226
rect 219430 22170 219498 22226
rect 219554 22170 219622 22226
rect 219678 22170 219774 22226
rect 219154 22102 219774 22170
rect 219154 22046 219250 22102
rect 219306 22046 219374 22102
rect 219430 22046 219498 22102
rect 219554 22046 219622 22102
rect 219678 22046 219774 22102
rect 219154 21978 219774 22046
rect 219154 21922 219250 21978
rect 219306 21922 219374 21978
rect 219430 21922 219498 21978
rect 219554 21922 219622 21978
rect 219678 21922 219774 21978
rect 215852 12674 215908 12684
rect 204874 10294 204970 10350
rect 205026 10294 205094 10350
rect 205150 10294 205218 10350
rect 205274 10294 205342 10350
rect 205398 10294 205494 10350
rect 204874 10226 205494 10294
rect 204874 10170 204970 10226
rect 205026 10170 205094 10226
rect 205150 10170 205218 10226
rect 205274 10170 205342 10226
rect 205398 10170 205494 10226
rect 204874 10102 205494 10170
rect 204874 10046 204970 10102
rect 205026 10046 205094 10102
rect 205150 10046 205218 10102
rect 205274 10046 205342 10102
rect 205398 10046 205494 10102
rect 204874 9978 205494 10046
rect 204874 9922 204970 9978
rect 205026 9922 205094 9978
rect 205150 9922 205218 9978
rect 205274 9922 205342 9978
rect 205398 9922 205494 9978
rect 204874 -1120 205494 9922
rect 204874 -1176 204970 -1120
rect 205026 -1176 205094 -1120
rect 205150 -1176 205218 -1120
rect 205274 -1176 205342 -1120
rect 205398 -1176 205494 -1120
rect 204874 -1244 205494 -1176
rect 204874 -1300 204970 -1244
rect 205026 -1300 205094 -1244
rect 205150 -1300 205218 -1244
rect 205274 -1300 205342 -1244
rect 205398 -1300 205494 -1244
rect 204874 -1368 205494 -1300
rect 204874 -1424 204970 -1368
rect 205026 -1424 205094 -1368
rect 205150 -1424 205218 -1368
rect 205274 -1424 205342 -1368
rect 205398 -1424 205494 -1368
rect 204874 -1492 205494 -1424
rect 204874 -1548 204970 -1492
rect 205026 -1548 205094 -1492
rect 205150 -1548 205218 -1492
rect 205274 -1548 205342 -1492
rect 205398 -1548 205494 -1492
rect 204874 -1644 205494 -1548
rect 219154 4350 219774 21922
rect 220108 10948 220164 28476
rect 221564 28532 221620 29582
rect 221564 28466 221620 28476
rect 220108 10882 220164 10892
rect 222874 28350 223494 31350
rect 222874 28294 222970 28350
rect 223026 28294 223094 28350
rect 223150 28294 223218 28350
rect 223274 28294 223342 28350
rect 223398 28294 223494 28350
rect 222874 28226 223494 28294
rect 222874 28170 222970 28226
rect 223026 28170 223094 28226
rect 223150 28170 223218 28226
rect 223274 28170 223342 28226
rect 223398 28170 223494 28226
rect 222874 28102 223494 28170
rect 222874 28046 222970 28102
rect 223026 28046 223094 28102
rect 223150 28046 223218 28102
rect 223274 28046 223342 28102
rect 223398 28046 223494 28102
rect 222874 27978 223494 28046
rect 222874 27922 222970 27978
rect 223026 27922 223094 27978
rect 223150 27922 223218 27978
rect 223274 27922 223342 27978
rect 223398 27922 223494 27978
rect 219154 4294 219250 4350
rect 219306 4294 219374 4350
rect 219430 4294 219498 4350
rect 219554 4294 219622 4350
rect 219678 4294 219774 4350
rect 219154 4226 219774 4294
rect 219154 4170 219250 4226
rect 219306 4170 219374 4226
rect 219430 4170 219498 4226
rect 219554 4170 219622 4226
rect 219678 4170 219774 4226
rect 219154 4102 219774 4170
rect 219154 4046 219250 4102
rect 219306 4046 219374 4102
rect 219430 4046 219498 4102
rect 219554 4046 219622 4102
rect 219678 4046 219774 4102
rect 219154 3978 219774 4046
rect 219154 3922 219250 3978
rect 219306 3922 219374 3978
rect 219430 3922 219498 3978
rect 219554 3922 219622 3978
rect 219678 3922 219774 3978
rect 219154 -160 219774 3922
rect 219154 -216 219250 -160
rect 219306 -216 219374 -160
rect 219430 -216 219498 -160
rect 219554 -216 219622 -160
rect 219678 -216 219774 -160
rect 219154 -284 219774 -216
rect 219154 -340 219250 -284
rect 219306 -340 219374 -284
rect 219430 -340 219498 -284
rect 219554 -340 219622 -284
rect 219678 -340 219774 -284
rect 219154 -408 219774 -340
rect 219154 -464 219250 -408
rect 219306 -464 219374 -408
rect 219430 -464 219498 -408
rect 219554 -464 219622 -408
rect 219678 -464 219774 -408
rect 219154 -532 219774 -464
rect 219154 -588 219250 -532
rect 219306 -588 219374 -532
rect 219430 -588 219498 -532
rect 219554 -588 219622 -532
rect 219678 -588 219774 -532
rect 219154 -1644 219774 -588
rect 222874 10350 223494 27922
rect 222874 10294 222970 10350
rect 223026 10294 223094 10350
rect 223150 10294 223218 10350
rect 223274 10294 223342 10350
rect 223398 10294 223494 10350
rect 222874 10226 223494 10294
rect 222874 10170 222970 10226
rect 223026 10170 223094 10226
rect 223150 10170 223218 10226
rect 223274 10170 223342 10226
rect 223398 10170 223494 10226
rect 222874 10102 223494 10170
rect 222874 10046 222970 10102
rect 223026 10046 223094 10102
rect 223150 10046 223218 10102
rect 223274 10046 223342 10102
rect 223398 10046 223494 10102
rect 222874 9978 223494 10046
rect 222874 9922 222970 9978
rect 223026 9922 223094 9978
rect 223150 9922 223218 9978
rect 223274 9922 223342 9978
rect 223398 9922 223494 9978
rect 222874 -1120 223494 9922
rect 222874 -1176 222970 -1120
rect 223026 -1176 223094 -1120
rect 223150 -1176 223218 -1120
rect 223274 -1176 223342 -1120
rect 223398 -1176 223494 -1120
rect 222874 -1244 223494 -1176
rect 222874 -1300 222970 -1244
rect 223026 -1300 223094 -1244
rect 223150 -1300 223218 -1244
rect 223274 -1300 223342 -1244
rect 223398 -1300 223494 -1244
rect 222874 -1368 223494 -1300
rect 222874 -1424 222970 -1368
rect 223026 -1424 223094 -1368
rect 223150 -1424 223218 -1368
rect 223274 -1424 223342 -1368
rect 223398 -1424 223494 -1368
rect 222874 -1492 223494 -1424
rect 222874 -1548 222970 -1492
rect 223026 -1548 223094 -1492
rect 223150 -1548 223218 -1492
rect 223274 -1548 223342 -1492
rect 223398 -1548 223494 -1492
rect 222874 -1644 223494 -1548
rect 237154 22350 237774 31350
rect 238476 27636 238532 34442
rect 238476 27570 238532 27580
rect 240874 28350 241494 45922
rect 242956 49364 243012 49374
rect 241948 43316 242004 43326
rect 241948 36820 242004 43260
rect 241948 36754 242004 36764
rect 242956 36708 243012 49308
rect 242956 36642 243012 36652
rect 244412 29638 244468 205772
rect 246092 164164 246148 218652
rect 252812 214676 252868 214686
rect 251132 210644 251188 210654
rect 247772 188468 247828 188478
rect 246092 164098 246148 164108
rect 246204 174356 246260 174366
rect 244524 162260 244580 162270
rect 244524 132804 244580 162204
rect 246204 139524 246260 174300
rect 247772 147364 247828 188412
rect 249452 184436 249508 184446
rect 247772 147298 247828 147308
rect 247884 166292 247940 166302
rect 246204 139458 246260 139468
rect 247884 135044 247940 166236
rect 249452 145124 249508 184380
rect 251132 159684 251188 210588
rect 251132 159618 251188 159628
rect 251244 180404 251300 180414
rect 249452 145058 249508 145068
rect 249676 145348 249732 145358
rect 247884 134978 247940 134988
rect 248108 136052 248164 136062
rect 244524 132738 244580 132748
rect 244524 130004 244580 130014
rect 244524 114884 244580 129948
rect 244524 114818 244580 114828
rect 246092 123956 246148 123966
rect 246092 113428 246148 123900
rect 248108 121828 248164 135996
rect 249676 126084 249732 145292
rect 251244 142884 251300 180348
rect 252812 161924 252868 214620
rect 255154 202350 255774 219922
rect 255154 202294 255250 202350
rect 255306 202294 255374 202350
rect 255430 202294 255498 202350
rect 255554 202294 255622 202350
rect 255678 202294 255774 202350
rect 255154 202226 255774 202294
rect 255154 202170 255250 202226
rect 255306 202170 255374 202226
rect 255430 202170 255498 202226
rect 255554 202170 255622 202226
rect 255678 202170 255774 202226
rect 255154 202102 255774 202170
rect 255154 202046 255250 202102
rect 255306 202046 255374 202102
rect 255430 202046 255498 202102
rect 255554 202046 255622 202102
rect 255678 202046 255774 202102
rect 255154 201978 255774 202046
rect 255154 201922 255250 201978
rect 255306 201922 255374 201978
rect 255430 201922 255498 201978
rect 255554 201922 255622 201978
rect 255678 201922 255774 201978
rect 255154 184350 255774 201922
rect 258874 226350 259494 243922
rect 258874 226294 258970 226350
rect 259026 226294 259094 226350
rect 259150 226294 259218 226350
rect 259274 226294 259342 226350
rect 259398 226294 259494 226350
rect 258874 226226 259494 226294
rect 258874 226170 258970 226226
rect 259026 226170 259094 226226
rect 259150 226170 259218 226226
rect 259274 226170 259342 226226
rect 259398 226170 259494 226226
rect 258874 226102 259494 226170
rect 258874 226046 258970 226102
rect 259026 226046 259094 226102
rect 259150 226046 259218 226102
rect 259274 226046 259342 226102
rect 259398 226046 259494 226102
rect 258874 225978 259494 226046
rect 258874 225922 258970 225978
rect 259026 225922 259094 225978
rect 259150 225922 259218 225978
rect 259274 225922 259342 225978
rect 259398 225922 259494 225978
rect 258874 208350 259494 225922
rect 273154 597212 273774 598268
rect 273154 597156 273250 597212
rect 273306 597156 273374 597212
rect 273430 597156 273498 597212
rect 273554 597156 273622 597212
rect 273678 597156 273774 597212
rect 273154 597088 273774 597156
rect 273154 597032 273250 597088
rect 273306 597032 273374 597088
rect 273430 597032 273498 597088
rect 273554 597032 273622 597088
rect 273678 597032 273774 597088
rect 273154 596964 273774 597032
rect 273154 596908 273250 596964
rect 273306 596908 273374 596964
rect 273430 596908 273498 596964
rect 273554 596908 273622 596964
rect 273678 596908 273774 596964
rect 273154 596840 273774 596908
rect 273154 596784 273250 596840
rect 273306 596784 273374 596840
rect 273430 596784 273498 596840
rect 273554 596784 273622 596840
rect 273678 596784 273774 596840
rect 273154 580350 273774 596784
rect 273154 580294 273250 580350
rect 273306 580294 273374 580350
rect 273430 580294 273498 580350
rect 273554 580294 273622 580350
rect 273678 580294 273774 580350
rect 273154 580226 273774 580294
rect 273154 580170 273250 580226
rect 273306 580170 273374 580226
rect 273430 580170 273498 580226
rect 273554 580170 273622 580226
rect 273678 580170 273774 580226
rect 273154 580102 273774 580170
rect 273154 580046 273250 580102
rect 273306 580046 273374 580102
rect 273430 580046 273498 580102
rect 273554 580046 273622 580102
rect 273678 580046 273774 580102
rect 273154 579978 273774 580046
rect 273154 579922 273250 579978
rect 273306 579922 273374 579978
rect 273430 579922 273498 579978
rect 273554 579922 273622 579978
rect 273678 579922 273774 579978
rect 273154 562350 273774 579922
rect 273154 562294 273250 562350
rect 273306 562294 273374 562350
rect 273430 562294 273498 562350
rect 273554 562294 273622 562350
rect 273678 562294 273774 562350
rect 273154 562226 273774 562294
rect 273154 562170 273250 562226
rect 273306 562170 273374 562226
rect 273430 562170 273498 562226
rect 273554 562170 273622 562226
rect 273678 562170 273774 562226
rect 273154 562102 273774 562170
rect 273154 562046 273250 562102
rect 273306 562046 273374 562102
rect 273430 562046 273498 562102
rect 273554 562046 273622 562102
rect 273678 562046 273774 562102
rect 273154 561978 273774 562046
rect 273154 561922 273250 561978
rect 273306 561922 273374 561978
rect 273430 561922 273498 561978
rect 273554 561922 273622 561978
rect 273678 561922 273774 561978
rect 273154 544350 273774 561922
rect 273154 544294 273250 544350
rect 273306 544294 273374 544350
rect 273430 544294 273498 544350
rect 273554 544294 273622 544350
rect 273678 544294 273774 544350
rect 273154 544226 273774 544294
rect 273154 544170 273250 544226
rect 273306 544170 273374 544226
rect 273430 544170 273498 544226
rect 273554 544170 273622 544226
rect 273678 544170 273774 544226
rect 273154 544102 273774 544170
rect 273154 544046 273250 544102
rect 273306 544046 273374 544102
rect 273430 544046 273498 544102
rect 273554 544046 273622 544102
rect 273678 544046 273774 544102
rect 273154 543978 273774 544046
rect 273154 543922 273250 543978
rect 273306 543922 273374 543978
rect 273430 543922 273498 543978
rect 273554 543922 273622 543978
rect 273678 543922 273774 543978
rect 273154 526350 273774 543922
rect 273154 526294 273250 526350
rect 273306 526294 273374 526350
rect 273430 526294 273498 526350
rect 273554 526294 273622 526350
rect 273678 526294 273774 526350
rect 273154 526226 273774 526294
rect 273154 526170 273250 526226
rect 273306 526170 273374 526226
rect 273430 526170 273498 526226
rect 273554 526170 273622 526226
rect 273678 526170 273774 526226
rect 273154 526102 273774 526170
rect 273154 526046 273250 526102
rect 273306 526046 273374 526102
rect 273430 526046 273498 526102
rect 273554 526046 273622 526102
rect 273678 526046 273774 526102
rect 273154 525978 273774 526046
rect 273154 525922 273250 525978
rect 273306 525922 273374 525978
rect 273430 525922 273498 525978
rect 273554 525922 273622 525978
rect 273678 525922 273774 525978
rect 273154 508350 273774 525922
rect 273154 508294 273250 508350
rect 273306 508294 273374 508350
rect 273430 508294 273498 508350
rect 273554 508294 273622 508350
rect 273678 508294 273774 508350
rect 273154 508226 273774 508294
rect 273154 508170 273250 508226
rect 273306 508170 273374 508226
rect 273430 508170 273498 508226
rect 273554 508170 273622 508226
rect 273678 508170 273774 508226
rect 273154 508102 273774 508170
rect 273154 508046 273250 508102
rect 273306 508046 273374 508102
rect 273430 508046 273498 508102
rect 273554 508046 273622 508102
rect 273678 508046 273774 508102
rect 273154 507978 273774 508046
rect 273154 507922 273250 507978
rect 273306 507922 273374 507978
rect 273430 507922 273498 507978
rect 273554 507922 273622 507978
rect 273678 507922 273774 507978
rect 273154 490350 273774 507922
rect 273154 490294 273250 490350
rect 273306 490294 273374 490350
rect 273430 490294 273498 490350
rect 273554 490294 273622 490350
rect 273678 490294 273774 490350
rect 273154 490226 273774 490294
rect 273154 490170 273250 490226
rect 273306 490170 273374 490226
rect 273430 490170 273498 490226
rect 273554 490170 273622 490226
rect 273678 490170 273774 490226
rect 273154 490102 273774 490170
rect 273154 490046 273250 490102
rect 273306 490046 273374 490102
rect 273430 490046 273498 490102
rect 273554 490046 273622 490102
rect 273678 490046 273774 490102
rect 273154 489978 273774 490046
rect 273154 489922 273250 489978
rect 273306 489922 273374 489978
rect 273430 489922 273498 489978
rect 273554 489922 273622 489978
rect 273678 489922 273774 489978
rect 273154 472350 273774 489922
rect 273154 472294 273250 472350
rect 273306 472294 273374 472350
rect 273430 472294 273498 472350
rect 273554 472294 273622 472350
rect 273678 472294 273774 472350
rect 273154 472226 273774 472294
rect 273154 472170 273250 472226
rect 273306 472170 273374 472226
rect 273430 472170 273498 472226
rect 273554 472170 273622 472226
rect 273678 472170 273774 472226
rect 273154 472102 273774 472170
rect 273154 472046 273250 472102
rect 273306 472046 273374 472102
rect 273430 472046 273498 472102
rect 273554 472046 273622 472102
rect 273678 472046 273774 472102
rect 273154 471978 273774 472046
rect 273154 471922 273250 471978
rect 273306 471922 273374 471978
rect 273430 471922 273498 471978
rect 273554 471922 273622 471978
rect 273678 471922 273774 471978
rect 273154 454350 273774 471922
rect 273154 454294 273250 454350
rect 273306 454294 273374 454350
rect 273430 454294 273498 454350
rect 273554 454294 273622 454350
rect 273678 454294 273774 454350
rect 273154 454226 273774 454294
rect 273154 454170 273250 454226
rect 273306 454170 273374 454226
rect 273430 454170 273498 454226
rect 273554 454170 273622 454226
rect 273678 454170 273774 454226
rect 273154 454102 273774 454170
rect 273154 454046 273250 454102
rect 273306 454046 273374 454102
rect 273430 454046 273498 454102
rect 273554 454046 273622 454102
rect 273678 454046 273774 454102
rect 273154 453978 273774 454046
rect 273154 453922 273250 453978
rect 273306 453922 273374 453978
rect 273430 453922 273498 453978
rect 273554 453922 273622 453978
rect 273678 453922 273774 453978
rect 273154 436350 273774 453922
rect 273154 436294 273250 436350
rect 273306 436294 273374 436350
rect 273430 436294 273498 436350
rect 273554 436294 273622 436350
rect 273678 436294 273774 436350
rect 273154 436226 273774 436294
rect 273154 436170 273250 436226
rect 273306 436170 273374 436226
rect 273430 436170 273498 436226
rect 273554 436170 273622 436226
rect 273678 436170 273774 436226
rect 273154 436102 273774 436170
rect 273154 436046 273250 436102
rect 273306 436046 273374 436102
rect 273430 436046 273498 436102
rect 273554 436046 273622 436102
rect 273678 436046 273774 436102
rect 273154 435978 273774 436046
rect 273154 435922 273250 435978
rect 273306 435922 273374 435978
rect 273430 435922 273498 435978
rect 273554 435922 273622 435978
rect 273678 435922 273774 435978
rect 273154 418350 273774 435922
rect 273154 418294 273250 418350
rect 273306 418294 273374 418350
rect 273430 418294 273498 418350
rect 273554 418294 273622 418350
rect 273678 418294 273774 418350
rect 273154 418226 273774 418294
rect 273154 418170 273250 418226
rect 273306 418170 273374 418226
rect 273430 418170 273498 418226
rect 273554 418170 273622 418226
rect 273678 418170 273774 418226
rect 273154 418102 273774 418170
rect 273154 418046 273250 418102
rect 273306 418046 273374 418102
rect 273430 418046 273498 418102
rect 273554 418046 273622 418102
rect 273678 418046 273774 418102
rect 273154 417978 273774 418046
rect 273154 417922 273250 417978
rect 273306 417922 273374 417978
rect 273430 417922 273498 417978
rect 273554 417922 273622 417978
rect 273678 417922 273774 417978
rect 273154 400350 273774 417922
rect 273154 400294 273250 400350
rect 273306 400294 273374 400350
rect 273430 400294 273498 400350
rect 273554 400294 273622 400350
rect 273678 400294 273774 400350
rect 273154 400226 273774 400294
rect 273154 400170 273250 400226
rect 273306 400170 273374 400226
rect 273430 400170 273498 400226
rect 273554 400170 273622 400226
rect 273678 400170 273774 400226
rect 273154 400102 273774 400170
rect 273154 400046 273250 400102
rect 273306 400046 273374 400102
rect 273430 400046 273498 400102
rect 273554 400046 273622 400102
rect 273678 400046 273774 400102
rect 273154 399978 273774 400046
rect 273154 399922 273250 399978
rect 273306 399922 273374 399978
rect 273430 399922 273498 399978
rect 273554 399922 273622 399978
rect 273678 399922 273774 399978
rect 273154 382350 273774 399922
rect 273154 382294 273250 382350
rect 273306 382294 273374 382350
rect 273430 382294 273498 382350
rect 273554 382294 273622 382350
rect 273678 382294 273774 382350
rect 273154 382226 273774 382294
rect 273154 382170 273250 382226
rect 273306 382170 273374 382226
rect 273430 382170 273498 382226
rect 273554 382170 273622 382226
rect 273678 382170 273774 382226
rect 273154 382102 273774 382170
rect 273154 382046 273250 382102
rect 273306 382046 273374 382102
rect 273430 382046 273498 382102
rect 273554 382046 273622 382102
rect 273678 382046 273774 382102
rect 273154 381978 273774 382046
rect 273154 381922 273250 381978
rect 273306 381922 273374 381978
rect 273430 381922 273498 381978
rect 273554 381922 273622 381978
rect 273678 381922 273774 381978
rect 273154 364350 273774 381922
rect 273154 364294 273250 364350
rect 273306 364294 273374 364350
rect 273430 364294 273498 364350
rect 273554 364294 273622 364350
rect 273678 364294 273774 364350
rect 273154 364226 273774 364294
rect 273154 364170 273250 364226
rect 273306 364170 273374 364226
rect 273430 364170 273498 364226
rect 273554 364170 273622 364226
rect 273678 364170 273774 364226
rect 273154 364102 273774 364170
rect 273154 364046 273250 364102
rect 273306 364046 273374 364102
rect 273430 364046 273498 364102
rect 273554 364046 273622 364102
rect 273678 364046 273774 364102
rect 273154 363978 273774 364046
rect 273154 363922 273250 363978
rect 273306 363922 273374 363978
rect 273430 363922 273498 363978
rect 273554 363922 273622 363978
rect 273678 363922 273774 363978
rect 273154 346350 273774 363922
rect 273154 346294 273250 346350
rect 273306 346294 273374 346350
rect 273430 346294 273498 346350
rect 273554 346294 273622 346350
rect 273678 346294 273774 346350
rect 273154 346226 273774 346294
rect 273154 346170 273250 346226
rect 273306 346170 273374 346226
rect 273430 346170 273498 346226
rect 273554 346170 273622 346226
rect 273678 346170 273774 346226
rect 273154 346102 273774 346170
rect 273154 346046 273250 346102
rect 273306 346046 273374 346102
rect 273430 346046 273498 346102
rect 273554 346046 273622 346102
rect 273678 346046 273774 346102
rect 273154 345978 273774 346046
rect 273154 345922 273250 345978
rect 273306 345922 273374 345978
rect 273430 345922 273498 345978
rect 273554 345922 273622 345978
rect 273678 345922 273774 345978
rect 273154 328350 273774 345922
rect 273154 328294 273250 328350
rect 273306 328294 273374 328350
rect 273430 328294 273498 328350
rect 273554 328294 273622 328350
rect 273678 328294 273774 328350
rect 273154 328226 273774 328294
rect 273154 328170 273250 328226
rect 273306 328170 273374 328226
rect 273430 328170 273498 328226
rect 273554 328170 273622 328226
rect 273678 328170 273774 328226
rect 273154 328102 273774 328170
rect 273154 328046 273250 328102
rect 273306 328046 273374 328102
rect 273430 328046 273498 328102
rect 273554 328046 273622 328102
rect 273678 328046 273774 328102
rect 273154 327978 273774 328046
rect 273154 327922 273250 327978
rect 273306 327922 273374 327978
rect 273430 327922 273498 327978
rect 273554 327922 273622 327978
rect 273678 327922 273774 327978
rect 273154 310350 273774 327922
rect 273154 310294 273250 310350
rect 273306 310294 273374 310350
rect 273430 310294 273498 310350
rect 273554 310294 273622 310350
rect 273678 310294 273774 310350
rect 273154 310226 273774 310294
rect 273154 310170 273250 310226
rect 273306 310170 273374 310226
rect 273430 310170 273498 310226
rect 273554 310170 273622 310226
rect 273678 310170 273774 310226
rect 273154 310102 273774 310170
rect 273154 310046 273250 310102
rect 273306 310046 273374 310102
rect 273430 310046 273498 310102
rect 273554 310046 273622 310102
rect 273678 310046 273774 310102
rect 273154 309978 273774 310046
rect 273154 309922 273250 309978
rect 273306 309922 273374 309978
rect 273430 309922 273498 309978
rect 273554 309922 273622 309978
rect 273678 309922 273774 309978
rect 273154 292350 273774 309922
rect 273154 292294 273250 292350
rect 273306 292294 273374 292350
rect 273430 292294 273498 292350
rect 273554 292294 273622 292350
rect 273678 292294 273774 292350
rect 273154 292226 273774 292294
rect 273154 292170 273250 292226
rect 273306 292170 273374 292226
rect 273430 292170 273498 292226
rect 273554 292170 273622 292226
rect 273678 292170 273774 292226
rect 273154 292102 273774 292170
rect 273154 292046 273250 292102
rect 273306 292046 273374 292102
rect 273430 292046 273498 292102
rect 273554 292046 273622 292102
rect 273678 292046 273774 292102
rect 273154 291978 273774 292046
rect 273154 291922 273250 291978
rect 273306 291922 273374 291978
rect 273430 291922 273498 291978
rect 273554 291922 273622 291978
rect 273678 291922 273774 291978
rect 273154 274350 273774 291922
rect 273154 274294 273250 274350
rect 273306 274294 273374 274350
rect 273430 274294 273498 274350
rect 273554 274294 273622 274350
rect 273678 274294 273774 274350
rect 273154 274226 273774 274294
rect 273154 274170 273250 274226
rect 273306 274170 273374 274226
rect 273430 274170 273498 274226
rect 273554 274170 273622 274226
rect 273678 274170 273774 274226
rect 273154 274102 273774 274170
rect 273154 274046 273250 274102
rect 273306 274046 273374 274102
rect 273430 274046 273498 274102
rect 273554 274046 273622 274102
rect 273678 274046 273774 274102
rect 273154 273978 273774 274046
rect 273154 273922 273250 273978
rect 273306 273922 273374 273978
rect 273430 273922 273498 273978
rect 273554 273922 273622 273978
rect 273678 273922 273774 273978
rect 273154 256350 273774 273922
rect 273154 256294 273250 256350
rect 273306 256294 273374 256350
rect 273430 256294 273498 256350
rect 273554 256294 273622 256350
rect 273678 256294 273774 256350
rect 273154 256226 273774 256294
rect 273154 256170 273250 256226
rect 273306 256170 273374 256226
rect 273430 256170 273498 256226
rect 273554 256170 273622 256226
rect 273678 256170 273774 256226
rect 273154 256102 273774 256170
rect 273154 256046 273250 256102
rect 273306 256046 273374 256102
rect 273430 256046 273498 256102
rect 273554 256046 273622 256102
rect 273678 256046 273774 256102
rect 273154 255978 273774 256046
rect 273154 255922 273250 255978
rect 273306 255922 273374 255978
rect 273430 255922 273498 255978
rect 273554 255922 273622 255978
rect 273678 255922 273774 255978
rect 273154 238350 273774 255922
rect 273154 238294 273250 238350
rect 273306 238294 273374 238350
rect 273430 238294 273498 238350
rect 273554 238294 273622 238350
rect 273678 238294 273774 238350
rect 273154 238226 273774 238294
rect 273154 238170 273250 238226
rect 273306 238170 273374 238226
rect 273430 238170 273498 238226
rect 273554 238170 273622 238226
rect 273678 238170 273774 238226
rect 273154 238102 273774 238170
rect 273154 238046 273250 238102
rect 273306 238046 273374 238102
rect 273430 238046 273498 238102
rect 273554 238046 273622 238102
rect 273678 238046 273774 238102
rect 273154 237978 273774 238046
rect 273154 237922 273250 237978
rect 273306 237922 273374 237978
rect 273430 237922 273498 237978
rect 273554 237922 273622 237978
rect 273678 237922 273774 237978
rect 273154 220350 273774 237922
rect 273154 220294 273250 220350
rect 273306 220294 273374 220350
rect 273430 220294 273498 220350
rect 273554 220294 273622 220350
rect 273678 220294 273774 220350
rect 273154 220226 273774 220294
rect 273154 220170 273250 220226
rect 273306 220170 273374 220226
rect 273430 220170 273498 220226
rect 273554 220170 273622 220226
rect 273678 220170 273774 220226
rect 273154 220102 273774 220170
rect 273154 220046 273250 220102
rect 273306 220046 273374 220102
rect 273430 220046 273498 220102
rect 273554 220046 273622 220102
rect 273678 220046 273774 220102
rect 273154 219978 273774 220046
rect 273154 219922 273250 219978
rect 273306 219922 273374 219978
rect 273430 219922 273498 219978
rect 273554 219922 273622 219978
rect 273678 219922 273774 219978
rect 258874 208294 258970 208350
rect 259026 208294 259094 208350
rect 259150 208294 259218 208350
rect 259274 208294 259342 208350
rect 259398 208294 259494 208350
rect 258874 208226 259494 208294
rect 258874 208170 258970 208226
rect 259026 208170 259094 208226
rect 259150 208170 259218 208226
rect 259274 208170 259342 208226
rect 259398 208170 259494 208226
rect 258874 208102 259494 208170
rect 258874 208046 258970 208102
rect 259026 208046 259094 208102
rect 259150 208046 259218 208102
rect 259274 208046 259342 208102
rect 259398 208046 259494 208102
rect 258874 207978 259494 208046
rect 258874 207922 258970 207978
rect 259026 207922 259094 207978
rect 259150 207922 259218 207978
rect 259274 207922 259342 207978
rect 259398 207922 259494 207978
rect 255154 184294 255250 184350
rect 255306 184294 255374 184350
rect 255430 184294 255498 184350
rect 255554 184294 255622 184350
rect 255678 184294 255774 184350
rect 255154 184226 255774 184294
rect 255154 184170 255250 184226
rect 255306 184170 255374 184226
rect 255430 184170 255498 184226
rect 255554 184170 255622 184226
rect 255678 184170 255774 184226
rect 255154 184102 255774 184170
rect 255154 184046 255250 184102
rect 255306 184046 255374 184102
rect 255430 184046 255498 184102
rect 255554 184046 255622 184102
rect 255678 184046 255774 184102
rect 255154 183978 255774 184046
rect 255154 183922 255250 183978
rect 255306 183922 255374 183978
rect 255430 183922 255498 183978
rect 255554 183922 255622 183978
rect 255678 183922 255774 183978
rect 252812 161858 252868 161868
rect 252924 178388 252980 178398
rect 251244 142818 251300 142828
rect 252924 141764 252980 178332
rect 252924 141698 252980 141708
rect 255154 166350 255774 183922
rect 255154 166294 255250 166350
rect 255306 166294 255374 166350
rect 255430 166294 255498 166350
rect 255554 166294 255622 166350
rect 255678 166294 255774 166350
rect 255154 166226 255774 166294
rect 255154 166170 255250 166226
rect 255306 166170 255374 166226
rect 255430 166170 255498 166226
rect 255554 166170 255622 166226
rect 255678 166170 255774 166226
rect 255154 166102 255774 166170
rect 255154 166046 255250 166102
rect 255306 166046 255374 166102
rect 255430 166046 255498 166102
rect 255554 166046 255622 166102
rect 255678 166046 255774 166102
rect 255154 165978 255774 166046
rect 255154 165922 255250 165978
rect 255306 165922 255374 165978
rect 255430 165922 255498 165978
rect 255554 165922 255622 165978
rect 255678 165922 255774 165978
rect 255154 148350 255774 165922
rect 257852 190484 257908 190494
rect 257852 148484 257908 190428
rect 258874 190350 259494 207922
rect 266252 216692 266308 216702
rect 264572 200564 264628 200574
rect 258874 190294 258970 190350
rect 259026 190294 259094 190350
rect 259150 190294 259218 190350
rect 259274 190294 259342 190350
rect 259398 190294 259494 190350
rect 258874 190226 259494 190294
rect 258874 190170 258970 190226
rect 259026 190170 259094 190226
rect 259150 190170 259218 190226
rect 259274 190170 259342 190226
rect 259398 190170 259494 190226
rect 258874 190102 259494 190170
rect 258874 190046 258970 190102
rect 259026 190046 259094 190102
rect 259150 190046 259218 190102
rect 259274 190046 259342 190102
rect 259398 190046 259494 190102
rect 258874 189978 259494 190046
rect 258874 189922 258970 189978
rect 259026 189922 259094 189978
rect 259150 189922 259218 189978
rect 259274 189922 259342 189978
rect 259398 189922 259494 189978
rect 258874 172350 259494 189922
rect 258874 172294 258970 172350
rect 259026 172294 259094 172350
rect 259150 172294 259218 172350
rect 259274 172294 259342 172350
rect 259398 172294 259494 172350
rect 258874 172226 259494 172294
rect 258874 172170 258970 172226
rect 259026 172170 259094 172226
rect 259150 172170 259218 172226
rect 259274 172170 259342 172226
rect 259398 172170 259494 172226
rect 258874 172102 259494 172170
rect 258874 172046 258970 172102
rect 259026 172046 259094 172102
rect 259150 172046 259218 172102
rect 259274 172046 259342 172102
rect 259398 172046 259494 172102
rect 258874 171978 259494 172046
rect 258874 171922 258970 171978
rect 259026 171922 259094 171978
rect 259150 171922 259218 171978
rect 259274 171922 259342 171978
rect 259398 171922 259494 171978
rect 257852 148418 257908 148428
rect 257964 158228 258020 158238
rect 255154 148294 255250 148350
rect 255306 148294 255374 148350
rect 255430 148294 255498 148350
rect 255554 148294 255622 148350
rect 255678 148294 255774 148350
rect 255154 148226 255774 148294
rect 255154 148170 255250 148226
rect 255306 148170 255374 148226
rect 255430 148170 255498 148226
rect 255554 148170 255622 148226
rect 255678 148170 255774 148226
rect 255154 148102 255774 148170
rect 255154 148046 255250 148102
rect 255306 148046 255374 148102
rect 255430 148046 255498 148102
rect 255554 148046 255622 148102
rect 255678 148046 255774 148102
rect 255154 147978 255774 148046
rect 255154 147922 255250 147978
rect 255306 147922 255374 147978
rect 255430 147922 255498 147978
rect 255554 147922 255622 147978
rect 255678 147922 255774 147978
rect 249676 126018 249732 126028
rect 252812 134036 252868 134046
rect 248108 121762 248164 121772
rect 252812 117124 252868 133980
rect 252812 117058 252868 117068
rect 255154 130350 255774 147922
rect 257964 131908 258020 158172
rect 258874 154350 259494 171922
rect 258874 154294 258970 154350
rect 259026 154294 259094 154350
rect 259150 154294 259218 154350
rect 259274 154294 259342 154350
rect 259398 154294 259494 154350
rect 258874 154226 259494 154294
rect 258874 154170 258970 154226
rect 259026 154170 259094 154226
rect 259150 154170 259218 154226
rect 259274 154170 259342 154226
rect 259398 154170 259494 154226
rect 258874 154102 259494 154170
rect 258874 154046 258970 154102
rect 259026 154046 259094 154102
rect 259150 154046 259218 154102
rect 259274 154046 259342 154102
rect 259398 154046 259494 154102
rect 258874 153978 259494 154046
rect 258874 153922 258970 153978
rect 259026 153922 259094 153978
rect 259150 153922 259218 153978
rect 259274 153922 259342 153978
rect 259398 153922 259494 153978
rect 258874 136350 259494 153922
rect 261212 196532 261268 196542
rect 261212 151844 261268 196476
rect 262892 192500 262948 192510
rect 261212 151778 261268 151788
rect 261324 168308 261380 168318
rect 261324 138628 261380 168252
rect 262892 149604 262948 192444
rect 262892 149538 262948 149548
rect 263004 164276 263060 164286
rect 261324 138562 261380 138572
rect 258874 136294 258970 136350
rect 259026 136294 259094 136350
rect 259150 136294 259218 136350
rect 259274 136294 259342 136350
rect 259398 136294 259494 136350
rect 258874 136226 259494 136294
rect 258874 136170 258970 136226
rect 259026 136170 259094 136226
rect 259150 136170 259218 136226
rect 259274 136170 259342 136226
rect 259398 136170 259494 136226
rect 258874 136102 259494 136170
rect 258874 136046 258970 136102
rect 259026 136046 259094 136102
rect 259150 136046 259218 136102
rect 259274 136046 259342 136102
rect 259398 136046 259494 136102
rect 258874 135978 259494 136046
rect 258874 135922 258970 135978
rect 259026 135922 259094 135978
rect 259150 135922 259218 135978
rect 259274 135922 259342 135978
rect 259398 135922 259494 135978
rect 257964 131842 258020 131852
rect 258188 132020 258244 132030
rect 255154 130294 255250 130350
rect 255306 130294 255374 130350
rect 255430 130294 255498 130350
rect 255554 130294 255622 130350
rect 255678 130294 255774 130350
rect 255154 130226 255774 130294
rect 255154 130170 255250 130226
rect 255306 130170 255374 130226
rect 255430 130170 255498 130226
rect 255554 130170 255622 130226
rect 255678 130170 255774 130226
rect 255154 130102 255774 130170
rect 255154 130046 255250 130102
rect 255306 130046 255374 130102
rect 255430 130046 255498 130102
rect 255554 130046 255622 130102
rect 255678 130046 255774 130102
rect 255154 129978 255774 130046
rect 255154 129922 255250 129978
rect 255306 129922 255374 129978
rect 255430 129922 255498 129978
rect 255554 129922 255622 129978
rect 255678 129922 255774 129978
rect 246092 113362 246148 113372
rect 255154 112350 255774 129922
rect 258188 116004 258244 131964
rect 258188 115938 258244 115948
rect 258874 118350 259494 135922
rect 263004 133924 263060 164220
rect 264572 155428 264628 200508
rect 264572 155362 264628 155372
rect 264684 182420 264740 182430
rect 263004 133858 263060 133868
rect 264572 152180 264628 152190
rect 264572 127204 264628 152124
rect 264684 144004 264740 182364
rect 266252 163044 266308 216636
rect 273154 202350 273774 219922
rect 276874 598172 277494 598268
rect 276874 598116 276970 598172
rect 277026 598116 277094 598172
rect 277150 598116 277218 598172
rect 277274 598116 277342 598172
rect 277398 598116 277494 598172
rect 276874 598048 277494 598116
rect 276874 597992 276970 598048
rect 277026 597992 277094 598048
rect 277150 597992 277218 598048
rect 277274 597992 277342 598048
rect 277398 597992 277494 598048
rect 276874 597924 277494 597992
rect 276874 597868 276970 597924
rect 277026 597868 277094 597924
rect 277150 597868 277218 597924
rect 277274 597868 277342 597924
rect 277398 597868 277494 597924
rect 276874 597800 277494 597868
rect 276874 597744 276970 597800
rect 277026 597744 277094 597800
rect 277150 597744 277218 597800
rect 277274 597744 277342 597800
rect 277398 597744 277494 597800
rect 276874 586350 277494 597744
rect 276874 586294 276970 586350
rect 277026 586294 277094 586350
rect 277150 586294 277218 586350
rect 277274 586294 277342 586350
rect 277398 586294 277494 586350
rect 276874 586226 277494 586294
rect 276874 586170 276970 586226
rect 277026 586170 277094 586226
rect 277150 586170 277218 586226
rect 277274 586170 277342 586226
rect 277398 586170 277494 586226
rect 276874 586102 277494 586170
rect 276874 586046 276970 586102
rect 277026 586046 277094 586102
rect 277150 586046 277218 586102
rect 277274 586046 277342 586102
rect 277398 586046 277494 586102
rect 276874 585978 277494 586046
rect 276874 585922 276970 585978
rect 277026 585922 277094 585978
rect 277150 585922 277218 585978
rect 277274 585922 277342 585978
rect 277398 585922 277494 585978
rect 276874 568350 277494 585922
rect 276874 568294 276970 568350
rect 277026 568294 277094 568350
rect 277150 568294 277218 568350
rect 277274 568294 277342 568350
rect 277398 568294 277494 568350
rect 276874 568226 277494 568294
rect 276874 568170 276970 568226
rect 277026 568170 277094 568226
rect 277150 568170 277218 568226
rect 277274 568170 277342 568226
rect 277398 568170 277494 568226
rect 276874 568102 277494 568170
rect 276874 568046 276970 568102
rect 277026 568046 277094 568102
rect 277150 568046 277218 568102
rect 277274 568046 277342 568102
rect 277398 568046 277494 568102
rect 276874 567978 277494 568046
rect 276874 567922 276970 567978
rect 277026 567922 277094 567978
rect 277150 567922 277218 567978
rect 277274 567922 277342 567978
rect 277398 567922 277494 567978
rect 276874 550350 277494 567922
rect 276874 550294 276970 550350
rect 277026 550294 277094 550350
rect 277150 550294 277218 550350
rect 277274 550294 277342 550350
rect 277398 550294 277494 550350
rect 276874 550226 277494 550294
rect 276874 550170 276970 550226
rect 277026 550170 277094 550226
rect 277150 550170 277218 550226
rect 277274 550170 277342 550226
rect 277398 550170 277494 550226
rect 276874 550102 277494 550170
rect 276874 550046 276970 550102
rect 277026 550046 277094 550102
rect 277150 550046 277218 550102
rect 277274 550046 277342 550102
rect 277398 550046 277494 550102
rect 276874 549978 277494 550046
rect 276874 549922 276970 549978
rect 277026 549922 277094 549978
rect 277150 549922 277218 549978
rect 277274 549922 277342 549978
rect 277398 549922 277494 549978
rect 276874 532350 277494 549922
rect 276874 532294 276970 532350
rect 277026 532294 277094 532350
rect 277150 532294 277218 532350
rect 277274 532294 277342 532350
rect 277398 532294 277494 532350
rect 276874 532226 277494 532294
rect 276874 532170 276970 532226
rect 277026 532170 277094 532226
rect 277150 532170 277218 532226
rect 277274 532170 277342 532226
rect 277398 532170 277494 532226
rect 276874 532102 277494 532170
rect 276874 532046 276970 532102
rect 277026 532046 277094 532102
rect 277150 532046 277218 532102
rect 277274 532046 277342 532102
rect 277398 532046 277494 532102
rect 276874 531978 277494 532046
rect 276874 531922 276970 531978
rect 277026 531922 277094 531978
rect 277150 531922 277218 531978
rect 277274 531922 277342 531978
rect 277398 531922 277494 531978
rect 276874 514350 277494 531922
rect 276874 514294 276970 514350
rect 277026 514294 277094 514350
rect 277150 514294 277218 514350
rect 277274 514294 277342 514350
rect 277398 514294 277494 514350
rect 276874 514226 277494 514294
rect 276874 514170 276970 514226
rect 277026 514170 277094 514226
rect 277150 514170 277218 514226
rect 277274 514170 277342 514226
rect 277398 514170 277494 514226
rect 276874 514102 277494 514170
rect 276874 514046 276970 514102
rect 277026 514046 277094 514102
rect 277150 514046 277218 514102
rect 277274 514046 277342 514102
rect 277398 514046 277494 514102
rect 276874 513978 277494 514046
rect 276874 513922 276970 513978
rect 277026 513922 277094 513978
rect 277150 513922 277218 513978
rect 277274 513922 277342 513978
rect 277398 513922 277494 513978
rect 276874 496350 277494 513922
rect 276874 496294 276970 496350
rect 277026 496294 277094 496350
rect 277150 496294 277218 496350
rect 277274 496294 277342 496350
rect 277398 496294 277494 496350
rect 276874 496226 277494 496294
rect 276874 496170 276970 496226
rect 277026 496170 277094 496226
rect 277150 496170 277218 496226
rect 277274 496170 277342 496226
rect 277398 496170 277494 496226
rect 276874 496102 277494 496170
rect 276874 496046 276970 496102
rect 277026 496046 277094 496102
rect 277150 496046 277218 496102
rect 277274 496046 277342 496102
rect 277398 496046 277494 496102
rect 276874 495978 277494 496046
rect 276874 495922 276970 495978
rect 277026 495922 277094 495978
rect 277150 495922 277218 495978
rect 277274 495922 277342 495978
rect 277398 495922 277494 495978
rect 276874 478350 277494 495922
rect 276874 478294 276970 478350
rect 277026 478294 277094 478350
rect 277150 478294 277218 478350
rect 277274 478294 277342 478350
rect 277398 478294 277494 478350
rect 276874 478226 277494 478294
rect 276874 478170 276970 478226
rect 277026 478170 277094 478226
rect 277150 478170 277218 478226
rect 277274 478170 277342 478226
rect 277398 478170 277494 478226
rect 276874 478102 277494 478170
rect 276874 478046 276970 478102
rect 277026 478046 277094 478102
rect 277150 478046 277218 478102
rect 277274 478046 277342 478102
rect 277398 478046 277494 478102
rect 276874 477978 277494 478046
rect 276874 477922 276970 477978
rect 277026 477922 277094 477978
rect 277150 477922 277218 477978
rect 277274 477922 277342 477978
rect 277398 477922 277494 477978
rect 276874 460350 277494 477922
rect 276874 460294 276970 460350
rect 277026 460294 277094 460350
rect 277150 460294 277218 460350
rect 277274 460294 277342 460350
rect 277398 460294 277494 460350
rect 276874 460226 277494 460294
rect 276874 460170 276970 460226
rect 277026 460170 277094 460226
rect 277150 460170 277218 460226
rect 277274 460170 277342 460226
rect 277398 460170 277494 460226
rect 276874 460102 277494 460170
rect 276874 460046 276970 460102
rect 277026 460046 277094 460102
rect 277150 460046 277218 460102
rect 277274 460046 277342 460102
rect 277398 460046 277494 460102
rect 276874 459978 277494 460046
rect 276874 459922 276970 459978
rect 277026 459922 277094 459978
rect 277150 459922 277218 459978
rect 277274 459922 277342 459978
rect 277398 459922 277494 459978
rect 276874 442350 277494 459922
rect 276874 442294 276970 442350
rect 277026 442294 277094 442350
rect 277150 442294 277218 442350
rect 277274 442294 277342 442350
rect 277398 442294 277494 442350
rect 276874 442226 277494 442294
rect 276874 442170 276970 442226
rect 277026 442170 277094 442226
rect 277150 442170 277218 442226
rect 277274 442170 277342 442226
rect 277398 442170 277494 442226
rect 276874 442102 277494 442170
rect 276874 442046 276970 442102
rect 277026 442046 277094 442102
rect 277150 442046 277218 442102
rect 277274 442046 277342 442102
rect 277398 442046 277494 442102
rect 276874 441978 277494 442046
rect 276874 441922 276970 441978
rect 277026 441922 277094 441978
rect 277150 441922 277218 441978
rect 277274 441922 277342 441978
rect 277398 441922 277494 441978
rect 276874 424350 277494 441922
rect 276874 424294 276970 424350
rect 277026 424294 277094 424350
rect 277150 424294 277218 424350
rect 277274 424294 277342 424350
rect 277398 424294 277494 424350
rect 276874 424226 277494 424294
rect 276874 424170 276970 424226
rect 277026 424170 277094 424226
rect 277150 424170 277218 424226
rect 277274 424170 277342 424226
rect 277398 424170 277494 424226
rect 276874 424102 277494 424170
rect 276874 424046 276970 424102
rect 277026 424046 277094 424102
rect 277150 424046 277218 424102
rect 277274 424046 277342 424102
rect 277398 424046 277494 424102
rect 276874 423978 277494 424046
rect 276874 423922 276970 423978
rect 277026 423922 277094 423978
rect 277150 423922 277218 423978
rect 277274 423922 277342 423978
rect 277398 423922 277494 423978
rect 276874 406350 277494 423922
rect 276874 406294 276970 406350
rect 277026 406294 277094 406350
rect 277150 406294 277218 406350
rect 277274 406294 277342 406350
rect 277398 406294 277494 406350
rect 276874 406226 277494 406294
rect 276874 406170 276970 406226
rect 277026 406170 277094 406226
rect 277150 406170 277218 406226
rect 277274 406170 277342 406226
rect 277398 406170 277494 406226
rect 276874 406102 277494 406170
rect 276874 406046 276970 406102
rect 277026 406046 277094 406102
rect 277150 406046 277218 406102
rect 277274 406046 277342 406102
rect 277398 406046 277494 406102
rect 276874 405978 277494 406046
rect 276874 405922 276970 405978
rect 277026 405922 277094 405978
rect 277150 405922 277218 405978
rect 277274 405922 277342 405978
rect 277398 405922 277494 405978
rect 276874 388350 277494 405922
rect 276874 388294 276970 388350
rect 277026 388294 277094 388350
rect 277150 388294 277218 388350
rect 277274 388294 277342 388350
rect 277398 388294 277494 388350
rect 276874 388226 277494 388294
rect 276874 388170 276970 388226
rect 277026 388170 277094 388226
rect 277150 388170 277218 388226
rect 277274 388170 277342 388226
rect 277398 388170 277494 388226
rect 276874 388102 277494 388170
rect 276874 388046 276970 388102
rect 277026 388046 277094 388102
rect 277150 388046 277218 388102
rect 277274 388046 277342 388102
rect 277398 388046 277494 388102
rect 276874 387978 277494 388046
rect 276874 387922 276970 387978
rect 277026 387922 277094 387978
rect 277150 387922 277218 387978
rect 277274 387922 277342 387978
rect 277398 387922 277494 387978
rect 276874 370350 277494 387922
rect 276874 370294 276970 370350
rect 277026 370294 277094 370350
rect 277150 370294 277218 370350
rect 277274 370294 277342 370350
rect 277398 370294 277494 370350
rect 276874 370226 277494 370294
rect 276874 370170 276970 370226
rect 277026 370170 277094 370226
rect 277150 370170 277218 370226
rect 277274 370170 277342 370226
rect 277398 370170 277494 370226
rect 276874 370102 277494 370170
rect 276874 370046 276970 370102
rect 277026 370046 277094 370102
rect 277150 370046 277218 370102
rect 277274 370046 277342 370102
rect 277398 370046 277494 370102
rect 276874 369978 277494 370046
rect 276874 369922 276970 369978
rect 277026 369922 277094 369978
rect 277150 369922 277218 369978
rect 277274 369922 277342 369978
rect 277398 369922 277494 369978
rect 276874 352350 277494 369922
rect 276874 352294 276970 352350
rect 277026 352294 277094 352350
rect 277150 352294 277218 352350
rect 277274 352294 277342 352350
rect 277398 352294 277494 352350
rect 276874 352226 277494 352294
rect 276874 352170 276970 352226
rect 277026 352170 277094 352226
rect 277150 352170 277218 352226
rect 277274 352170 277342 352226
rect 277398 352170 277494 352226
rect 276874 352102 277494 352170
rect 276874 352046 276970 352102
rect 277026 352046 277094 352102
rect 277150 352046 277218 352102
rect 277274 352046 277342 352102
rect 277398 352046 277494 352102
rect 276874 351978 277494 352046
rect 276874 351922 276970 351978
rect 277026 351922 277094 351978
rect 277150 351922 277218 351978
rect 277274 351922 277342 351978
rect 277398 351922 277494 351978
rect 276874 334350 277494 351922
rect 276874 334294 276970 334350
rect 277026 334294 277094 334350
rect 277150 334294 277218 334350
rect 277274 334294 277342 334350
rect 277398 334294 277494 334350
rect 276874 334226 277494 334294
rect 276874 334170 276970 334226
rect 277026 334170 277094 334226
rect 277150 334170 277218 334226
rect 277274 334170 277342 334226
rect 277398 334170 277494 334226
rect 276874 334102 277494 334170
rect 276874 334046 276970 334102
rect 277026 334046 277094 334102
rect 277150 334046 277218 334102
rect 277274 334046 277342 334102
rect 277398 334046 277494 334102
rect 276874 333978 277494 334046
rect 276874 333922 276970 333978
rect 277026 333922 277094 333978
rect 277150 333922 277218 333978
rect 277274 333922 277342 333978
rect 277398 333922 277494 333978
rect 276874 316350 277494 333922
rect 276874 316294 276970 316350
rect 277026 316294 277094 316350
rect 277150 316294 277218 316350
rect 277274 316294 277342 316350
rect 277398 316294 277494 316350
rect 276874 316226 277494 316294
rect 276874 316170 276970 316226
rect 277026 316170 277094 316226
rect 277150 316170 277218 316226
rect 277274 316170 277342 316226
rect 277398 316170 277494 316226
rect 276874 316102 277494 316170
rect 276874 316046 276970 316102
rect 277026 316046 277094 316102
rect 277150 316046 277218 316102
rect 277274 316046 277342 316102
rect 277398 316046 277494 316102
rect 276874 315978 277494 316046
rect 276874 315922 276970 315978
rect 277026 315922 277094 315978
rect 277150 315922 277218 315978
rect 277274 315922 277342 315978
rect 277398 315922 277494 315978
rect 276874 298350 277494 315922
rect 276874 298294 276970 298350
rect 277026 298294 277094 298350
rect 277150 298294 277218 298350
rect 277274 298294 277342 298350
rect 277398 298294 277494 298350
rect 276874 298226 277494 298294
rect 276874 298170 276970 298226
rect 277026 298170 277094 298226
rect 277150 298170 277218 298226
rect 277274 298170 277342 298226
rect 277398 298170 277494 298226
rect 276874 298102 277494 298170
rect 276874 298046 276970 298102
rect 277026 298046 277094 298102
rect 277150 298046 277218 298102
rect 277274 298046 277342 298102
rect 277398 298046 277494 298102
rect 276874 297978 277494 298046
rect 276874 297922 276970 297978
rect 277026 297922 277094 297978
rect 277150 297922 277218 297978
rect 277274 297922 277342 297978
rect 277398 297922 277494 297978
rect 276874 280350 277494 297922
rect 276874 280294 276970 280350
rect 277026 280294 277094 280350
rect 277150 280294 277218 280350
rect 277274 280294 277342 280350
rect 277398 280294 277494 280350
rect 276874 280226 277494 280294
rect 276874 280170 276970 280226
rect 277026 280170 277094 280226
rect 277150 280170 277218 280226
rect 277274 280170 277342 280226
rect 277398 280170 277494 280226
rect 276874 280102 277494 280170
rect 276874 280046 276970 280102
rect 277026 280046 277094 280102
rect 277150 280046 277218 280102
rect 277274 280046 277342 280102
rect 277398 280046 277494 280102
rect 276874 279978 277494 280046
rect 276874 279922 276970 279978
rect 277026 279922 277094 279978
rect 277150 279922 277218 279978
rect 277274 279922 277342 279978
rect 277398 279922 277494 279978
rect 276874 262350 277494 279922
rect 276874 262294 276970 262350
rect 277026 262294 277094 262350
rect 277150 262294 277218 262350
rect 277274 262294 277342 262350
rect 277398 262294 277494 262350
rect 276874 262226 277494 262294
rect 276874 262170 276970 262226
rect 277026 262170 277094 262226
rect 277150 262170 277218 262226
rect 277274 262170 277342 262226
rect 277398 262170 277494 262226
rect 276874 262102 277494 262170
rect 276874 262046 276970 262102
rect 277026 262046 277094 262102
rect 277150 262046 277218 262102
rect 277274 262046 277342 262102
rect 277398 262046 277494 262102
rect 276874 261978 277494 262046
rect 276874 261922 276970 261978
rect 277026 261922 277094 261978
rect 277150 261922 277218 261978
rect 277274 261922 277342 261978
rect 277398 261922 277494 261978
rect 276874 244350 277494 261922
rect 276874 244294 276970 244350
rect 277026 244294 277094 244350
rect 277150 244294 277218 244350
rect 277274 244294 277342 244350
rect 277398 244294 277494 244350
rect 276874 244226 277494 244294
rect 276874 244170 276970 244226
rect 277026 244170 277094 244226
rect 277150 244170 277218 244226
rect 277274 244170 277342 244226
rect 277398 244170 277494 244226
rect 276874 244102 277494 244170
rect 276874 244046 276970 244102
rect 277026 244046 277094 244102
rect 277150 244046 277218 244102
rect 277274 244046 277342 244102
rect 277398 244046 277494 244102
rect 276874 243978 277494 244046
rect 276874 243922 276970 243978
rect 277026 243922 277094 243978
rect 277150 243922 277218 243978
rect 277274 243922 277342 243978
rect 277398 243922 277494 243978
rect 276874 226350 277494 243922
rect 276874 226294 276970 226350
rect 277026 226294 277094 226350
rect 277150 226294 277218 226350
rect 277274 226294 277342 226350
rect 277398 226294 277494 226350
rect 276874 226226 277494 226294
rect 276874 226170 276970 226226
rect 277026 226170 277094 226226
rect 277150 226170 277218 226226
rect 277274 226170 277342 226226
rect 277398 226170 277494 226226
rect 276874 226102 277494 226170
rect 276874 226046 276970 226102
rect 277026 226046 277094 226102
rect 277150 226046 277218 226102
rect 277274 226046 277342 226102
rect 277398 226046 277494 226102
rect 276874 225978 277494 226046
rect 276874 225922 276970 225978
rect 277026 225922 277094 225978
rect 277150 225922 277218 225978
rect 277274 225922 277342 225978
rect 277398 225922 277494 225978
rect 273154 202294 273250 202350
rect 273306 202294 273374 202350
rect 273430 202294 273498 202350
rect 273554 202294 273622 202350
rect 273678 202294 273774 202350
rect 273154 202226 273774 202294
rect 273154 202170 273250 202226
rect 273306 202170 273374 202226
rect 273430 202170 273498 202226
rect 273554 202170 273622 202226
rect 273678 202170 273774 202226
rect 273154 202102 273774 202170
rect 273154 202046 273250 202102
rect 273306 202046 273374 202102
rect 273430 202046 273498 202102
rect 273554 202046 273622 202102
rect 273678 202046 273774 202102
rect 273154 201978 273774 202046
rect 273154 201922 273250 201978
rect 273306 201922 273374 201978
rect 273430 201922 273498 201978
rect 273554 201922 273622 201978
rect 273678 201922 273774 201978
rect 271292 198548 271348 198558
rect 269612 194516 269668 194526
rect 267932 186452 267988 186462
rect 266252 162978 266308 162988
rect 266364 170548 266420 170558
rect 264684 143938 264740 143948
rect 266364 138404 266420 170492
rect 267932 146244 267988 186396
rect 269612 150724 269668 194460
rect 269612 150658 269668 150668
rect 269724 160244 269780 160254
rect 267932 146178 267988 146188
rect 268044 150388 268100 150398
rect 266364 138338 266420 138348
rect 268044 128324 268100 150332
rect 269724 131684 269780 160188
rect 271292 152964 271348 198492
rect 273154 184350 273774 201922
rect 273154 184294 273250 184350
rect 273306 184294 273374 184350
rect 273430 184294 273498 184350
rect 273554 184294 273622 184350
rect 273678 184294 273774 184350
rect 273154 184226 273774 184294
rect 273154 184170 273250 184226
rect 273306 184170 273374 184226
rect 273430 184170 273498 184226
rect 273554 184170 273622 184226
rect 273678 184170 273774 184226
rect 273154 184102 273774 184170
rect 273154 184046 273250 184102
rect 273306 184046 273374 184102
rect 273430 184046 273498 184102
rect 273554 184046 273622 184102
rect 273678 184046 273774 184102
rect 273154 183978 273774 184046
rect 273154 183922 273250 183978
rect 273306 183922 273374 183978
rect 273430 183922 273498 183978
rect 273554 183922 273622 183978
rect 273678 183922 273774 183978
rect 271292 152898 271348 152908
rect 271404 170324 271460 170334
rect 271404 137284 271460 170268
rect 271404 137218 271460 137228
rect 273154 166350 273774 183922
rect 273154 166294 273250 166350
rect 273306 166294 273374 166350
rect 273430 166294 273498 166350
rect 273554 166294 273622 166350
rect 273678 166294 273774 166350
rect 273154 166226 273774 166294
rect 273154 166170 273250 166226
rect 273306 166170 273374 166226
rect 273430 166170 273498 166226
rect 273554 166170 273622 166226
rect 273678 166170 273774 166226
rect 273154 166102 273774 166170
rect 273154 166046 273250 166102
rect 273306 166046 273374 166102
rect 273430 166046 273498 166102
rect 273554 166046 273622 166102
rect 273678 166046 273774 166102
rect 273154 165978 273774 166046
rect 273154 165922 273250 165978
rect 273306 165922 273374 165978
rect 273430 165922 273498 165978
rect 273554 165922 273622 165978
rect 273678 165922 273774 165978
rect 273154 148350 273774 165922
rect 274652 217812 274708 217822
rect 274652 165284 274708 217756
rect 276874 208350 277494 225922
rect 276874 208294 276970 208350
rect 277026 208294 277094 208350
rect 277150 208294 277218 208350
rect 277274 208294 277342 208350
rect 277398 208294 277494 208350
rect 276874 208226 277494 208294
rect 276874 208170 276970 208226
rect 277026 208170 277094 208226
rect 277150 208170 277218 208226
rect 277274 208170 277342 208226
rect 277398 208170 277494 208226
rect 276874 208102 277494 208170
rect 276874 208046 276970 208102
rect 277026 208046 277094 208102
rect 277150 208046 277218 208102
rect 277274 208046 277342 208102
rect 277398 208046 277494 208102
rect 276874 207978 277494 208046
rect 276874 207922 276970 207978
rect 277026 207922 277094 207978
rect 277150 207922 277218 207978
rect 277274 207922 277342 207978
rect 277398 207922 277494 207978
rect 276874 190350 277494 207922
rect 276874 190294 276970 190350
rect 277026 190294 277094 190350
rect 277150 190294 277218 190350
rect 277274 190294 277342 190350
rect 277398 190294 277494 190350
rect 276874 190226 277494 190294
rect 276874 190170 276970 190226
rect 277026 190170 277094 190226
rect 277150 190170 277218 190226
rect 277274 190170 277342 190226
rect 277398 190170 277494 190226
rect 276874 190102 277494 190170
rect 276874 190046 276970 190102
rect 277026 190046 277094 190102
rect 277150 190046 277218 190102
rect 277274 190046 277342 190102
rect 277398 190046 277494 190102
rect 276874 189978 277494 190046
rect 276874 189922 276970 189978
rect 277026 189922 277094 189978
rect 277150 189922 277218 189978
rect 277274 189922 277342 189978
rect 277398 189922 277494 189978
rect 276332 189028 276388 189038
rect 274652 165218 274708 165228
rect 274764 176372 274820 176382
rect 273154 148294 273250 148350
rect 273306 148294 273374 148350
rect 273430 148294 273498 148350
rect 273554 148294 273622 148350
rect 273678 148294 273774 148350
rect 273154 148226 273774 148294
rect 273154 148170 273250 148226
rect 273306 148170 273374 148226
rect 273430 148170 273498 148226
rect 273554 148170 273622 148226
rect 273678 148170 273774 148226
rect 273154 148102 273774 148170
rect 273154 148046 273250 148102
rect 273306 148046 273374 148102
rect 273430 148046 273498 148102
rect 273554 148046 273622 148102
rect 273678 148046 273774 148102
rect 273154 147978 273774 148046
rect 273154 147922 273250 147978
rect 273306 147922 273374 147978
rect 273430 147922 273498 147978
rect 273554 147922 273622 147978
rect 273678 147922 273774 147978
rect 269724 131618 269780 131628
rect 268044 128258 268100 128268
rect 273154 130350 273774 147922
rect 273154 130294 273250 130350
rect 273306 130294 273374 130350
rect 273430 130294 273498 130350
rect 273554 130294 273622 130350
rect 273678 130294 273774 130350
rect 273154 130226 273774 130294
rect 273154 130170 273250 130226
rect 273306 130170 273374 130226
rect 273430 130170 273498 130226
rect 273554 130170 273622 130226
rect 273678 130170 273774 130226
rect 273154 130102 273774 130170
rect 273154 130046 273250 130102
rect 273306 130046 273374 130102
rect 273430 130046 273498 130102
rect 273554 130046 273622 130102
rect 273678 130046 273774 130102
rect 273154 129978 273774 130046
rect 273154 129922 273250 129978
rect 273306 129922 273374 129978
rect 273430 129922 273498 129978
rect 273554 129922 273622 129978
rect 273678 129922 273774 129978
rect 264572 127138 264628 127148
rect 268268 127988 268324 127998
rect 258874 118294 258970 118350
rect 259026 118294 259094 118350
rect 259150 118294 259218 118350
rect 259274 118294 259342 118350
rect 259398 118294 259494 118350
rect 258874 118226 259494 118294
rect 258874 118170 258970 118226
rect 259026 118170 259094 118226
rect 259150 118170 259218 118226
rect 259274 118170 259342 118226
rect 259398 118170 259494 118226
rect 258874 118102 259494 118170
rect 258874 118046 258970 118102
rect 259026 118046 259094 118102
rect 259150 118046 259218 118102
rect 259274 118046 259342 118102
rect 259398 118046 259494 118102
rect 258874 117978 259494 118046
rect 258874 117922 258970 117978
rect 259026 117922 259094 117978
rect 259150 117922 259218 117978
rect 259274 117922 259342 117978
rect 259398 117922 259494 117978
rect 255154 112294 255250 112350
rect 255306 112294 255374 112350
rect 255430 112294 255498 112350
rect 255554 112294 255622 112350
rect 255678 112294 255774 112350
rect 255154 112226 255774 112294
rect 255154 112170 255250 112226
rect 255306 112170 255374 112226
rect 255430 112170 255498 112226
rect 255554 112170 255622 112226
rect 255678 112170 255774 112226
rect 255154 112102 255774 112170
rect 255154 112046 255250 112102
rect 255306 112046 255374 112102
rect 255430 112046 255498 112102
rect 255554 112046 255622 112102
rect 255678 112046 255774 112102
rect 255154 111978 255774 112046
rect 255154 111922 255250 111978
rect 255306 111922 255374 111978
rect 255430 111922 255498 111978
rect 255554 111922 255622 111978
rect 255678 111922 255774 111978
rect 255154 94350 255774 111922
rect 255154 94294 255250 94350
rect 255306 94294 255374 94350
rect 255430 94294 255498 94350
rect 255554 94294 255622 94350
rect 255678 94294 255774 94350
rect 255154 94226 255774 94294
rect 255154 94170 255250 94226
rect 255306 94170 255374 94226
rect 255430 94170 255498 94226
rect 255554 94170 255622 94226
rect 255678 94170 255774 94226
rect 255154 94102 255774 94170
rect 255154 94046 255250 94102
rect 255306 94046 255374 94102
rect 255430 94046 255498 94102
rect 255554 94046 255622 94102
rect 255678 94046 255774 94102
rect 255154 93978 255774 94046
rect 255154 93922 255250 93978
rect 255306 93922 255374 93978
rect 255430 93922 255498 93978
rect 255554 93922 255622 93978
rect 255678 93922 255774 93978
rect 244524 84644 244580 84654
rect 244524 75572 244580 84588
rect 244524 75506 244580 75516
rect 255154 76350 255774 93922
rect 255154 76294 255250 76350
rect 255306 76294 255374 76350
rect 255430 76294 255498 76350
rect 255554 76294 255622 76350
rect 255678 76294 255774 76350
rect 255154 76226 255774 76294
rect 255154 76170 255250 76226
rect 255306 76170 255374 76226
rect 255430 76170 255498 76226
rect 255554 76170 255622 76226
rect 255678 76170 255774 76226
rect 255154 76102 255774 76170
rect 255154 76046 255250 76102
rect 255306 76046 255374 76102
rect 255430 76046 255498 76102
rect 255554 76046 255622 76102
rect 255678 76046 255774 76102
rect 255154 75978 255774 76046
rect 255154 75922 255250 75978
rect 255306 75922 255374 75978
rect 255430 75922 255498 75978
rect 255554 75922 255622 75978
rect 255678 75922 255774 75978
rect 244524 73108 244580 73118
rect 244524 61460 244580 73052
rect 244524 61394 244580 61404
rect 244412 29572 244468 29582
rect 255154 58350 255774 75922
rect 255154 58294 255250 58350
rect 255306 58294 255374 58350
rect 255430 58294 255498 58350
rect 255554 58294 255622 58350
rect 255678 58294 255774 58350
rect 255154 58226 255774 58294
rect 255154 58170 255250 58226
rect 255306 58170 255374 58226
rect 255430 58170 255498 58226
rect 255554 58170 255622 58226
rect 255678 58170 255774 58226
rect 255154 58102 255774 58170
rect 255154 58046 255250 58102
rect 255306 58046 255374 58102
rect 255430 58046 255498 58102
rect 255554 58046 255622 58102
rect 255678 58046 255774 58102
rect 255154 57978 255774 58046
rect 255154 57922 255250 57978
rect 255306 57922 255374 57978
rect 255430 57922 255498 57978
rect 255554 57922 255622 57978
rect 255678 57922 255774 57978
rect 255154 40350 255774 57922
rect 255154 40294 255250 40350
rect 255306 40294 255374 40350
rect 255430 40294 255498 40350
rect 255554 40294 255622 40350
rect 255678 40294 255774 40350
rect 255154 40226 255774 40294
rect 255154 40170 255250 40226
rect 255306 40170 255374 40226
rect 255430 40170 255498 40226
rect 255554 40170 255622 40226
rect 255678 40170 255774 40226
rect 255154 40102 255774 40170
rect 255154 40046 255250 40102
rect 255306 40046 255374 40102
rect 255430 40046 255498 40102
rect 255554 40046 255622 40102
rect 255678 40046 255774 40102
rect 255154 39978 255774 40046
rect 255154 39922 255250 39978
rect 255306 39922 255374 39978
rect 255430 39922 255498 39978
rect 255554 39922 255622 39978
rect 255678 39922 255774 39978
rect 240874 28294 240970 28350
rect 241026 28294 241094 28350
rect 241150 28294 241218 28350
rect 241274 28294 241342 28350
rect 241398 28294 241494 28350
rect 240874 28226 241494 28294
rect 240874 28170 240970 28226
rect 241026 28170 241094 28226
rect 241150 28170 241218 28226
rect 241274 28170 241342 28226
rect 241398 28170 241494 28226
rect 240874 28102 241494 28170
rect 240874 28046 240970 28102
rect 241026 28046 241094 28102
rect 241150 28046 241218 28102
rect 241274 28046 241342 28102
rect 241398 28046 241494 28102
rect 240874 27978 241494 28046
rect 240874 27922 240970 27978
rect 241026 27922 241094 27978
rect 241150 27922 241218 27978
rect 241274 27922 241342 27978
rect 241398 27922 241494 27978
rect 237154 22294 237250 22350
rect 237306 22294 237374 22350
rect 237430 22294 237498 22350
rect 237554 22294 237622 22350
rect 237678 22294 237774 22350
rect 237154 22226 237774 22294
rect 237154 22170 237250 22226
rect 237306 22170 237374 22226
rect 237430 22170 237498 22226
rect 237554 22170 237622 22226
rect 237678 22170 237774 22226
rect 237154 22102 237774 22170
rect 237154 22046 237250 22102
rect 237306 22046 237374 22102
rect 237430 22046 237498 22102
rect 237554 22046 237622 22102
rect 237678 22046 237774 22102
rect 237154 21978 237774 22046
rect 237154 21922 237250 21978
rect 237306 21922 237374 21978
rect 237430 21922 237498 21978
rect 237554 21922 237622 21978
rect 237678 21922 237774 21978
rect 237154 4350 237774 21922
rect 237154 4294 237250 4350
rect 237306 4294 237374 4350
rect 237430 4294 237498 4350
rect 237554 4294 237622 4350
rect 237678 4294 237774 4350
rect 237154 4226 237774 4294
rect 237154 4170 237250 4226
rect 237306 4170 237374 4226
rect 237430 4170 237498 4226
rect 237554 4170 237622 4226
rect 237678 4170 237774 4226
rect 237154 4102 237774 4170
rect 237154 4046 237250 4102
rect 237306 4046 237374 4102
rect 237430 4046 237498 4102
rect 237554 4046 237622 4102
rect 237678 4046 237774 4102
rect 237154 3978 237774 4046
rect 237154 3922 237250 3978
rect 237306 3922 237374 3978
rect 237430 3922 237498 3978
rect 237554 3922 237622 3978
rect 237678 3922 237774 3978
rect 237154 -160 237774 3922
rect 237154 -216 237250 -160
rect 237306 -216 237374 -160
rect 237430 -216 237498 -160
rect 237554 -216 237622 -160
rect 237678 -216 237774 -160
rect 237154 -284 237774 -216
rect 237154 -340 237250 -284
rect 237306 -340 237374 -284
rect 237430 -340 237498 -284
rect 237554 -340 237622 -284
rect 237678 -340 237774 -284
rect 237154 -408 237774 -340
rect 237154 -464 237250 -408
rect 237306 -464 237374 -408
rect 237430 -464 237498 -408
rect 237554 -464 237622 -408
rect 237678 -464 237774 -408
rect 237154 -532 237774 -464
rect 237154 -588 237250 -532
rect 237306 -588 237374 -532
rect 237430 -588 237498 -532
rect 237554 -588 237622 -532
rect 237678 -588 237774 -532
rect 237154 -1644 237774 -588
rect 240874 10350 241494 27922
rect 240874 10294 240970 10350
rect 241026 10294 241094 10350
rect 241150 10294 241218 10350
rect 241274 10294 241342 10350
rect 241398 10294 241494 10350
rect 240874 10226 241494 10294
rect 240874 10170 240970 10226
rect 241026 10170 241094 10226
rect 241150 10170 241218 10226
rect 241274 10170 241342 10226
rect 241398 10170 241494 10226
rect 240874 10102 241494 10170
rect 240874 10046 240970 10102
rect 241026 10046 241094 10102
rect 241150 10046 241218 10102
rect 241274 10046 241342 10102
rect 241398 10046 241494 10102
rect 240874 9978 241494 10046
rect 240874 9922 240970 9978
rect 241026 9922 241094 9978
rect 241150 9922 241218 9978
rect 241274 9922 241342 9978
rect 241398 9922 241494 9978
rect 240874 -1120 241494 9922
rect 240874 -1176 240970 -1120
rect 241026 -1176 241094 -1120
rect 241150 -1176 241218 -1120
rect 241274 -1176 241342 -1120
rect 241398 -1176 241494 -1120
rect 240874 -1244 241494 -1176
rect 240874 -1300 240970 -1244
rect 241026 -1300 241094 -1244
rect 241150 -1300 241218 -1244
rect 241274 -1300 241342 -1244
rect 241398 -1300 241494 -1244
rect 240874 -1368 241494 -1300
rect 240874 -1424 240970 -1368
rect 241026 -1424 241094 -1368
rect 241150 -1424 241218 -1368
rect 241274 -1424 241342 -1368
rect 241398 -1424 241494 -1368
rect 240874 -1492 241494 -1424
rect 240874 -1548 240970 -1492
rect 241026 -1548 241094 -1492
rect 241150 -1548 241218 -1492
rect 241274 -1548 241342 -1492
rect 241398 -1548 241494 -1492
rect 240874 -1644 241494 -1548
rect 255154 22350 255774 39922
rect 255154 22294 255250 22350
rect 255306 22294 255374 22350
rect 255430 22294 255498 22350
rect 255554 22294 255622 22350
rect 255678 22294 255774 22350
rect 255154 22226 255774 22294
rect 255154 22170 255250 22226
rect 255306 22170 255374 22226
rect 255430 22170 255498 22226
rect 255554 22170 255622 22226
rect 255678 22170 255774 22226
rect 255154 22102 255774 22170
rect 255154 22046 255250 22102
rect 255306 22046 255374 22102
rect 255430 22046 255498 22102
rect 255554 22046 255622 22102
rect 255678 22046 255774 22102
rect 255154 21978 255774 22046
rect 255154 21922 255250 21978
rect 255306 21922 255374 21978
rect 255430 21922 255498 21978
rect 255554 21922 255622 21978
rect 255678 21922 255774 21978
rect 255154 4350 255774 21922
rect 255154 4294 255250 4350
rect 255306 4294 255374 4350
rect 255430 4294 255498 4350
rect 255554 4294 255622 4350
rect 255678 4294 255774 4350
rect 255154 4226 255774 4294
rect 255154 4170 255250 4226
rect 255306 4170 255374 4226
rect 255430 4170 255498 4226
rect 255554 4170 255622 4226
rect 255678 4170 255774 4226
rect 255154 4102 255774 4170
rect 255154 4046 255250 4102
rect 255306 4046 255374 4102
rect 255430 4046 255498 4102
rect 255554 4046 255622 4102
rect 255678 4046 255774 4102
rect 255154 3978 255774 4046
rect 255154 3922 255250 3978
rect 255306 3922 255374 3978
rect 255430 3922 255498 3978
rect 255554 3922 255622 3978
rect 255678 3922 255774 3978
rect 255154 -160 255774 3922
rect 255154 -216 255250 -160
rect 255306 -216 255374 -160
rect 255430 -216 255498 -160
rect 255554 -216 255622 -160
rect 255678 -216 255774 -160
rect 255154 -284 255774 -216
rect 255154 -340 255250 -284
rect 255306 -340 255374 -284
rect 255430 -340 255498 -284
rect 255554 -340 255622 -284
rect 255678 -340 255774 -284
rect 255154 -408 255774 -340
rect 255154 -464 255250 -408
rect 255306 -464 255374 -408
rect 255430 -464 255498 -408
rect 255554 -464 255622 -408
rect 255678 -464 255774 -408
rect 255154 -532 255774 -464
rect 255154 -588 255250 -532
rect 255306 -588 255374 -532
rect 255430 -588 255498 -532
rect 255554 -588 255622 -532
rect 255678 -588 255774 -532
rect 255154 -1644 255774 -588
rect 258874 100350 259494 117922
rect 268268 113764 268324 127932
rect 268268 113698 268324 113708
rect 258874 100294 258970 100350
rect 259026 100294 259094 100350
rect 259150 100294 259218 100350
rect 259274 100294 259342 100350
rect 259398 100294 259494 100350
rect 258874 100226 259494 100294
rect 258874 100170 258970 100226
rect 259026 100170 259094 100226
rect 259150 100170 259218 100226
rect 259274 100170 259342 100226
rect 259398 100170 259494 100226
rect 258874 100102 259494 100170
rect 258874 100046 258970 100102
rect 259026 100046 259094 100102
rect 259150 100046 259218 100102
rect 259274 100046 259342 100102
rect 259398 100046 259494 100102
rect 258874 99978 259494 100046
rect 258874 99922 258970 99978
rect 259026 99922 259094 99978
rect 259150 99922 259218 99978
rect 259274 99922 259342 99978
rect 259398 99922 259494 99978
rect 258874 82350 259494 99922
rect 258874 82294 258970 82350
rect 259026 82294 259094 82350
rect 259150 82294 259218 82350
rect 259274 82294 259342 82350
rect 259398 82294 259494 82350
rect 258874 82226 259494 82294
rect 258874 82170 258970 82226
rect 259026 82170 259094 82226
rect 259150 82170 259218 82226
rect 259274 82170 259342 82226
rect 259398 82170 259494 82226
rect 258874 82102 259494 82170
rect 258874 82046 258970 82102
rect 259026 82046 259094 82102
rect 259150 82046 259218 82102
rect 259274 82046 259342 82102
rect 259398 82046 259494 82102
rect 258874 81978 259494 82046
rect 258874 81922 258970 81978
rect 259026 81922 259094 81978
rect 259150 81922 259218 81978
rect 259274 81922 259342 81978
rect 259398 81922 259494 81978
rect 258874 64350 259494 81922
rect 258874 64294 258970 64350
rect 259026 64294 259094 64350
rect 259150 64294 259218 64350
rect 259274 64294 259342 64350
rect 259398 64294 259494 64350
rect 258874 64226 259494 64294
rect 258874 64170 258970 64226
rect 259026 64170 259094 64226
rect 259150 64170 259218 64226
rect 259274 64170 259342 64226
rect 259398 64170 259494 64226
rect 258874 64102 259494 64170
rect 258874 64046 258970 64102
rect 259026 64046 259094 64102
rect 259150 64046 259218 64102
rect 259274 64046 259342 64102
rect 259398 64046 259494 64102
rect 258874 63978 259494 64046
rect 258874 63922 258970 63978
rect 259026 63922 259094 63978
rect 259150 63922 259218 63978
rect 259274 63922 259342 63978
rect 259398 63922 259494 63978
rect 258874 46350 259494 63922
rect 258874 46294 258970 46350
rect 259026 46294 259094 46350
rect 259150 46294 259218 46350
rect 259274 46294 259342 46350
rect 259398 46294 259494 46350
rect 258874 46226 259494 46294
rect 258874 46170 258970 46226
rect 259026 46170 259094 46226
rect 259150 46170 259218 46226
rect 259274 46170 259342 46226
rect 259398 46170 259494 46226
rect 258874 46102 259494 46170
rect 258874 46046 258970 46102
rect 259026 46046 259094 46102
rect 259150 46046 259218 46102
rect 259274 46046 259342 46102
rect 259398 46046 259494 46102
rect 258874 45978 259494 46046
rect 258874 45922 258970 45978
rect 259026 45922 259094 45978
rect 259150 45922 259218 45978
rect 259274 45922 259342 45978
rect 259398 45922 259494 45978
rect 258874 28350 259494 45922
rect 258874 28294 258970 28350
rect 259026 28294 259094 28350
rect 259150 28294 259218 28350
rect 259274 28294 259342 28350
rect 259398 28294 259494 28350
rect 258874 28226 259494 28294
rect 258874 28170 258970 28226
rect 259026 28170 259094 28226
rect 259150 28170 259218 28226
rect 259274 28170 259342 28226
rect 259398 28170 259494 28226
rect 258874 28102 259494 28170
rect 258874 28046 258970 28102
rect 259026 28046 259094 28102
rect 259150 28046 259218 28102
rect 259274 28046 259342 28102
rect 259398 28046 259494 28102
rect 258874 27978 259494 28046
rect 258874 27922 258970 27978
rect 259026 27922 259094 27978
rect 259150 27922 259218 27978
rect 259274 27922 259342 27978
rect 259398 27922 259494 27978
rect 258874 10350 259494 27922
rect 258874 10294 258970 10350
rect 259026 10294 259094 10350
rect 259150 10294 259218 10350
rect 259274 10294 259342 10350
rect 259398 10294 259494 10350
rect 258874 10226 259494 10294
rect 258874 10170 258970 10226
rect 259026 10170 259094 10226
rect 259150 10170 259218 10226
rect 259274 10170 259342 10226
rect 259398 10170 259494 10226
rect 258874 10102 259494 10170
rect 258874 10046 258970 10102
rect 259026 10046 259094 10102
rect 259150 10046 259218 10102
rect 259274 10046 259342 10102
rect 259398 10046 259494 10102
rect 258874 9978 259494 10046
rect 258874 9922 258970 9978
rect 259026 9922 259094 9978
rect 259150 9922 259218 9978
rect 259274 9922 259342 9978
rect 259398 9922 259494 9978
rect 258874 -1120 259494 9922
rect 258874 -1176 258970 -1120
rect 259026 -1176 259094 -1120
rect 259150 -1176 259218 -1120
rect 259274 -1176 259342 -1120
rect 259398 -1176 259494 -1120
rect 258874 -1244 259494 -1176
rect 258874 -1300 258970 -1244
rect 259026 -1300 259094 -1244
rect 259150 -1300 259218 -1244
rect 259274 -1300 259342 -1244
rect 259398 -1300 259494 -1244
rect 258874 -1368 259494 -1300
rect 258874 -1424 258970 -1368
rect 259026 -1424 259094 -1368
rect 259150 -1424 259218 -1368
rect 259274 -1424 259342 -1368
rect 259398 -1424 259494 -1368
rect 258874 -1492 259494 -1424
rect 258874 -1548 258970 -1492
rect 259026 -1548 259094 -1492
rect 259150 -1548 259218 -1492
rect 259274 -1548 259342 -1492
rect 259398 -1548 259494 -1492
rect 258874 -1644 259494 -1548
rect 273154 112350 273774 129922
rect 274652 156212 274708 156222
rect 274652 129444 274708 156156
rect 274764 140644 274820 176316
rect 275548 155428 275604 155438
rect 275548 154084 275604 155372
rect 276332 155204 276388 188972
rect 276444 185668 276500 185678
rect 276444 157444 276500 185612
rect 276556 175588 276612 175598
rect 276556 160804 276612 175532
rect 276556 160738 276612 160748
rect 276874 172350 277494 189922
rect 276874 172294 276970 172350
rect 277026 172294 277094 172350
rect 277150 172294 277218 172350
rect 277274 172294 277342 172350
rect 277398 172294 277494 172350
rect 276874 172226 277494 172294
rect 276874 172170 276970 172226
rect 277026 172170 277094 172226
rect 277150 172170 277218 172226
rect 277274 172170 277342 172226
rect 277398 172170 277494 172226
rect 276874 172102 277494 172170
rect 276874 172046 276970 172102
rect 277026 172046 277094 172102
rect 277150 172046 277218 172102
rect 277274 172046 277342 172102
rect 277398 172046 277494 172102
rect 276874 171978 277494 172046
rect 276874 171922 276970 171978
rect 277026 171922 277094 171978
rect 277150 171922 277218 171978
rect 277274 171922 277342 171978
rect 277398 171922 277494 171978
rect 276444 157378 276500 157388
rect 276332 155138 276388 155148
rect 275548 154018 275604 154028
rect 276874 154350 277494 171922
rect 291154 597212 291774 598268
rect 291154 597156 291250 597212
rect 291306 597156 291374 597212
rect 291430 597156 291498 597212
rect 291554 597156 291622 597212
rect 291678 597156 291774 597212
rect 291154 597088 291774 597156
rect 291154 597032 291250 597088
rect 291306 597032 291374 597088
rect 291430 597032 291498 597088
rect 291554 597032 291622 597088
rect 291678 597032 291774 597088
rect 291154 596964 291774 597032
rect 291154 596908 291250 596964
rect 291306 596908 291374 596964
rect 291430 596908 291498 596964
rect 291554 596908 291622 596964
rect 291678 596908 291774 596964
rect 291154 596840 291774 596908
rect 291154 596784 291250 596840
rect 291306 596784 291374 596840
rect 291430 596784 291498 596840
rect 291554 596784 291622 596840
rect 291678 596784 291774 596840
rect 291154 580350 291774 596784
rect 291154 580294 291250 580350
rect 291306 580294 291374 580350
rect 291430 580294 291498 580350
rect 291554 580294 291622 580350
rect 291678 580294 291774 580350
rect 291154 580226 291774 580294
rect 291154 580170 291250 580226
rect 291306 580170 291374 580226
rect 291430 580170 291498 580226
rect 291554 580170 291622 580226
rect 291678 580170 291774 580226
rect 291154 580102 291774 580170
rect 291154 580046 291250 580102
rect 291306 580046 291374 580102
rect 291430 580046 291498 580102
rect 291554 580046 291622 580102
rect 291678 580046 291774 580102
rect 291154 579978 291774 580046
rect 291154 579922 291250 579978
rect 291306 579922 291374 579978
rect 291430 579922 291498 579978
rect 291554 579922 291622 579978
rect 291678 579922 291774 579978
rect 291154 562350 291774 579922
rect 291154 562294 291250 562350
rect 291306 562294 291374 562350
rect 291430 562294 291498 562350
rect 291554 562294 291622 562350
rect 291678 562294 291774 562350
rect 291154 562226 291774 562294
rect 291154 562170 291250 562226
rect 291306 562170 291374 562226
rect 291430 562170 291498 562226
rect 291554 562170 291622 562226
rect 291678 562170 291774 562226
rect 291154 562102 291774 562170
rect 291154 562046 291250 562102
rect 291306 562046 291374 562102
rect 291430 562046 291498 562102
rect 291554 562046 291622 562102
rect 291678 562046 291774 562102
rect 291154 561978 291774 562046
rect 291154 561922 291250 561978
rect 291306 561922 291374 561978
rect 291430 561922 291498 561978
rect 291554 561922 291622 561978
rect 291678 561922 291774 561978
rect 291154 544350 291774 561922
rect 291154 544294 291250 544350
rect 291306 544294 291374 544350
rect 291430 544294 291498 544350
rect 291554 544294 291622 544350
rect 291678 544294 291774 544350
rect 291154 544226 291774 544294
rect 291154 544170 291250 544226
rect 291306 544170 291374 544226
rect 291430 544170 291498 544226
rect 291554 544170 291622 544226
rect 291678 544170 291774 544226
rect 291154 544102 291774 544170
rect 291154 544046 291250 544102
rect 291306 544046 291374 544102
rect 291430 544046 291498 544102
rect 291554 544046 291622 544102
rect 291678 544046 291774 544102
rect 291154 543978 291774 544046
rect 291154 543922 291250 543978
rect 291306 543922 291374 543978
rect 291430 543922 291498 543978
rect 291554 543922 291622 543978
rect 291678 543922 291774 543978
rect 291154 526350 291774 543922
rect 291154 526294 291250 526350
rect 291306 526294 291374 526350
rect 291430 526294 291498 526350
rect 291554 526294 291622 526350
rect 291678 526294 291774 526350
rect 291154 526226 291774 526294
rect 291154 526170 291250 526226
rect 291306 526170 291374 526226
rect 291430 526170 291498 526226
rect 291554 526170 291622 526226
rect 291678 526170 291774 526226
rect 291154 526102 291774 526170
rect 291154 526046 291250 526102
rect 291306 526046 291374 526102
rect 291430 526046 291498 526102
rect 291554 526046 291622 526102
rect 291678 526046 291774 526102
rect 291154 525978 291774 526046
rect 291154 525922 291250 525978
rect 291306 525922 291374 525978
rect 291430 525922 291498 525978
rect 291554 525922 291622 525978
rect 291678 525922 291774 525978
rect 291154 508350 291774 525922
rect 291154 508294 291250 508350
rect 291306 508294 291374 508350
rect 291430 508294 291498 508350
rect 291554 508294 291622 508350
rect 291678 508294 291774 508350
rect 291154 508226 291774 508294
rect 291154 508170 291250 508226
rect 291306 508170 291374 508226
rect 291430 508170 291498 508226
rect 291554 508170 291622 508226
rect 291678 508170 291774 508226
rect 291154 508102 291774 508170
rect 291154 508046 291250 508102
rect 291306 508046 291374 508102
rect 291430 508046 291498 508102
rect 291554 508046 291622 508102
rect 291678 508046 291774 508102
rect 291154 507978 291774 508046
rect 291154 507922 291250 507978
rect 291306 507922 291374 507978
rect 291430 507922 291498 507978
rect 291554 507922 291622 507978
rect 291678 507922 291774 507978
rect 291154 490350 291774 507922
rect 291154 490294 291250 490350
rect 291306 490294 291374 490350
rect 291430 490294 291498 490350
rect 291554 490294 291622 490350
rect 291678 490294 291774 490350
rect 291154 490226 291774 490294
rect 291154 490170 291250 490226
rect 291306 490170 291374 490226
rect 291430 490170 291498 490226
rect 291554 490170 291622 490226
rect 291678 490170 291774 490226
rect 291154 490102 291774 490170
rect 291154 490046 291250 490102
rect 291306 490046 291374 490102
rect 291430 490046 291498 490102
rect 291554 490046 291622 490102
rect 291678 490046 291774 490102
rect 291154 489978 291774 490046
rect 291154 489922 291250 489978
rect 291306 489922 291374 489978
rect 291430 489922 291498 489978
rect 291554 489922 291622 489978
rect 291678 489922 291774 489978
rect 291154 472350 291774 489922
rect 291154 472294 291250 472350
rect 291306 472294 291374 472350
rect 291430 472294 291498 472350
rect 291554 472294 291622 472350
rect 291678 472294 291774 472350
rect 291154 472226 291774 472294
rect 291154 472170 291250 472226
rect 291306 472170 291374 472226
rect 291430 472170 291498 472226
rect 291554 472170 291622 472226
rect 291678 472170 291774 472226
rect 291154 472102 291774 472170
rect 291154 472046 291250 472102
rect 291306 472046 291374 472102
rect 291430 472046 291498 472102
rect 291554 472046 291622 472102
rect 291678 472046 291774 472102
rect 291154 471978 291774 472046
rect 291154 471922 291250 471978
rect 291306 471922 291374 471978
rect 291430 471922 291498 471978
rect 291554 471922 291622 471978
rect 291678 471922 291774 471978
rect 291154 454350 291774 471922
rect 291154 454294 291250 454350
rect 291306 454294 291374 454350
rect 291430 454294 291498 454350
rect 291554 454294 291622 454350
rect 291678 454294 291774 454350
rect 291154 454226 291774 454294
rect 291154 454170 291250 454226
rect 291306 454170 291374 454226
rect 291430 454170 291498 454226
rect 291554 454170 291622 454226
rect 291678 454170 291774 454226
rect 291154 454102 291774 454170
rect 291154 454046 291250 454102
rect 291306 454046 291374 454102
rect 291430 454046 291498 454102
rect 291554 454046 291622 454102
rect 291678 454046 291774 454102
rect 291154 453978 291774 454046
rect 291154 453922 291250 453978
rect 291306 453922 291374 453978
rect 291430 453922 291498 453978
rect 291554 453922 291622 453978
rect 291678 453922 291774 453978
rect 291154 436350 291774 453922
rect 291154 436294 291250 436350
rect 291306 436294 291374 436350
rect 291430 436294 291498 436350
rect 291554 436294 291622 436350
rect 291678 436294 291774 436350
rect 291154 436226 291774 436294
rect 291154 436170 291250 436226
rect 291306 436170 291374 436226
rect 291430 436170 291498 436226
rect 291554 436170 291622 436226
rect 291678 436170 291774 436226
rect 291154 436102 291774 436170
rect 291154 436046 291250 436102
rect 291306 436046 291374 436102
rect 291430 436046 291498 436102
rect 291554 436046 291622 436102
rect 291678 436046 291774 436102
rect 291154 435978 291774 436046
rect 291154 435922 291250 435978
rect 291306 435922 291374 435978
rect 291430 435922 291498 435978
rect 291554 435922 291622 435978
rect 291678 435922 291774 435978
rect 291154 418350 291774 435922
rect 291154 418294 291250 418350
rect 291306 418294 291374 418350
rect 291430 418294 291498 418350
rect 291554 418294 291622 418350
rect 291678 418294 291774 418350
rect 291154 418226 291774 418294
rect 291154 418170 291250 418226
rect 291306 418170 291374 418226
rect 291430 418170 291498 418226
rect 291554 418170 291622 418226
rect 291678 418170 291774 418226
rect 291154 418102 291774 418170
rect 291154 418046 291250 418102
rect 291306 418046 291374 418102
rect 291430 418046 291498 418102
rect 291554 418046 291622 418102
rect 291678 418046 291774 418102
rect 291154 417978 291774 418046
rect 291154 417922 291250 417978
rect 291306 417922 291374 417978
rect 291430 417922 291498 417978
rect 291554 417922 291622 417978
rect 291678 417922 291774 417978
rect 291154 400350 291774 417922
rect 291154 400294 291250 400350
rect 291306 400294 291374 400350
rect 291430 400294 291498 400350
rect 291554 400294 291622 400350
rect 291678 400294 291774 400350
rect 291154 400226 291774 400294
rect 291154 400170 291250 400226
rect 291306 400170 291374 400226
rect 291430 400170 291498 400226
rect 291554 400170 291622 400226
rect 291678 400170 291774 400226
rect 291154 400102 291774 400170
rect 291154 400046 291250 400102
rect 291306 400046 291374 400102
rect 291430 400046 291498 400102
rect 291554 400046 291622 400102
rect 291678 400046 291774 400102
rect 291154 399978 291774 400046
rect 291154 399922 291250 399978
rect 291306 399922 291374 399978
rect 291430 399922 291498 399978
rect 291554 399922 291622 399978
rect 291678 399922 291774 399978
rect 291154 382350 291774 399922
rect 291154 382294 291250 382350
rect 291306 382294 291374 382350
rect 291430 382294 291498 382350
rect 291554 382294 291622 382350
rect 291678 382294 291774 382350
rect 291154 382226 291774 382294
rect 291154 382170 291250 382226
rect 291306 382170 291374 382226
rect 291430 382170 291498 382226
rect 291554 382170 291622 382226
rect 291678 382170 291774 382226
rect 291154 382102 291774 382170
rect 291154 382046 291250 382102
rect 291306 382046 291374 382102
rect 291430 382046 291498 382102
rect 291554 382046 291622 382102
rect 291678 382046 291774 382102
rect 291154 381978 291774 382046
rect 291154 381922 291250 381978
rect 291306 381922 291374 381978
rect 291430 381922 291498 381978
rect 291554 381922 291622 381978
rect 291678 381922 291774 381978
rect 291154 364350 291774 381922
rect 291154 364294 291250 364350
rect 291306 364294 291374 364350
rect 291430 364294 291498 364350
rect 291554 364294 291622 364350
rect 291678 364294 291774 364350
rect 291154 364226 291774 364294
rect 291154 364170 291250 364226
rect 291306 364170 291374 364226
rect 291430 364170 291498 364226
rect 291554 364170 291622 364226
rect 291678 364170 291774 364226
rect 291154 364102 291774 364170
rect 291154 364046 291250 364102
rect 291306 364046 291374 364102
rect 291430 364046 291498 364102
rect 291554 364046 291622 364102
rect 291678 364046 291774 364102
rect 291154 363978 291774 364046
rect 291154 363922 291250 363978
rect 291306 363922 291374 363978
rect 291430 363922 291498 363978
rect 291554 363922 291622 363978
rect 291678 363922 291774 363978
rect 291154 346350 291774 363922
rect 291154 346294 291250 346350
rect 291306 346294 291374 346350
rect 291430 346294 291498 346350
rect 291554 346294 291622 346350
rect 291678 346294 291774 346350
rect 291154 346226 291774 346294
rect 291154 346170 291250 346226
rect 291306 346170 291374 346226
rect 291430 346170 291498 346226
rect 291554 346170 291622 346226
rect 291678 346170 291774 346226
rect 291154 346102 291774 346170
rect 291154 346046 291250 346102
rect 291306 346046 291374 346102
rect 291430 346046 291498 346102
rect 291554 346046 291622 346102
rect 291678 346046 291774 346102
rect 291154 345978 291774 346046
rect 291154 345922 291250 345978
rect 291306 345922 291374 345978
rect 291430 345922 291498 345978
rect 291554 345922 291622 345978
rect 291678 345922 291774 345978
rect 291154 328350 291774 345922
rect 291154 328294 291250 328350
rect 291306 328294 291374 328350
rect 291430 328294 291498 328350
rect 291554 328294 291622 328350
rect 291678 328294 291774 328350
rect 291154 328226 291774 328294
rect 291154 328170 291250 328226
rect 291306 328170 291374 328226
rect 291430 328170 291498 328226
rect 291554 328170 291622 328226
rect 291678 328170 291774 328226
rect 291154 328102 291774 328170
rect 291154 328046 291250 328102
rect 291306 328046 291374 328102
rect 291430 328046 291498 328102
rect 291554 328046 291622 328102
rect 291678 328046 291774 328102
rect 291154 327978 291774 328046
rect 291154 327922 291250 327978
rect 291306 327922 291374 327978
rect 291430 327922 291498 327978
rect 291554 327922 291622 327978
rect 291678 327922 291774 327978
rect 291154 310350 291774 327922
rect 291154 310294 291250 310350
rect 291306 310294 291374 310350
rect 291430 310294 291498 310350
rect 291554 310294 291622 310350
rect 291678 310294 291774 310350
rect 291154 310226 291774 310294
rect 291154 310170 291250 310226
rect 291306 310170 291374 310226
rect 291430 310170 291498 310226
rect 291554 310170 291622 310226
rect 291678 310170 291774 310226
rect 291154 310102 291774 310170
rect 291154 310046 291250 310102
rect 291306 310046 291374 310102
rect 291430 310046 291498 310102
rect 291554 310046 291622 310102
rect 291678 310046 291774 310102
rect 291154 309978 291774 310046
rect 291154 309922 291250 309978
rect 291306 309922 291374 309978
rect 291430 309922 291498 309978
rect 291554 309922 291622 309978
rect 291678 309922 291774 309978
rect 291154 292350 291774 309922
rect 291154 292294 291250 292350
rect 291306 292294 291374 292350
rect 291430 292294 291498 292350
rect 291554 292294 291622 292350
rect 291678 292294 291774 292350
rect 291154 292226 291774 292294
rect 291154 292170 291250 292226
rect 291306 292170 291374 292226
rect 291430 292170 291498 292226
rect 291554 292170 291622 292226
rect 291678 292170 291774 292226
rect 291154 292102 291774 292170
rect 291154 292046 291250 292102
rect 291306 292046 291374 292102
rect 291430 292046 291498 292102
rect 291554 292046 291622 292102
rect 291678 292046 291774 292102
rect 291154 291978 291774 292046
rect 291154 291922 291250 291978
rect 291306 291922 291374 291978
rect 291430 291922 291498 291978
rect 291554 291922 291622 291978
rect 291678 291922 291774 291978
rect 291154 274350 291774 291922
rect 291154 274294 291250 274350
rect 291306 274294 291374 274350
rect 291430 274294 291498 274350
rect 291554 274294 291622 274350
rect 291678 274294 291774 274350
rect 291154 274226 291774 274294
rect 291154 274170 291250 274226
rect 291306 274170 291374 274226
rect 291430 274170 291498 274226
rect 291554 274170 291622 274226
rect 291678 274170 291774 274226
rect 291154 274102 291774 274170
rect 291154 274046 291250 274102
rect 291306 274046 291374 274102
rect 291430 274046 291498 274102
rect 291554 274046 291622 274102
rect 291678 274046 291774 274102
rect 291154 273978 291774 274046
rect 291154 273922 291250 273978
rect 291306 273922 291374 273978
rect 291430 273922 291498 273978
rect 291554 273922 291622 273978
rect 291678 273922 291774 273978
rect 291154 256350 291774 273922
rect 291154 256294 291250 256350
rect 291306 256294 291374 256350
rect 291430 256294 291498 256350
rect 291554 256294 291622 256350
rect 291678 256294 291774 256350
rect 291154 256226 291774 256294
rect 291154 256170 291250 256226
rect 291306 256170 291374 256226
rect 291430 256170 291498 256226
rect 291554 256170 291622 256226
rect 291678 256170 291774 256226
rect 291154 256102 291774 256170
rect 291154 256046 291250 256102
rect 291306 256046 291374 256102
rect 291430 256046 291498 256102
rect 291554 256046 291622 256102
rect 291678 256046 291774 256102
rect 291154 255978 291774 256046
rect 291154 255922 291250 255978
rect 291306 255922 291374 255978
rect 291430 255922 291498 255978
rect 291554 255922 291622 255978
rect 291678 255922 291774 255978
rect 291154 238350 291774 255922
rect 309154 597212 309774 598268
rect 309154 597156 309250 597212
rect 309306 597156 309374 597212
rect 309430 597156 309498 597212
rect 309554 597156 309622 597212
rect 309678 597156 309774 597212
rect 309154 597088 309774 597156
rect 309154 597032 309250 597088
rect 309306 597032 309374 597088
rect 309430 597032 309498 597088
rect 309554 597032 309622 597088
rect 309678 597032 309774 597088
rect 309154 596964 309774 597032
rect 309154 596908 309250 596964
rect 309306 596908 309374 596964
rect 309430 596908 309498 596964
rect 309554 596908 309622 596964
rect 309678 596908 309774 596964
rect 309154 596840 309774 596908
rect 309154 596784 309250 596840
rect 309306 596784 309374 596840
rect 309430 596784 309498 596840
rect 309554 596784 309622 596840
rect 309678 596784 309774 596840
rect 309154 580350 309774 596784
rect 309154 580294 309250 580350
rect 309306 580294 309374 580350
rect 309430 580294 309498 580350
rect 309554 580294 309622 580350
rect 309678 580294 309774 580350
rect 309154 580226 309774 580294
rect 309154 580170 309250 580226
rect 309306 580170 309374 580226
rect 309430 580170 309498 580226
rect 309554 580170 309622 580226
rect 309678 580170 309774 580226
rect 309154 580102 309774 580170
rect 309154 580046 309250 580102
rect 309306 580046 309374 580102
rect 309430 580046 309498 580102
rect 309554 580046 309622 580102
rect 309678 580046 309774 580102
rect 309154 579978 309774 580046
rect 309154 579922 309250 579978
rect 309306 579922 309374 579978
rect 309430 579922 309498 579978
rect 309554 579922 309622 579978
rect 309678 579922 309774 579978
rect 309154 562350 309774 579922
rect 309154 562294 309250 562350
rect 309306 562294 309374 562350
rect 309430 562294 309498 562350
rect 309554 562294 309622 562350
rect 309678 562294 309774 562350
rect 309154 562226 309774 562294
rect 309154 562170 309250 562226
rect 309306 562170 309374 562226
rect 309430 562170 309498 562226
rect 309554 562170 309622 562226
rect 309678 562170 309774 562226
rect 309154 562102 309774 562170
rect 309154 562046 309250 562102
rect 309306 562046 309374 562102
rect 309430 562046 309498 562102
rect 309554 562046 309622 562102
rect 309678 562046 309774 562102
rect 309154 561978 309774 562046
rect 309154 561922 309250 561978
rect 309306 561922 309374 561978
rect 309430 561922 309498 561978
rect 309554 561922 309622 561978
rect 309678 561922 309774 561978
rect 309154 544350 309774 561922
rect 309154 544294 309250 544350
rect 309306 544294 309374 544350
rect 309430 544294 309498 544350
rect 309554 544294 309622 544350
rect 309678 544294 309774 544350
rect 309154 544226 309774 544294
rect 309154 544170 309250 544226
rect 309306 544170 309374 544226
rect 309430 544170 309498 544226
rect 309554 544170 309622 544226
rect 309678 544170 309774 544226
rect 309154 544102 309774 544170
rect 309154 544046 309250 544102
rect 309306 544046 309374 544102
rect 309430 544046 309498 544102
rect 309554 544046 309622 544102
rect 309678 544046 309774 544102
rect 309154 543978 309774 544046
rect 309154 543922 309250 543978
rect 309306 543922 309374 543978
rect 309430 543922 309498 543978
rect 309554 543922 309622 543978
rect 309678 543922 309774 543978
rect 309154 526350 309774 543922
rect 309154 526294 309250 526350
rect 309306 526294 309374 526350
rect 309430 526294 309498 526350
rect 309554 526294 309622 526350
rect 309678 526294 309774 526350
rect 309154 526226 309774 526294
rect 309154 526170 309250 526226
rect 309306 526170 309374 526226
rect 309430 526170 309498 526226
rect 309554 526170 309622 526226
rect 309678 526170 309774 526226
rect 309154 526102 309774 526170
rect 309154 526046 309250 526102
rect 309306 526046 309374 526102
rect 309430 526046 309498 526102
rect 309554 526046 309622 526102
rect 309678 526046 309774 526102
rect 309154 525978 309774 526046
rect 309154 525922 309250 525978
rect 309306 525922 309374 525978
rect 309430 525922 309498 525978
rect 309554 525922 309622 525978
rect 309678 525922 309774 525978
rect 309154 508350 309774 525922
rect 309154 508294 309250 508350
rect 309306 508294 309374 508350
rect 309430 508294 309498 508350
rect 309554 508294 309622 508350
rect 309678 508294 309774 508350
rect 309154 508226 309774 508294
rect 309154 508170 309250 508226
rect 309306 508170 309374 508226
rect 309430 508170 309498 508226
rect 309554 508170 309622 508226
rect 309678 508170 309774 508226
rect 309154 508102 309774 508170
rect 309154 508046 309250 508102
rect 309306 508046 309374 508102
rect 309430 508046 309498 508102
rect 309554 508046 309622 508102
rect 309678 508046 309774 508102
rect 309154 507978 309774 508046
rect 309154 507922 309250 507978
rect 309306 507922 309374 507978
rect 309430 507922 309498 507978
rect 309554 507922 309622 507978
rect 309678 507922 309774 507978
rect 309154 490350 309774 507922
rect 309154 490294 309250 490350
rect 309306 490294 309374 490350
rect 309430 490294 309498 490350
rect 309554 490294 309622 490350
rect 309678 490294 309774 490350
rect 309154 490226 309774 490294
rect 309154 490170 309250 490226
rect 309306 490170 309374 490226
rect 309430 490170 309498 490226
rect 309554 490170 309622 490226
rect 309678 490170 309774 490226
rect 309154 490102 309774 490170
rect 309154 490046 309250 490102
rect 309306 490046 309374 490102
rect 309430 490046 309498 490102
rect 309554 490046 309622 490102
rect 309678 490046 309774 490102
rect 309154 489978 309774 490046
rect 309154 489922 309250 489978
rect 309306 489922 309374 489978
rect 309430 489922 309498 489978
rect 309554 489922 309622 489978
rect 309678 489922 309774 489978
rect 309154 472350 309774 489922
rect 309154 472294 309250 472350
rect 309306 472294 309374 472350
rect 309430 472294 309498 472350
rect 309554 472294 309622 472350
rect 309678 472294 309774 472350
rect 309154 472226 309774 472294
rect 309154 472170 309250 472226
rect 309306 472170 309374 472226
rect 309430 472170 309498 472226
rect 309554 472170 309622 472226
rect 309678 472170 309774 472226
rect 309154 472102 309774 472170
rect 309154 472046 309250 472102
rect 309306 472046 309374 472102
rect 309430 472046 309498 472102
rect 309554 472046 309622 472102
rect 309678 472046 309774 472102
rect 309154 471978 309774 472046
rect 309154 471922 309250 471978
rect 309306 471922 309374 471978
rect 309430 471922 309498 471978
rect 309554 471922 309622 471978
rect 309678 471922 309774 471978
rect 309154 454350 309774 471922
rect 309154 454294 309250 454350
rect 309306 454294 309374 454350
rect 309430 454294 309498 454350
rect 309554 454294 309622 454350
rect 309678 454294 309774 454350
rect 309154 454226 309774 454294
rect 309154 454170 309250 454226
rect 309306 454170 309374 454226
rect 309430 454170 309498 454226
rect 309554 454170 309622 454226
rect 309678 454170 309774 454226
rect 309154 454102 309774 454170
rect 309154 454046 309250 454102
rect 309306 454046 309374 454102
rect 309430 454046 309498 454102
rect 309554 454046 309622 454102
rect 309678 454046 309774 454102
rect 309154 453978 309774 454046
rect 309154 453922 309250 453978
rect 309306 453922 309374 453978
rect 309430 453922 309498 453978
rect 309554 453922 309622 453978
rect 309678 453922 309774 453978
rect 309154 436350 309774 453922
rect 309154 436294 309250 436350
rect 309306 436294 309374 436350
rect 309430 436294 309498 436350
rect 309554 436294 309622 436350
rect 309678 436294 309774 436350
rect 309154 436226 309774 436294
rect 309154 436170 309250 436226
rect 309306 436170 309374 436226
rect 309430 436170 309498 436226
rect 309554 436170 309622 436226
rect 309678 436170 309774 436226
rect 309154 436102 309774 436170
rect 309154 436046 309250 436102
rect 309306 436046 309374 436102
rect 309430 436046 309498 436102
rect 309554 436046 309622 436102
rect 309678 436046 309774 436102
rect 309154 435978 309774 436046
rect 309154 435922 309250 435978
rect 309306 435922 309374 435978
rect 309430 435922 309498 435978
rect 309554 435922 309622 435978
rect 309678 435922 309774 435978
rect 309154 418350 309774 435922
rect 309154 418294 309250 418350
rect 309306 418294 309374 418350
rect 309430 418294 309498 418350
rect 309554 418294 309622 418350
rect 309678 418294 309774 418350
rect 309154 418226 309774 418294
rect 309154 418170 309250 418226
rect 309306 418170 309374 418226
rect 309430 418170 309498 418226
rect 309554 418170 309622 418226
rect 309678 418170 309774 418226
rect 309154 418102 309774 418170
rect 309154 418046 309250 418102
rect 309306 418046 309374 418102
rect 309430 418046 309498 418102
rect 309554 418046 309622 418102
rect 309678 418046 309774 418102
rect 309154 417978 309774 418046
rect 309154 417922 309250 417978
rect 309306 417922 309374 417978
rect 309430 417922 309498 417978
rect 309554 417922 309622 417978
rect 309678 417922 309774 417978
rect 309154 400350 309774 417922
rect 309154 400294 309250 400350
rect 309306 400294 309374 400350
rect 309430 400294 309498 400350
rect 309554 400294 309622 400350
rect 309678 400294 309774 400350
rect 309154 400226 309774 400294
rect 309154 400170 309250 400226
rect 309306 400170 309374 400226
rect 309430 400170 309498 400226
rect 309554 400170 309622 400226
rect 309678 400170 309774 400226
rect 309154 400102 309774 400170
rect 309154 400046 309250 400102
rect 309306 400046 309374 400102
rect 309430 400046 309498 400102
rect 309554 400046 309622 400102
rect 309678 400046 309774 400102
rect 309154 399978 309774 400046
rect 309154 399922 309250 399978
rect 309306 399922 309374 399978
rect 309430 399922 309498 399978
rect 309554 399922 309622 399978
rect 309678 399922 309774 399978
rect 309154 382350 309774 399922
rect 309154 382294 309250 382350
rect 309306 382294 309374 382350
rect 309430 382294 309498 382350
rect 309554 382294 309622 382350
rect 309678 382294 309774 382350
rect 309154 382226 309774 382294
rect 309154 382170 309250 382226
rect 309306 382170 309374 382226
rect 309430 382170 309498 382226
rect 309554 382170 309622 382226
rect 309678 382170 309774 382226
rect 309154 382102 309774 382170
rect 309154 382046 309250 382102
rect 309306 382046 309374 382102
rect 309430 382046 309498 382102
rect 309554 382046 309622 382102
rect 309678 382046 309774 382102
rect 309154 381978 309774 382046
rect 309154 381922 309250 381978
rect 309306 381922 309374 381978
rect 309430 381922 309498 381978
rect 309554 381922 309622 381978
rect 309678 381922 309774 381978
rect 309154 364350 309774 381922
rect 309154 364294 309250 364350
rect 309306 364294 309374 364350
rect 309430 364294 309498 364350
rect 309554 364294 309622 364350
rect 309678 364294 309774 364350
rect 309154 364226 309774 364294
rect 309154 364170 309250 364226
rect 309306 364170 309374 364226
rect 309430 364170 309498 364226
rect 309554 364170 309622 364226
rect 309678 364170 309774 364226
rect 309154 364102 309774 364170
rect 309154 364046 309250 364102
rect 309306 364046 309374 364102
rect 309430 364046 309498 364102
rect 309554 364046 309622 364102
rect 309678 364046 309774 364102
rect 309154 363978 309774 364046
rect 309154 363922 309250 363978
rect 309306 363922 309374 363978
rect 309430 363922 309498 363978
rect 309554 363922 309622 363978
rect 309678 363922 309774 363978
rect 309154 346350 309774 363922
rect 309154 346294 309250 346350
rect 309306 346294 309374 346350
rect 309430 346294 309498 346350
rect 309554 346294 309622 346350
rect 309678 346294 309774 346350
rect 309154 346226 309774 346294
rect 309154 346170 309250 346226
rect 309306 346170 309374 346226
rect 309430 346170 309498 346226
rect 309554 346170 309622 346226
rect 309678 346170 309774 346226
rect 309154 346102 309774 346170
rect 309154 346046 309250 346102
rect 309306 346046 309374 346102
rect 309430 346046 309498 346102
rect 309554 346046 309622 346102
rect 309678 346046 309774 346102
rect 309154 345978 309774 346046
rect 309154 345922 309250 345978
rect 309306 345922 309374 345978
rect 309430 345922 309498 345978
rect 309554 345922 309622 345978
rect 309678 345922 309774 345978
rect 309154 328350 309774 345922
rect 309154 328294 309250 328350
rect 309306 328294 309374 328350
rect 309430 328294 309498 328350
rect 309554 328294 309622 328350
rect 309678 328294 309774 328350
rect 309154 328226 309774 328294
rect 309154 328170 309250 328226
rect 309306 328170 309374 328226
rect 309430 328170 309498 328226
rect 309554 328170 309622 328226
rect 309678 328170 309774 328226
rect 309154 328102 309774 328170
rect 309154 328046 309250 328102
rect 309306 328046 309374 328102
rect 309430 328046 309498 328102
rect 309554 328046 309622 328102
rect 309678 328046 309774 328102
rect 309154 327978 309774 328046
rect 309154 327922 309250 327978
rect 309306 327922 309374 327978
rect 309430 327922 309498 327978
rect 309554 327922 309622 327978
rect 309678 327922 309774 327978
rect 309154 310350 309774 327922
rect 309154 310294 309250 310350
rect 309306 310294 309374 310350
rect 309430 310294 309498 310350
rect 309554 310294 309622 310350
rect 309678 310294 309774 310350
rect 309154 310226 309774 310294
rect 309154 310170 309250 310226
rect 309306 310170 309374 310226
rect 309430 310170 309498 310226
rect 309554 310170 309622 310226
rect 309678 310170 309774 310226
rect 309154 310102 309774 310170
rect 309154 310046 309250 310102
rect 309306 310046 309374 310102
rect 309430 310046 309498 310102
rect 309554 310046 309622 310102
rect 309678 310046 309774 310102
rect 309154 309978 309774 310046
rect 309154 309922 309250 309978
rect 309306 309922 309374 309978
rect 309430 309922 309498 309978
rect 309554 309922 309622 309978
rect 309678 309922 309774 309978
rect 309154 292350 309774 309922
rect 309154 292294 309250 292350
rect 309306 292294 309374 292350
rect 309430 292294 309498 292350
rect 309554 292294 309622 292350
rect 309678 292294 309774 292350
rect 309154 292226 309774 292294
rect 309154 292170 309250 292226
rect 309306 292170 309374 292226
rect 309430 292170 309498 292226
rect 309554 292170 309622 292226
rect 309678 292170 309774 292226
rect 309154 292102 309774 292170
rect 309154 292046 309250 292102
rect 309306 292046 309374 292102
rect 309430 292046 309498 292102
rect 309554 292046 309622 292102
rect 309678 292046 309774 292102
rect 309154 291978 309774 292046
rect 309154 291922 309250 291978
rect 309306 291922 309374 291978
rect 309430 291922 309498 291978
rect 309554 291922 309622 291978
rect 309678 291922 309774 291978
rect 309154 274350 309774 291922
rect 309154 274294 309250 274350
rect 309306 274294 309374 274350
rect 309430 274294 309498 274350
rect 309554 274294 309622 274350
rect 309678 274294 309774 274350
rect 309154 274226 309774 274294
rect 309154 274170 309250 274226
rect 309306 274170 309374 274226
rect 309430 274170 309498 274226
rect 309554 274170 309622 274226
rect 309678 274170 309774 274226
rect 309154 274102 309774 274170
rect 309154 274046 309250 274102
rect 309306 274046 309374 274102
rect 309430 274046 309498 274102
rect 309554 274046 309622 274102
rect 309678 274046 309774 274102
rect 309154 273978 309774 274046
rect 309154 273922 309250 273978
rect 309306 273922 309374 273978
rect 309430 273922 309498 273978
rect 309554 273922 309622 273978
rect 309678 273922 309774 273978
rect 309154 256350 309774 273922
rect 309154 256294 309250 256350
rect 309306 256294 309374 256350
rect 309430 256294 309498 256350
rect 309554 256294 309622 256350
rect 309678 256294 309774 256350
rect 309154 256226 309774 256294
rect 309154 256170 309250 256226
rect 309306 256170 309374 256226
rect 309430 256170 309498 256226
rect 309554 256170 309622 256226
rect 309678 256170 309774 256226
rect 309154 256102 309774 256170
rect 309154 256046 309250 256102
rect 309306 256046 309374 256102
rect 309430 256046 309498 256102
rect 309554 256046 309622 256102
rect 309678 256046 309774 256102
rect 309154 255978 309774 256046
rect 309154 255922 309250 255978
rect 309306 255922 309374 255978
rect 309430 255922 309498 255978
rect 309554 255922 309622 255978
rect 309678 255922 309774 255978
rect 291154 238294 291250 238350
rect 291306 238294 291374 238350
rect 291430 238294 291498 238350
rect 291554 238294 291622 238350
rect 291678 238294 291774 238350
rect 291154 238226 291774 238294
rect 291154 238170 291250 238226
rect 291306 238170 291374 238226
rect 291430 238170 291498 238226
rect 291554 238170 291622 238226
rect 291678 238170 291774 238226
rect 291154 238102 291774 238170
rect 291154 238046 291250 238102
rect 291306 238046 291374 238102
rect 291430 238046 291498 238102
rect 291554 238046 291622 238102
rect 291678 238046 291774 238102
rect 291154 237978 291774 238046
rect 291154 237922 291250 237978
rect 291306 237922 291374 237978
rect 291430 237922 291498 237978
rect 291554 237922 291622 237978
rect 291678 237922 291774 237978
rect 291154 220350 291774 237922
rect 291154 220294 291250 220350
rect 291306 220294 291374 220350
rect 291430 220294 291498 220350
rect 291554 220294 291622 220350
rect 291678 220294 291774 220350
rect 291154 220226 291774 220294
rect 291154 220170 291250 220226
rect 291306 220170 291374 220226
rect 291430 220170 291498 220226
rect 291554 220170 291622 220226
rect 291678 220170 291774 220226
rect 291154 220102 291774 220170
rect 291154 220046 291250 220102
rect 291306 220046 291374 220102
rect 291430 220046 291498 220102
rect 291554 220046 291622 220102
rect 291678 220046 291774 220102
rect 291154 219978 291774 220046
rect 291154 219922 291250 219978
rect 291306 219922 291374 219978
rect 291430 219922 291498 219978
rect 291554 219922 291622 219978
rect 291678 219922 291774 219978
rect 291154 202350 291774 219922
rect 291154 202294 291250 202350
rect 291306 202294 291374 202350
rect 291430 202294 291498 202350
rect 291554 202294 291622 202350
rect 291678 202294 291774 202350
rect 291154 202226 291774 202294
rect 291154 202170 291250 202226
rect 291306 202170 291374 202226
rect 291430 202170 291498 202226
rect 291554 202170 291622 202226
rect 291678 202170 291774 202226
rect 291154 202102 291774 202170
rect 291154 202046 291250 202102
rect 291306 202046 291374 202102
rect 291430 202046 291498 202102
rect 291554 202046 291622 202102
rect 291678 202046 291774 202102
rect 291154 201978 291774 202046
rect 291154 201922 291250 201978
rect 291306 201922 291374 201978
rect 291430 201922 291498 201978
rect 291554 201922 291622 201978
rect 291678 201922 291774 201978
rect 291154 184350 291774 201922
rect 291154 184294 291250 184350
rect 291306 184294 291374 184350
rect 291430 184294 291498 184350
rect 291554 184294 291622 184350
rect 291678 184294 291774 184350
rect 291154 184226 291774 184294
rect 291154 184170 291250 184226
rect 291306 184170 291374 184226
rect 291430 184170 291498 184226
rect 291554 184170 291622 184226
rect 291678 184170 291774 184226
rect 291154 184102 291774 184170
rect 291154 184046 291250 184102
rect 291306 184046 291374 184102
rect 291430 184046 291498 184102
rect 291554 184046 291622 184102
rect 291678 184046 291774 184102
rect 291154 183978 291774 184046
rect 291154 183922 291250 183978
rect 291306 183922 291374 183978
rect 291430 183922 291498 183978
rect 291554 183922 291622 183978
rect 291678 183922 291774 183978
rect 283988 166412 285228 166446
rect 283988 166356 284022 166412
rect 284078 166356 284146 166412
rect 284202 166356 284270 166412
rect 284326 166356 284394 166412
rect 284450 166356 284518 166412
rect 284574 166356 284642 166412
rect 284698 166356 284766 166412
rect 284822 166356 284890 166412
rect 284946 166356 285014 166412
rect 285070 166356 285138 166412
rect 285194 166356 285228 166412
rect 283988 166288 285228 166356
rect 283988 166232 284022 166288
rect 284078 166232 284146 166288
rect 284202 166232 284270 166288
rect 284326 166232 284394 166288
rect 284450 166232 284518 166288
rect 284574 166232 284642 166288
rect 284698 166232 284766 166288
rect 284822 166232 284890 166288
rect 284946 166232 285014 166288
rect 285070 166232 285138 166288
rect 285194 166232 285228 166288
rect 283988 166164 285228 166232
rect 283988 166108 284022 166164
rect 284078 166108 284146 166164
rect 284202 166108 284270 166164
rect 284326 166108 284394 166164
rect 284450 166108 284518 166164
rect 284574 166108 284642 166164
rect 284698 166108 284766 166164
rect 284822 166108 284890 166164
rect 284946 166108 285014 166164
rect 285070 166108 285138 166164
rect 285194 166108 285228 166164
rect 283988 166040 285228 166108
rect 283988 165984 284022 166040
rect 284078 165984 284146 166040
rect 284202 165984 284270 166040
rect 284326 165984 284394 166040
rect 284450 165984 284518 166040
rect 284574 165984 284642 166040
rect 284698 165984 284766 166040
rect 284822 165984 284890 166040
rect 284946 165984 285014 166040
rect 285070 165984 285138 166040
rect 285194 165984 285228 166040
rect 283988 165916 285228 165984
rect 283988 165860 284022 165916
rect 284078 165860 284146 165916
rect 284202 165860 284270 165916
rect 284326 165860 284394 165916
rect 284450 165860 284518 165916
rect 284574 165860 284642 165916
rect 284698 165860 284766 165916
rect 284822 165860 284890 165916
rect 284946 165860 285014 165916
rect 285070 165860 285138 165916
rect 285194 165860 285228 165916
rect 283988 165826 285228 165860
rect 291154 166350 291774 183922
rect 294874 226350 295494 242964
rect 294874 226294 294970 226350
rect 295026 226294 295094 226350
rect 295150 226294 295218 226350
rect 295274 226294 295342 226350
rect 295398 226294 295494 226350
rect 294874 226226 295494 226294
rect 294874 226170 294970 226226
rect 295026 226170 295094 226226
rect 295150 226170 295218 226226
rect 295274 226170 295342 226226
rect 295398 226170 295494 226226
rect 294874 226102 295494 226170
rect 294874 226046 294970 226102
rect 295026 226046 295094 226102
rect 295150 226046 295218 226102
rect 295274 226046 295342 226102
rect 295398 226046 295494 226102
rect 294874 225978 295494 226046
rect 294874 225922 294970 225978
rect 295026 225922 295094 225978
rect 295150 225922 295218 225978
rect 295274 225922 295342 225978
rect 295398 225922 295494 225978
rect 294874 208350 295494 225922
rect 294874 208294 294970 208350
rect 295026 208294 295094 208350
rect 295150 208294 295218 208350
rect 295274 208294 295342 208350
rect 295398 208294 295494 208350
rect 294874 208226 295494 208294
rect 294874 208170 294970 208226
rect 295026 208170 295094 208226
rect 295150 208170 295218 208226
rect 295274 208170 295342 208226
rect 295398 208170 295494 208226
rect 294874 208102 295494 208170
rect 294874 208046 294970 208102
rect 295026 208046 295094 208102
rect 295150 208046 295218 208102
rect 295274 208046 295342 208102
rect 295398 208046 295494 208102
rect 294874 207978 295494 208046
rect 294874 207922 294970 207978
rect 295026 207922 295094 207978
rect 295150 207922 295218 207978
rect 295274 207922 295342 207978
rect 295398 207922 295494 207978
rect 294874 190350 295494 207922
rect 294874 190294 294970 190350
rect 295026 190294 295094 190350
rect 295150 190294 295218 190350
rect 295274 190294 295342 190350
rect 295398 190294 295494 190350
rect 294874 190226 295494 190294
rect 294874 190170 294970 190226
rect 295026 190170 295094 190226
rect 295150 190170 295218 190226
rect 295274 190170 295342 190226
rect 295398 190170 295494 190226
rect 294874 190102 295494 190170
rect 294874 190046 294970 190102
rect 295026 190046 295094 190102
rect 295150 190046 295218 190102
rect 295274 190046 295342 190102
rect 295398 190046 295494 190102
rect 294874 189978 295494 190046
rect 294874 189922 294970 189978
rect 295026 189922 295094 189978
rect 295150 189922 295218 189978
rect 295274 189922 295342 189978
rect 295398 189922 295494 189978
rect 294874 172350 295494 189922
rect 294874 172294 294970 172350
rect 295026 172294 295094 172350
rect 295150 172294 295218 172350
rect 295274 172294 295342 172350
rect 295398 172294 295494 172350
rect 294874 172226 295494 172294
rect 294874 172170 294970 172226
rect 295026 172170 295094 172226
rect 295150 172170 295218 172226
rect 295274 172170 295342 172226
rect 295398 172170 295494 172226
rect 294874 172102 295494 172170
rect 294874 172046 294970 172102
rect 295026 172046 295094 172102
rect 295150 172046 295218 172102
rect 295274 172046 295342 172102
rect 295398 172046 295494 172102
rect 294874 171978 295494 172046
rect 294874 171922 294970 171978
rect 295026 171922 295094 171978
rect 295150 171922 295218 171978
rect 295274 171922 295342 171978
rect 295398 171922 295494 171978
rect 294874 168604 295494 171922
rect 309154 238350 309774 255922
rect 309154 238294 309250 238350
rect 309306 238294 309374 238350
rect 309430 238294 309498 238350
rect 309554 238294 309622 238350
rect 309678 238294 309774 238350
rect 309154 238226 309774 238294
rect 309154 238170 309250 238226
rect 309306 238170 309374 238226
rect 309430 238170 309498 238226
rect 309554 238170 309622 238226
rect 309678 238170 309774 238226
rect 309154 238102 309774 238170
rect 309154 238046 309250 238102
rect 309306 238046 309374 238102
rect 309430 238046 309498 238102
rect 309554 238046 309622 238102
rect 309678 238046 309774 238102
rect 309154 237978 309774 238046
rect 309154 237922 309250 237978
rect 309306 237922 309374 237978
rect 309430 237922 309498 237978
rect 309554 237922 309622 237978
rect 309678 237922 309774 237978
rect 309154 220350 309774 237922
rect 309154 220294 309250 220350
rect 309306 220294 309374 220350
rect 309430 220294 309498 220350
rect 309554 220294 309622 220350
rect 309678 220294 309774 220350
rect 309154 220226 309774 220294
rect 309154 220170 309250 220226
rect 309306 220170 309374 220226
rect 309430 220170 309498 220226
rect 309554 220170 309622 220226
rect 309678 220170 309774 220226
rect 309154 220102 309774 220170
rect 309154 220046 309250 220102
rect 309306 220046 309374 220102
rect 309430 220046 309498 220102
rect 309554 220046 309622 220102
rect 309678 220046 309774 220102
rect 309154 219978 309774 220046
rect 309154 219922 309250 219978
rect 309306 219922 309374 219978
rect 309430 219922 309498 219978
rect 309554 219922 309622 219978
rect 309678 219922 309774 219978
rect 309154 202350 309774 219922
rect 309154 202294 309250 202350
rect 309306 202294 309374 202350
rect 309430 202294 309498 202350
rect 309554 202294 309622 202350
rect 309678 202294 309774 202350
rect 309154 202226 309774 202294
rect 309154 202170 309250 202226
rect 309306 202170 309374 202226
rect 309430 202170 309498 202226
rect 309554 202170 309622 202226
rect 309678 202170 309774 202226
rect 309154 202102 309774 202170
rect 309154 202046 309250 202102
rect 309306 202046 309374 202102
rect 309430 202046 309498 202102
rect 309554 202046 309622 202102
rect 309678 202046 309774 202102
rect 309154 201978 309774 202046
rect 309154 201922 309250 201978
rect 309306 201922 309374 201978
rect 309430 201922 309498 201978
rect 309554 201922 309622 201978
rect 309678 201922 309774 201978
rect 309154 184350 309774 201922
rect 309154 184294 309250 184350
rect 309306 184294 309374 184350
rect 309430 184294 309498 184350
rect 309554 184294 309622 184350
rect 309678 184294 309774 184350
rect 309154 184226 309774 184294
rect 309154 184170 309250 184226
rect 309306 184170 309374 184226
rect 309430 184170 309498 184226
rect 309554 184170 309622 184226
rect 309678 184170 309774 184226
rect 309154 184102 309774 184170
rect 309154 184046 309250 184102
rect 309306 184046 309374 184102
rect 309430 184046 309498 184102
rect 309554 184046 309622 184102
rect 309678 184046 309774 184102
rect 309154 183978 309774 184046
rect 309154 183922 309250 183978
rect 309306 183922 309374 183978
rect 309430 183922 309498 183978
rect 309554 183922 309622 183978
rect 309678 183922 309774 183978
rect 291154 166294 291250 166350
rect 291306 166294 291374 166350
rect 291430 166294 291498 166350
rect 291554 166294 291622 166350
rect 291678 166294 291774 166350
rect 291154 166226 291774 166294
rect 291154 166170 291250 166226
rect 291306 166170 291374 166226
rect 291430 166170 291498 166226
rect 291554 166170 291622 166226
rect 291678 166170 291774 166226
rect 291154 166102 291774 166170
rect 291154 166046 291250 166102
rect 291306 166046 291374 166102
rect 291430 166046 291498 166102
rect 291554 166046 291622 166102
rect 291678 166046 291774 166102
rect 291154 165978 291774 166046
rect 291154 165922 291250 165978
rect 291306 165922 291374 165978
rect 291430 165922 291498 165978
rect 291554 165922 291622 165978
rect 291678 165922 291774 165978
rect 291154 158782 291774 165922
rect 303988 166412 305228 166446
rect 303988 166356 304022 166412
rect 304078 166356 304146 166412
rect 304202 166356 304270 166412
rect 304326 166356 304394 166412
rect 304450 166356 304518 166412
rect 304574 166356 304642 166412
rect 304698 166356 304766 166412
rect 304822 166356 304890 166412
rect 304946 166356 305014 166412
rect 305070 166356 305138 166412
rect 305194 166356 305228 166412
rect 303988 166288 305228 166356
rect 303988 166232 304022 166288
rect 304078 166232 304146 166288
rect 304202 166232 304270 166288
rect 304326 166232 304394 166288
rect 304450 166232 304518 166288
rect 304574 166232 304642 166288
rect 304698 166232 304766 166288
rect 304822 166232 304890 166288
rect 304946 166232 305014 166288
rect 305070 166232 305138 166288
rect 305194 166232 305228 166288
rect 303988 166164 305228 166232
rect 303988 166108 304022 166164
rect 304078 166108 304146 166164
rect 304202 166108 304270 166164
rect 304326 166108 304394 166164
rect 304450 166108 304518 166164
rect 304574 166108 304642 166164
rect 304698 166108 304766 166164
rect 304822 166108 304890 166164
rect 304946 166108 305014 166164
rect 305070 166108 305138 166164
rect 305194 166108 305228 166164
rect 303988 166040 305228 166108
rect 303988 165984 304022 166040
rect 304078 165984 304146 166040
rect 304202 165984 304270 166040
rect 304326 165984 304394 166040
rect 304450 165984 304518 166040
rect 304574 165984 304642 166040
rect 304698 165984 304766 166040
rect 304822 165984 304890 166040
rect 304946 165984 305014 166040
rect 305070 165984 305138 166040
rect 305194 165984 305228 166040
rect 303988 165916 305228 165984
rect 303988 165860 304022 165916
rect 304078 165860 304146 165916
rect 304202 165860 304270 165916
rect 304326 165860 304394 165916
rect 304450 165860 304518 165916
rect 304574 165860 304642 165916
rect 304698 165860 304766 165916
rect 304822 165860 304890 165916
rect 304946 165860 305014 165916
rect 305070 165860 305138 165916
rect 305194 165860 305228 165916
rect 303988 165826 305228 165860
rect 309154 166350 309774 183922
rect 309154 166294 309250 166350
rect 309306 166294 309374 166350
rect 309430 166294 309498 166350
rect 309554 166294 309622 166350
rect 309678 166294 309774 166350
rect 309154 166226 309774 166294
rect 309154 166170 309250 166226
rect 309306 166170 309374 166226
rect 309430 166170 309498 166226
rect 309554 166170 309622 166226
rect 309678 166170 309774 166226
rect 309154 166102 309774 166170
rect 309154 166046 309250 166102
rect 309306 166046 309374 166102
rect 309430 166046 309498 166102
rect 309554 166046 309622 166102
rect 309678 166046 309774 166102
rect 309154 165978 309774 166046
rect 309154 165922 309250 165978
rect 309306 165922 309374 165978
rect 309430 165922 309498 165978
rect 309554 165922 309622 165978
rect 309678 165922 309774 165978
rect 309154 158782 309774 165922
rect 312874 598172 313494 598268
rect 312874 598116 312970 598172
rect 313026 598116 313094 598172
rect 313150 598116 313218 598172
rect 313274 598116 313342 598172
rect 313398 598116 313494 598172
rect 312874 598048 313494 598116
rect 312874 597992 312970 598048
rect 313026 597992 313094 598048
rect 313150 597992 313218 598048
rect 313274 597992 313342 598048
rect 313398 597992 313494 598048
rect 312874 597924 313494 597992
rect 312874 597868 312970 597924
rect 313026 597868 313094 597924
rect 313150 597868 313218 597924
rect 313274 597868 313342 597924
rect 313398 597868 313494 597924
rect 312874 597800 313494 597868
rect 312874 597744 312970 597800
rect 313026 597744 313094 597800
rect 313150 597744 313218 597800
rect 313274 597744 313342 597800
rect 313398 597744 313494 597800
rect 312874 586350 313494 597744
rect 312874 586294 312970 586350
rect 313026 586294 313094 586350
rect 313150 586294 313218 586350
rect 313274 586294 313342 586350
rect 313398 586294 313494 586350
rect 312874 586226 313494 586294
rect 312874 586170 312970 586226
rect 313026 586170 313094 586226
rect 313150 586170 313218 586226
rect 313274 586170 313342 586226
rect 313398 586170 313494 586226
rect 312874 586102 313494 586170
rect 312874 586046 312970 586102
rect 313026 586046 313094 586102
rect 313150 586046 313218 586102
rect 313274 586046 313342 586102
rect 313398 586046 313494 586102
rect 312874 585978 313494 586046
rect 312874 585922 312970 585978
rect 313026 585922 313094 585978
rect 313150 585922 313218 585978
rect 313274 585922 313342 585978
rect 313398 585922 313494 585978
rect 312874 568350 313494 585922
rect 312874 568294 312970 568350
rect 313026 568294 313094 568350
rect 313150 568294 313218 568350
rect 313274 568294 313342 568350
rect 313398 568294 313494 568350
rect 312874 568226 313494 568294
rect 312874 568170 312970 568226
rect 313026 568170 313094 568226
rect 313150 568170 313218 568226
rect 313274 568170 313342 568226
rect 313398 568170 313494 568226
rect 312874 568102 313494 568170
rect 312874 568046 312970 568102
rect 313026 568046 313094 568102
rect 313150 568046 313218 568102
rect 313274 568046 313342 568102
rect 313398 568046 313494 568102
rect 312874 567978 313494 568046
rect 312874 567922 312970 567978
rect 313026 567922 313094 567978
rect 313150 567922 313218 567978
rect 313274 567922 313342 567978
rect 313398 567922 313494 567978
rect 312874 550350 313494 567922
rect 312874 550294 312970 550350
rect 313026 550294 313094 550350
rect 313150 550294 313218 550350
rect 313274 550294 313342 550350
rect 313398 550294 313494 550350
rect 312874 550226 313494 550294
rect 312874 550170 312970 550226
rect 313026 550170 313094 550226
rect 313150 550170 313218 550226
rect 313274 550170 313342 550226
rect 313398 550170 313494 550226
rect 312874 550102 313494 550170
rect 312874 550046 312970 550102
rect 313026 550046 313094 550102
rect 313150 550046 313218 550102
rect 313274 550046 313342 550102
rect 313398 550046 313494 550102
rect 312874 549978 313494 550046
rect 312874 549922 312970 549978
rect 313026 549922 313094 549978
rect 313150 549922 313218 549978
rect 313274 549922 313342 549978
rect 313398 549922 313494 549978
rect 312874 532350 313494 549922
rect 312874 532294 312970 532350
rect 313026 532294 313094 532350
rect 313150 532294 313218 532350
rect 313274 532294 313342 532350
rect 313398 532294 313494 532350
rect 312874 532226 313494 532294
rect 312874 532170 312970 532226
rect 313026 532170 313094 532226
rect 313150 532170 313218 532226
rect 313274 532170 313342 532226
rect 313398 532170 313494 532226
rect 312874 532102 313494 532170
rect 312874 532046 312970 532102
rect 313026 532046 313094 532102
rect 313150 532046 313218 532102
rect 313274 532046 313342 532102
rect 313398 532046 313494 532102
rect 312874 531978 313494 532046
rect 312874 531922 312970 531978
rect 313026 531922 313094 531978
rect 313150 531922 313218 531978
rect 313274 531922 313342 531978
rect 313398 531922 313494 531978
rect 312874 514350 313494 531922
rect 312874 514294 312970 514350
rect 313026 514294 313094 514350
rect 313150 514294 313218 514350
rect 313274 514294 313342 514350
rect 313398 514294 313494 514350
rect 312874 514226 313494 514294
rect 312874 514170 312970 514226
rect 313026 514170 313094 514226
rect 313150 514170 313218 514226
rect 313274 514170 313342 514226
rect 313398 514170 313494 514226
rect 312874 514102 313494 514170
rect 312874 514046 312970 514102
rect 313026 514046 313094 514102
rect 313150 514046 313218 514102
rect 313274 514046 313342 514102
rect 313398 514046 313494 514102
rect 312874 513978 313494 514046
rect 312874 513922 312970 513978
rect 313026 513922 313094 513978
rect 313150 513922 313218 513978
rect 313274 513922 313342 513978
rect 313398 513922 313494 513978
rect 312874 496350 313494 513922
rect 312874 496294 312970 496350
rect 313026 496294 313094 496350
rect 313150 496294 313218 496350
rect 313274 496294 313342 496350
rect 313398 496294 313494 496350
rect 312874 496226 313494 496294
rect 312874 496170 312970 496226
rect 313026 496170 313094 496226
rect 313150 496170 313218 496226
rect 313274 496170 313342 496226
rect 313398 496170 313494 496226
rect 312874 496102 313494 496170
rect 312874 496046 312970 496102
rect 313026 496046 313094 496102
rect 313150 496046 313218 496102
rect 313274 496046 313342 496102
rect 313398 496046 313494 496102
rect 312874 495978 313494 496046
rect 312874 495922 312970 495978
rect 313026 495922 313094 495978
rect 313150 495922 313218 495978
rect 313274 495922 313342 495978
rect 313398 495922 313494 495978
rect 312874 478350 313494 495922
rect 312874 478294 312970 478350
rect 313026 478294 313094 478350
rect 313150 478294 313218 478350
rect 313274 478294 313342 478350
rect 313398 478294 313494 478350
rect 312874 478226 313494 478294
rect 312874 478170 312970 478226
rect 313026 478170 313094 478226
rect 313150 478170 313218 478226
rect 313274 478170 313342 478226
rect 313398 478170 313494 478226
rect 312874 478102 313494 478170
rect 312874 478046 312970 478102
rect 313026 478046 313094 478102
rect 313150 478046 313218 478102
rect 313274 478046 313342 478102
rect 313398 478046 313494 478102
rect 312874 477978 313494 478046
rect 312874 477922 312970 477978
rect 313026 477922 313094 477978
rect 313150 477922 313218 477978
rect 313274 477922 313342 477978
rect 313398 477922 313494 477978
rect 312874 460350 313494 477922
rect 312874 460294 312970 460350
rect 313026 460294 313094 460350
rect 313150 460294 313218 460350
rect 313274 460294 313342 460350
rect 313398 460294 313494 460350
rect 312874 460226 313494 460294
rect 312874 460170 312970 460226
rect 313026 460170 313094 460226
rect 313150 460170 313218 460226
rect 313274 460170 313342 460226
rect 313398 460170 313494 460226
rect 312874 460102 313494 460170
rect 312874 460046 312970 460102
rect 313026 460046 313094 460102
rect 313150 460046 313218 460102
rect 313274 460046 313342 460102
rect 313398 460046 313494 460102
rect 312874 459978 313494 460046
rect 312874 459922 312970 459978
rect 313026 459922 313094 459978
rect 313150 459922 313218 459978
rect 313274 459922 313342 459978
rect 313398 459922 313494 459978
rect 312874 442350 313494 459922
rect 312874 442294 312970 442350
rect 313026 442294 313094 442350
rect 313150 442294 313218 442350
rect 313274 442294 313342 442350
rect 313398 442294 313494 442350
rect 312874 442226 313494 442294
rect 312874 442170 312970 442226
rect 313026 442170 313094 442226
rect 313150 442170 313218 442226
rect 313274 442170 313342 442226
rect 313398 442170 313494 442226
rect 312874 442102 313494 442170
rect 312874 442046 312970 442102
rect 313026 442046 313094 442102
rect 313150 442046 313218 442102
rect 313274 442046 313342 442102
rect 313398 442046 313494 442102
rect 312874 441978 313494 442046
rect 312874 441922 312970 441978
rect 313026 441922 313094 441978
rect 313150 441922 313218 441978
rect 313274 441922 313342 441978
rect 313398 441922 313494 441978
rect 312874 424350 313494 441922
rect 312874 424294 312970 424350
rect 313026 424294 313094 424350
rect 313150 424294 313218 424350
rect 313274 424294 313342 424350
rect 313398 424294 313494 424350
rect 312874 424226 313494 424294
rect 312874 424170 312970 424226
rect 313026 424170 313094 424226
rect 313150 424170 313218 424226
rect 313274 424170 313342 424226
rect 313398 424170 313494 424226
rect 312874 424102 313494 424170
rect 312874 424046 312970 424102
rect 313026 424046 313094 424102
rect 313150 424046 313218 424102
rect 313274 424046 313342 424102
rect 313398 424046 313494 424102
rect 312874 423978 313494 424046
rect 312874 423922 312970 423978
rect 313026 423922 313094 423978
rect 313150 423922 313218 423978
rect 313274 423922 313342 423978
rect 313398 423922 313494 423978
rect 312874 406350 313494 423922
rect 312874 406294 312970 406350
rect 313026 406294 313094 406350
rect 313150 406294 313218 406350
rect 313274 406294 313342 406350
rect 313398 406294 313494 406350
rect 312874 406226 313494 406294
rect 312874 406170 312970 406226
rect 313026 406170 313094 406226
rect 313150 406170 313218 406226
rect 313274 406170 313342 406226
rect 313398 406170 313494 406226
rect 312874 406102 313494 406170
rect 312874 406046 312970 406102
rect 313026 406046 313094 406102
rect 313150 406046 313218 406102
rect 313274 406046 313342 406102
rect 313398 406046 313494 406102
rect 312874 405978 313494 406046
rect 312874 405922 312970 405978
rect 313026 405922 313094 405978
rect 313150 405922 313218 405978
rect 313274 405922 313342 405978
rect 313398 405922 313494 405978
rect 312874 388350 313494 405922
rect 312874 388294 312970 388350
rect 313026 388294 313094 388350
rect 313150 388294 313218 388350
rect 313274 388294 313342 388350
rect 313398 388294 313494 388350
rect 312874 388226 313494 388294
rect 312874 388170 312970 388226
rect 313026 388170 313094 388226
rect 313150 388170 313218 388226
rect 313274 388170 313342 388226
rect 313398 388170 313494 388226
rect 312874 388102 313494 388170
rect 312874 388046 312970 388102
rect 313026 388046 313094 388102
rect 313150 388046 313218 388102
rect 313274 388046 313342 388102
rect 313398 388046 313494 388102
rect 312874 387978 313494 388046
rect 312874 387922 312970 387978
rect 313026 387922 313094 387978
rect 313150 387922 313218 387978
rect 313274 387922 313342 387978
rect 313398 387922 313494 387978
rect 312874 370350 313494 387922
rect 312874 370294 312970 370350
rect 313026 370294 313094 370350
rect 313150 370294 313218 370350
rect 313274 370294 313342 370350
rect 313398 370294 313494 370350
rect 312874 370226 313494 370294
rect 312874 370170 312970 370226
rect 313026 370170 313094 370226
rect 313150 370170 313218 370226
rect 313274 370170 313342 370226
rect 313398 370170 313494 370226
rect 312874 370102 313494 370170
rect 312874 370046 312970 370102
rect 313026 370046 313094 370102
rect 313150 370046 313218 370102
rect 313274 370046 313342 370102
rect 313398 370046 313494 370102
rect 312874 369978 313494 370046
rect 312874 369922 312970 369978
rect 313026 369922 313094 369978
rect 313150 369922 313218 369978
rect 313274 369922 313342 369978
rect 313398 369922 313494 369978
rect 312874 352350 313494 369922
rect 312874 352294 312970 352350
rect 313026 352294 313094 352350
rect 313150 352294 313218 352350
rect 313274 352294 313342 352350
rect 313398 352294 313494 352350
rect 312874 352226 313494 352294
rect 312874 352170 312970 352226
rect 313026 352170 313094 352226
rect 313150 352170 313218 352226
rect 313274 352170 313342 352226
rect 313398 352170 313494 352226
rect 312874 352102 313494 352170
rect 312874 352046 312970 352102
rect 313026 352046 313094 352102
rect 313150 352046 313218 352102
rect 313274 352046 313342 352102
rect 313398 352046 313494 352102
rect 312874 351978 313494 352046
rect 312874 351922 312970 351978
rect 313026 351922 313094 351978
rect 313150 351922 313218 351978
rect 313274 351922 313342 351978
rect 313398 351922 313494 351978
rect 312874 334350 313494 351922
rect 312874 334294 312970 334350
rect 313026 334294 313094 334350
rect 313150 334294 313218 334350
rect 313274 334294 313342 334350
rect 313398 334294 313494 334350
rect 312874 334226 313494 334294
rect 312874 334170 312970 334226
rect 313026 334170 313094 334226
rect 313150 334170 313218 334226
rect 313274 334170 313342 334226
rect 313398 334170 313494 334226
rect 312874 334102 313494 334170
rect 312874 334046 312970 334102
rect 313026 334046 313094 334102
rect 313150 334046 313218 334102
rect 313274 334046 313342 334102
rect 313398 334046 313494 334102
rect 312874 333978 313494 334046
rect 312874 333922 312970 333978
rect 313026 333922 313094 333978
rect 313150 333922 313218 333978
rect 313274 333922 313342 333978
rect 313398 333922 313494 333978
rect 312874 316350 313494 333922
rect 312874 316294 312970 316350
rect 313026 316294 313094 316350
rect 313150 316294 313218 316350
rect 313274 316294 313342 316350
rect 313398 316294 313494 316350
rect 312874 316226 313494 316294
rect 312874 316170 312970 316226
rect 313026 316170 313094 316226
rect 313150 316170 313218 316226
rect 313274 316170 313342 316226
rect 313398 316170 313494 316226
rect 312874 316102 313494 316170
rect 312874 316046 312970 316102
rect 313026 316046 313094 316102
rect 313150 316046 313218 316102
rect 313274 316046 313342 316102
rect 313398 316046 313494 316102
rect 312874 315978 313494 316046
rect 312874 315922 312970 315978
rect 313026 315922 313094 315978
rect 313150 315922 313218 315978
rect 313274 315922 313342 315978
rect 313398 315922 313494 315978
rect 312874 298350 313494 315922
rect 312874 298294 312970 298350
rect 313026 298294 313094 298350
rect 313150 298294 313218 298350
rect 313274 298294 313342 298350
rect 313398 298294 313494 298350
rect 312874 298226 313494 298294
rect 312874 298170 312970 298226
rect 313026 298170 313094 298226
rect 313150 298170 313218 298226
rect 313274 298170 313342 298226
rect 313398 298170 313494 298226
rect 312874 298102 313494 298170
rect 312874 298046 312970 298102
rect 313026 298046 313094 298102
rect 313150 298046 313218 298102
rect 313274 298046 313342 298102
rect 313398 298046 313494 298102
rect 312874 297978 313494 298046
rect 312874 297922 312970 297978
rect 313026 297922 313094 297978
rect 313150 297922 313218 297978
rect 313274 297922 313342 297978
rect 313398 297922 313494 297978
rect 312874 280350 313494 297922
rect 312874 280294 312970 280350
rect 313026 280294 313094 280350
rect 313150 280294 313218 280350
rect 313274 280294 313342 280350
rect 313398 280294 313494 280350
rect 312874 280226 313494 280294
rect 312874 280170 312970 280226
rect 313026 280170 313094 280226
rect 313150 280170 313218 280226
rect 313274 280170 313342 280226
rect 313398 280170 313494 280226
rect 312874 280102 313494 280170
rect 312874 280046 312970 280102
rect 313026 280046 313094 280102
rect 313150 280046 313218 280102
rect 313274 280046 313342 280102
rect 313398 280046 313494 280102
rect 312874 279978 313494 280046
rect 312874 279922 312970 279978
rect 313026 279922 313094 279978
rect 313150 279922 313218 279978
rect 313274 279922 313342 279978
rect 313398 279922 313494 279978
rect 312874 262350 313494 279922
rect 312874 262294 312970 262350
rect 313026 262294 313094 262350
rect 313150 262294 313218 262350
rect 313274 262294 313342 262350
rect 313398 262294 313494 262350
rect 312874 262226 313494 262294
rect 312874 262170 312970 262226
rect 313026 262170 313094 262226
rect 313150 262170 313218 262226
rect 313274 262170 313342 262226
rect 313398 262170 313494 262226
rect 312874 262102 313494 262170
rect 312874 262046 312970 262102
rect 313026 262046 313094 262102
rect 313150 262046 313218 262102
rect 313274 262046 313342 262102
rect 313398 262046 313494 262102
rect 312874 261978 313494 262046
rect 312874 261922 312970 261978
rect 313026 261922 313094 261978
rect 313150 261922 313218 261978
rect 313274 261922 313342 261978
rect 313398 261922 313494 261978
rect 312874 244350 313494 261922
rect 312874 244294 312970 244350
rect 313026 244294 313094 244350
rect 313150 244294 313218 244350
rect 313274 244294 313342 244350
rect 313398 244294 313494 244350
rect 312874 244226 313494 244294
rect 312874 244170 312970 244226
rect 313026 244170 313094 244226
rect 313150 244170 313218 244226
rect 313274 244170 313342 244226
rect 313398 244170 313494 244226
rect 312874 244102 313494 244170
rect 312874 244046 312970 244102
rect 313026 244046 313094 244102
rect 313150 244046 313218 244102
rect 313274 244046 313342 244102
rect 313398 244046 313494 244102
rect 312874 243978 313494 244046
rect 312874 243922 312970 243978
rect 313026 243922 313094 243978
rect 313150 243922 313218 243978
rect 313274 243922 313342 243978
rect 313398 243922 313494 243978
rect 312874 226350 313494 243922
rect 312874 226294 312970 226350
rect 313026 226294 313094 226350
rect 313150 226294 313218 226350
rect 313274 226294 313342 226350
rect 313398 226294 313494 226350
rect 312874 226226 313494 226294
rect 312874 226170 312970 226226
rect 313026 226170 313094 226226
rect 313150 226170 313218 226226
rect 313274 226170 313342 226226
rect 313398 226170 313494 226226
rect 312874 226102 313494 226170
rect 312874 226046 312970 226102
rect 313026 226046 313094 226102
rect 313150 226046 313218 226102
rect 313274 226046 313342 226102
rect 313398 226046 313494 226102
rect 312874 225978 313494 226046
rect 312874 225922 312970 225978
rect 313026 225922 313094 225978
rect 313150 225922 313218 225978
rect 313274 225922 313342 225978
rect 313398 225922 313494 225978
rect 312874 208350 313494 225922
rect 312874 208294 312970 208350
rect 313026 208294 313094 208350
rect 313150 208294 313218 208350
rect 313274 208294 313342 208350
rect 313398 208294 313494 208350
rect 312874 208226 313494 208294
rect 312874 208170 312970 208226
rect 313026 208170 313094 208226
rect 313150 208170 313218 208226
rect 313274 208170 313342 208226
rect 313398 208170 313494 208226
rect 312874 208102 313494 208170
rect 312874 208046 312970 208102
rect 313026 208046 313094 208102
rect 313150 208046 313218 208102
rect 313274 208046 313342 208102
rect 313398 208046 313494 208102
rect 312874 207978 313494 208046
rect 312874 207922 312970 207978
rect 313026 207922 313094 207978
rect 313150 207922 313218 207978
rect 313274 207922 313342 207978
rect 313398 207922 313494 207978
rect 312874 190350 313494 207922
rect 312874 190294 312970 190350
rect 313026 190294 313094 190350
rect 313150 190294 313218 190350
rect 313274 190294 313342 190350
rect 313398 190294 313494 190350
rect 312874 190226 313494 190294
rect 312874 190170 312970 190226
rect 313026 190170 313094 190226
rect 313150 190170 313218 190226
rect 313274 190170 313342 190226
rect 313398 190170 313494 190226
rect 312874 190102 313494 190170
rect 312874 190046 312970 190102
rect 313026 190046 313094 190102
rect 313150 190046 313218 190102
rect 313274 190046 313342 190102
rect 313398 190046 313494 190102
rect 312874 189978 313494 190046
rect 312874 189922 312970 189978
rect 313026 189922 313094 189978
rect 313150 189922 313218 189978
rect 313274 189922 313342 189978
rect 313398 189922 313494 189978
rect 312874 172350 313494 189922
rect 312874 172294 312970 172350
rect 313026 172294 313094 172350
rect 313150 172294 313218 172350
rect 313274 172294 313342 172350
rect 313398 172294 313494 172350
rect 312874 172226 313494 172294
rect 312874 172170 312970 172226
rect 313026 172170 313094 172226
rect 313150 172170 313218 172226
rect 313274 172170 313342 172226
rect 313398 172170 313494 172226
rect 312874 172102 313494 172170
rect 312874 172046 312970 172102
rect 313026 172046 313094 172102
rect 313150 172046 313218 172102
rect 313274 172046 313342 172102
rect 313398 172046 313494 172102
rect 312874 171978 313494 172046
rect 312874 171922 312970 171978
rect 313026 171922 313094 171978
rect 313150 171922 313218 171978
rect 313274 171922 313342 171978
rect 313398 171922 313494 171978
rect 312874 158782 313494 171922
rect 327154 597212 327774 598268
rect 327154 597156 327250 597212
rect 327306 597156 327374 597212
rect 327430 597156 327498 597212
rect 327554 597156 327622 597212
rect 327678 597156 327774 597212
rect 327154 597088 327774 597156
rect 327154 597032 327250 597088
rect 327306 597032 327374 597088
rect 327430 597032 327498 597088
rect 327554 597032 327622 597088
rect 327678 597032 327774 597088
rect 327154 596964 327774 597032
rect 327154 596908 327250 596964
rect 327306 596908 327374 596964
rect 327430 596908 327498 596964
rect 327554 596908 327622 596964
rect 327678 596908 327774 596964
rect 327154 596840 327774 596908
rect 327154 596784 327250 596840
rect 327306 596784 327374 596840
rect 327430 596784 327498 596840
rect 327554 596784 327622 596840
rect 327678 596784 327774 596840
rect 327154 580350 327774 596784
rect 327154 580294 327250 580350
rect 327306 580294 327374 580350
rect 327430 580294 327498 580350
rect 327554 580294 327622 580350
rect 327678 580294 327774 580350
rect 327154 580226 327774 580294
rect 327154 580170 327250 580226
rect 327306 580170 327374 580226
rect 327430 580170 327498 580226
rect 327554 580170 327622 580226
rect 327678 580170 327774 580226
rect 327154 580102 327774 580170
rect 327154 580046 327250 580102
rect 327306 580046 327374 580102
rect 327430 580046 327498 580102
rect 327554 580046 327622 580102
rect 327678 580046 327774 580102
rect 327154 579978 327774 580046
rect 327154 579922 327250 579978
rect 327306 579922 327374 579978
rect 327430 579922 327498 579978
rect 327554 579922 327622 579978
rect 327678 579922 327774 579978
rect 327154 562350 327774 579922
rect 327154 562294 327250 562350
rect 327306 562294 327374 562350
rect 327430 562294 327498 562350
rect 327554 562294 327622 562350
rect 327678 562294 327774 562350
rect 327154 562226 327774 562294
rect 327154 562170 327250 562226
rect 327306 562170 327374 562226
rect 327430 562170 327498 562226
rect 327554 562170 327622 562226
rect 327678 562170 327774 562226
rect 327154 562102 327774 562170
rect 327154 562046 327250 562102
rect 327306 562046 327374 562102
rect 327430 562046 327498 562102
rect 327554 562046 327622 562102
rect 327678 562046 327774 562102
rect 327154 561978 327774 562046
rect 327154 561922 327250 561978
rect 327306 561922 327374 561978
rect 327430 561922 327498 561978
rect 327554 561922 327622 561978
rect 327678 561922 327774 561978
rect 327154 544350 327774 561922
rect 327154 544294 327250 544350
rect 327306 544294 327374 544350
rect 327430 544294 327498 544350
rect 327554 544294 327622 544350
rect 327678 544294 327774 544350
rect 327154 544226 327774 544294
rect 327154 544170 327250 544226
rect 327306 544170 327374 544226
rect 327430 544170 327498 544226
rect 327554 544170 327622 544226
rect 327678 544170 327774 544226
rect 327154 544102 327774 544170
rect 327154 544046 327250 544102
rect 327306 544046 327374 544102
rect 327430 544046 327498 544102
rect 327554 544046 327622 544102
rect 327678 544046 327774 544102
rect 327154 543978 327774 544046
rect 327154 543922 327250 543978
rect 327306 543922 327374 543978
rect 327430 543922 327498 543978
rect 327554 543922 327622 543978
rect 327678 543922 327774 543978
rect 327154 526350 327774 543922
rect 327154 526294 327250 526350
rect 327306 526294 327374 526350
rect 327430 526294 327498 526350
rect 327554 526294 327622 526350
rect 327678 526294 327774 526350
rect 327154 526226 327774 526294
rect 327154 526170 327250 526226
rect 327306 526170 327374 526226
rect 327430 526170 327498 526226
rect 327554 526170 327622 526226
rect 327678 526170 327774 526226
rect 327154 526102 327774 526170
rect 327154 526046 327250 526102
rect 327306 526046 327374 526102
rect 327430 526046 327498 526102
rect 327554 526046 327622 526102
rect 327678 526046 327774 526102
rect 327154 525978 327774 526046
rect 327154 525922 327250 525978
rect 327306 525922 327374 525978
rect 327430 525922 327498 525978
rect 327554 525922 327622 525978
rect 327678 525922 327774 525978
rect 327154 508350 327774 525922
rect 327154 508294 327250 508350
rect 327306 508294 327374 508350
rect 327430 508294 327498 508350
rect 327554 508294 327622 508350
rect 327678 508294 327774 508350
rect 327154 508226 327774 508294
rect 327154 508170 327250 508226
rect 327306 508170 327374 508226
rect 327430 508170 327498 508226
rect 327554 508170 327622 508226
rect 327678 508170 327774 508226
rect 327154 508102 327774 508170
rect 327154 508046 327250 508102
rect 327306 508046 327374 508102
rect 327430 508046 327498 508102
rect 327554 508046 327622 508102
rect 327678 508046 327774 508102
rect 327154 507978 327774 508046
rect 327154 507922 327250 507978
rect 327306 507922 327374 507978
rect 327430 507922 327498 507978
rect 327554 507922 327622 507978
rect 327678 507922 327774 507978
rect 327154 490350 327774 507922
rect 327154 490294 327250 490350
rect 327306 490294 327374 490350
rect 327430 490294 327498 490350
rect 327554 490294 327622 490350
rect 327678 490294 327774 490350
rect 327154 490226 327774 490294
rect 327154 490170 327250 490226
rect 327306 490170 327374 490226
rect 327430 490170 327498 490226
rect 327554 490170 327622 490226
rect 327678 490170 327774 490226
rect 327154 490102 327774 490170
rect 327154 490046 327250 490102
rect 327306 490046 327374 490102
rect 327430 490046 327498 490102
rect 327554 490046 327622 490102
rect 327678 490046 327774 490102
rect 327154 489978 327774 490046
rect 327154 489922 327250 489978
rect 327306 489922 327374 489978
rect 327430 489922 327498 489978
rect 327554 489922 327622 489978
rect 327678 489922 327774 489978
rect 327154 472350 327774 489922
rect 327154 472294 327250 472350
rect 327306 472294 327374 472350
rect 327430 472294 327498 472350
rect 327554 472294 327622 472350
rect 327678 472294 327774 472350
rect 327154 472226 327774 472294
rect 327154 472170 327250 472226
rect 327306 472170 327374 472226
rect 327430 472170 327498 472226
rect 327554 472170 327622 472226
rect 327678 472170 327774 472226
rect 327154 472102 327774 472170
rect 327154 472046 327250 472102
rect 327306 472046 327374 472102
rect 327430 472046 327498 472102
rect 327554 472046 327622 472102
rect 327678 472046 327774 472102
rect 327154 471978 327774 472046
rect 327154 471922 327250 471978
rect 327306 471922 327374 471978
rect 327430 471922 327498 471978
rect 327554 471922 327622 471978
rect 327678 471922 327774 471978
rect 327154 454350 327774 471922
rect 327154 454294 327250 454350
rect 327306 454294 327374 454350
rect 327430 454294 327498 454350
rect 327554 454294 327622 454350
rect 327678 454294 327774 454350
rect 327154 454226 327774 454294
rect 327154 454170 327250 454226
rect 327306 454170 327374 454226
rect 327430 454170 327498 454226
rect 327554 454170 327622 454226
rect 327678 454170 327774 454226
rect 327154 454102 327774 454170
rect 327154 454046 327250 454102
rect 327306 454046 327374 454102
rect 327430 454046 327498 454102
rect 327554 454046 327622 454102
rect 327678 454046 327774 454102
rect 327154 453978 327774 454046
rect 327154 453922 327250 453978
rect 327306 453922 327374 453978
rect 327430 453922 327498 453978
rect 327554 453922 327622 453978
rect 327678 453922 327774 453978
rect 327154 436350 327774 453922
rect 327154 436294 327250 436350
rect 327306 436294 327374 436350
rect 327430 436294 327498 436350
rect 327554 436294 327622 436350
rect 327678 436294 327774 436350
rect 327154 436226 327774 436294
rect 327154 436170 327250 436226
rect 327306 436170 327374 436226
rect 327430 436170 327498 436226
rect 327554 436170 327622 436226
rect 327678 436170 327774 436226
rect 327154 436102 327774 436170
rect 327154 436046 327250 436102
rect 327306 436046 327374 436102
rect 327430 436046 327498 436102
rect 327554 436046 327622 436102
rect 327678 436046 327774 436102
rect 327154 435978 327774 436046
rect 327154 435922 327250 435978
rect 327306 435922 327374 435978
rect 327430 435922 327498 435978
rect 327554 435922 327622 435978
rect 327678 435922 327774 435978
rect 327154 418350 327774 435922
rect 327154 418294 327250 418350
rect 327306 418294 327374 418350
rect 327430 418294 327498 418350
rect 327554 418294 327622 418350
rect 327678 418294 327774 418350
rect 327154 418226 327774 418294
rect 327154 418170 327250 418226
rect 327306 418170 327374 418226
rect 327430 418170 327498 418226
rect 327554 418170 327622 418226
rect 327678 418170 327774 418226
rect 327154 418102 327774 418170
rect 327154 418046 327250 418102
rect 327306 418046 327374 418102
rect 327430 418046 327498 418102
rect 327554 418046 327622 418102
rect 327678 418046 327774 418102
rect 327154 417978 327774 418046
rect 327154 417922 327250 417978
rect 327306 417922 327374 417978
rect 327430 417922 327498 417978
rect 327554 417922 327622 417978
rect 327678 417922 327774 417978
rect 327154 400350 327774 417922
rect 327154 400294 327250 400350
rect 327306 400294 327374 400350
rect 327430 400294 327498 400350
rect 327554 400294 327622 400350
rect 327678 400294 327774 400350
rect 327154 400226 327774 400294
rect 327154 400170 327250 400226
rect 327306 400170 327374 400226
rect 327430 400170 327498 400226
rect 327554 400170 327622 400226
rect 327678 400170 327774 400226
rect 327154 400102 327774 400170
rect 327154 400046 327250 400102
rect 327306 400046 327374 400102
rect 327430 400046 327498 400102
rect 327554 400046 327622 400102
rect 327678 400046 327774 400102
rect 327154 399978 327774 400046
rect 327154 399922 327250 399978
rect 327306 399922 327374 399978
rect 327430 399922 327498 399978
rect 327554 399922 327622 399978
rect 327678 399922 327774 399978
rect 327154 382350 327774 399922
rect 327154 382294 327250 382350
rect 327306 382294 327374 382350
rect 327430 382294 327498 382350
rect 327554 382294 327622 382350
rect 327678 382294 327774 382350
rect 327154 382226 327774 382294
rect 327154 382170 327250 382226
rect 327306 382170 327374 382226
rect 327430 382170 327498 382226
rect 327554 382170 327622 382226
rect 327678 382170 327774 382226
rect 327154 382102 327774 382170
rect 327154 382046 327250 382102
rect 327306 382046 327374 382102
rect 327430 382046 327498 382102
rect 327554 382046 327622 382102
rect 327678 382046 327774 382102
rect 327154 381978 327774 382046
rect 327154 381922 327250 381978
rect 327306 381922 327374 381978
rect 327430 381922 327498 381978
rect 327554 381922 327622 381978
rect 327678 381922 327774 381978
rect 327154 364350 327774 381922
rect 327154 364294 327250 364350
rect 327306 364294 327374 364350
rect 327430 364294 327498 364350
rect 327554 364294 327622 364350
rect 327678 364294 327774 364350
rect 327154 364226 327774 364294
rect 327154 364170 327250 364226
rect 327306 364170 327374 364226
rect 327430 364170 327498 364226
rect 327554 364170 327622 364226
rect 327678 364170 327774 364226
rect 327154 364102 327774 364170
rect 327154 364046 327250 364102
rect 327306 364046 327374 364102
rect 327430 364046 327498 364102
rect 327554 364046 327622 364102
rect 327678 364046 327774 364102
rect 327154 363978 327774 364046
rect 327154 363922 327250 363978
rect 327306 363922 327374 363978
rect 327430 363922 327498 363978
rect 327554 363922 327622 363978
rect 327678 363922 327774 363978
rect 327154 346350 327774 363922
rect 327154 346294 327250 346350
rect 327306 346294 327374 346350
rect 327430 346294 327498 346350
rect 327554 346294 327622 346350
rect 327678 346294 327774 346350
rect 327154 346226 327774 346294
rect 327154 346170 327250 346226
rect 327306 346170 327374 346226
rect 327430 346170 327498 346226
rect 327554 346170 327622 346226
rect 327678 346170 327774 346226
rect 327154 346102 327774 346170
rect 327154 346046 327250 346102
rect 327306 346046 327374 346102
rect 327430 346046 327498 346102
rect 327554 346046 327622 346102
rect 327678 346046 327774 346102
rect 327154 345978 327774 346046
rect 327154 345922 327250 345978
rect 327306 345922 327374 345978
rect 327430 345922 327498 345978
rect 327554 345922 327622 345978
rect 327678 345922 327774 345978
rect 327154 328350 327774 345922
rect 327154 328294 327250 328350
rect 327306 328294 327374 328350
rect 327430 328294 327498 328350
rect 327554 328294 327622 328350
rect 327678 328294 327774 328350
rect 327154 328226 327774 328294
rect 327154 328170 327250 328226
rect 327306 328170 327374 328226
rect 327430 328170 327498 328226
rect 327554 328170 327622 328226
rect 327678 328170 327774 328226
rect 327154 328102 327774 328170
rect 327154 328046 327250 328102
rect 327306 328046 327374 328102
rect 327430 328046 327498 328102
rect 327554 328046 327622 328102
rect 327678 328046 327774 328102
rect 327154 327978 327774 328046
rect 327154 327922 327250 327978
rect 327306 327922 327374 327978
rect 327430 327922 327498 327978
rect 327554 327922 327622 327978
rect 327678 327922 327774 327978
rect 327154 310350 327774 327922
rect 327154 310294 327250 310350
rect 327306 310294 327374 310350
rect 327430 310294 327498 310350
rect 327554 310294 327622 310350
rect 327678 310294 327774 310350
rect 327154 310226 327774 310294
rect 327154 310170 327250 310226
rect 327306 310170 327374 310226
rect 327430 310170 327498 310226
rect 327554 310170 327622 310226
rect 327678 310170 327774 310226
rect 327154 310102 327774 310170
rect 327154 310046 327250 310102
rect 327306 310046 327374 310102
rect 327430 310046 327498 310102
rect 327554 310046 327622 310102
rect 327678 310046 327774 310102
rect 327154 309978 327774 310046
rect 327154 309922 327250 309978
rect 327306 309922 327374 309978
rect 327430 309922 327498 309978
rect 327554 309922 327622 309978
rect 327678 309922 327774 309978
rect 327154 292350 327774 309922
rect 327154 292294 327250 292350
rect 327306 292294 327374 292350
rect 327430 292294 327498 292350
rect 327554 292294 327622 292350
rect 327678 292294 327774 292350
rect 327154 292226 327774 292294
rect 327154 292170 327250 292226
rect 327306 292170 327374 292226
rect 327430 292170 327498 292226
rect 327554 292170 327622 292226
rect 327678 292170 327774 292226
rect 327154 292102 327774 292170
rect 327154 292046 327250 292102
rect 327306 292046 327374 292102
rect 327430 292046 327498 292102
rect 327554 292046 327622 292102
rect 327678 292046 327774 292102
rect 327154 291978 327774 292046
rect 327154 291922 327250 291978
rect 327306 291922 327374 291978
rect 327430 291922 327498 291978
rect 327554 291922 327622 291978
rect 327678 291922 327774 291978
rect 327154 274350 327774 291922
rect 327154 274294 327250 274350
rect 327306 274294 327374 274350
rect 327430 274294 327498 274350
rect 327554 274294 327622 274350
rect 327678 274294 327774 274350
rect 327154 274226 327774 274294
rect 327154 274170 327250 274226
rect 327306 274170 327374 274226
rect 327430 274170 327498 274226
rect 327554 274170 327622 274226
rect 327678 274170 327774 274226
rect 327154 274102 327774 274170
rect 327154 274046 327250 274102
rect 327306 274046 327374 274102
rect 327430 274046 327498 274102
rect 327554 274046 327622 274102
rect 327678 274046 327774 274102
rect 327154 273978 327774 274046
rect 327154 273922 327250 273978
rect 327306 273922 327374 273978
rect 327430 273922 327498 273978
rect 327554 273922 327622 273978
rect 327678 273922 327774 273978
rect 327154 256350 327774 273922
rect 327154 256294 327250 256350
rect 327306 256294 327374 256350
rect 327430 256294 327498 256350
rect 327554 256294 327622 256350
rect 327678 256294 327774 256350
rect 327154 256226 327774 256294
rect 327154 256170 327250 256226
rect 327306 256170 327374 256226
rect 327430 256170 327498 256226
rect 327554 256170 327622 256226
rect 327678 256170 327774 256226
rect 327154 256102 327774 256170
rect 327154 256046 327250 256102
rect 327306 256046 327374 256102
rect 327430 256046 327498 256102
rect 327554 256046 327622 256102
rect 327678 256046 327774 256102
rect 327154 255978 327774 256046
rect 327154 255922 327250 255978
rect 327306 255922 327374 255978
rect 327430 255922 327498 255978
rect 327554 255922 327622 255978
rect 327678 255922 327774 255978
rect 327154 238350 327774 255922
rect 327154 238294 327250 238350
rect 327306 238294 327374 238350
rect 327430 238294 327498 238350
rect 327554 238294 327622 238350
rect 327678 238294 327774 238350
rect 327154 238226 327774 238294
rect 327154 238170 327250 238226
rect 327306 238170 327374 238226
rect 327430 238170 327498 238226
rect 327554 238170 327622 238226
rect 327678 238170 327774 238226
rect 327154 238102 327774 238170
rect 327154 238046 327250 238102
rect 327306 238046 327374 238102
rect 327430 238046 327498 238102
rect 327554 238046 327622 238102
rect 327678 238046 327774 238102
rect 327154 237978 327774 238046
rect 327154 237922 327250 237978
rect 327306 237922 327374 237978
rect 327430 237922 327498 237978
rect 327554 237922 327622 237978
rect 327678 237922 327774 237978
rect 327154 220350 327774 237922
rect 327154 220294 327250 220350
rect 327306 220294 327374 220350
rect 327430 220294 327498 220350
rect 327554 220294 327622 220350
rect 327678 220294 327774 220350
rect 327154 220226 327774 220294
rect 327154 220170 327250 220226
rect 327306 220170 327374 220226
rect 327430 220170 327498 220226
rect 327554 220170 327622 220226
rect 327678 220170 327774 220226
rect 327154 220102 327774 220170
rect 327154 220046 327250 220102
rect 327306 220046 327374 220102
rect 327430 220046 327498 220102
rect 327554 220046 327622 220102
rect 327678 220046 327774 220102
rect 327154 219978 327774 220046
rect 327154 219922 327250 219978
rect 327306 219922 327374 219978
rect 327430 219922 327498 219978
rect 327554 219922 327622 219978
rect 327678 219922 327774 219978
rect 327154 202350 327774 219922
rect 327154 202294 327250 202350
rect 327306 202294 327374 202350
rect 327430 202294 327498 202350
rect 327554 202294 327622 202350
rect 327678 202294 327774 202350
rect 327154 202226 327774 202294
rect 327154 202170 327250 202226
rect 327306 202170 327374 202226
rect 327430 202170 327498 202226
rect 327554 202170 327622 202226
rect 327678 202170 327774 202226
rect 327154 202102 327774 202170
rect 327154 202046 327250 202102
rect 327306 202046 327374 202102
rect 327430 202046 327498 202102
rect 327554 202046 327622 202102
rect 327678 202046 327774 202102
rect 327154 201978 327774 202046
rect 327154 201922 327250 201978
rect 327306 201922 327374 201978
rect 327430 201922 327498 201978
rect 327554 201922 327622 201978
rect 327678 201922 327774 201978
rect 327154 184350 327774 201922
rect 327154 184294 327250 184350
rect 327306 184294 327374 184350
rect 327430 184294 327498 184350
rect 327554 184294 327622 184350
rect 327678 184294 327774 184350
rect 327154 184226 327774 184294
rect 327154 184170 327250 184226
rect 327306 184170 327374 184226
rect 327430 184170 327498 184226
rect 327554 184170 327622 184226
rect 327678 184170 327774 184226
rect 327154 184102 327774 184170
rect 327154 184046 327250 184102
rect 327306 184046 327374 184102
rect 327430 184046 327498 184102
rect 327554 184046 327622 184102
rect 327678 184046 327774 184102
rect 327154 183978 327774 184046
rect 327154 183922 327250 183978
rect 327306 183922 327374 183978
rect 327430 183922 327498 183978
rect 327554 183922 327622 183978
rect 327678 183922 327774 183978
rect 327154 166350 327774 183922
rect 327154 166294 327250 166350
rect 327306 166294 327374 166350
rect 327430 166294 327498 166350
rect 327554 166294 327622 166350
rect 327678 166294 327774 166350
rect 327154 166226 327774 166294
rect 327154 166170 327250 166226
rect 327306 166170 327374 166226
rect 327430 166170 327498 166226
rect 327554 166170 327622 166226
rect 327678 166170 327774 166226
rect 327154 166102 327774 166170
rect 327154 166046 327250 166102
rect 327306 166046 327374 166102
rect 327430 166046 327498 166102
rect 327554 166046 327622 166102
rect 327678 166046 327774 166102
rect 327154 165978 327774 166046
rect 327154 165922 327250 165978
rect 327306 165922 327374 165978
rect 327430 165922 327498 165978
rect 327554 165922 327622 165978
rect 327678 165922 327774 165978
rect 276874 154294 276970 154350
rect 277026 154294 277094 154350
rect 277150 154294 277218 154350
rect 277274 154294 277342 154350
rect 277398 154294 277494 154350
rect 276874 154226 277494 154294
rect 276874 154170 276970 154226
rect 277026 154170 277094 154226
rect 277150 154170 277218 154226
rect 277274 154170 277342 154226
rect 277398 154170 277494 154226
rect 276874 154102 277494 154170
rect 276874 154046 276970 154102
rect 277026 154046 277094 154102
rect 277150 154046 277218 154102
rect 277274 154046 277342 154102
rect 277398 154046 277494 154102
rect 274764 140578 274820 140588
rect 276874 153978 277494 154046
rect 276874 153922 276970 153978
rect 277026 153922 277094 153978
rect 277150 153922 277218 153978
rect 277274 153922 277342 153978
rect 277398 153922 277494 153978
rect 275548 138628 275604 138638
rect 275548 136164 275604 138572
rect 275548 136098 275604 136108
rect 276874 136350 277494 153922
rect 293988 154412 295228 154446
rect 293988 154356 294022 154412
rect 294078 154356 294146 154412
rect 294202 154356 294270 154412
rect 294326 154356 294394 154412
rect 294450 154356 294518 154412
rect 294574 154356 294642 154412
rect 294698 154356 294766 154412
rect 294822 154356 294890 154412
rect 294946 154356 295014 154412
rect 295070 154356 295138 154412
rect 295194 154356 295228 154412
rect 293988 154288 295228 154356
rect 293988 154232 294022 154288
rect 294078 154232 294146 154288
rect 294202 154232 294270 154288
rect 294326 154232 294394 154288
rect 294450 154232 294518 154288
rect 294574 154232 294642 154288
rect 294698 154232 294766 154288
rect 294822 154232 294890 154288
rect 294946 154232 295014 154288
rect 295070 154232 295138 154288
rect 295194 154232 295228 154288
rect 293988 154164 295228 154232
rect 293988 154108 294022 154164
rect 294078 154108 294146 154164
rect 294202 154108 294270 154164
rect 294326 154108 294394 154164
rect 294450 154108 294518 154164
rect 294574 154108 294642 154164
rect 294698 154108 294766 154164
rect 294822 154108 294890 154164
rect 294946 154108 295014 154164
rect 295070 154108 295138 154164
rect 295194 154108 295228 154164
rect 293988 154040 295228 154108
rect 293988 153984 294022 154040
rect 294078 153984 294146 154040
rect 294202 153984 294270 154040
rect 294326 153984 294394 154040
rect 294450 153984 294518 154040
rect 294574 153984 294642 154040
rect 294698 153984 294766 154040
rect 294822 153984 294890 154040
rect 294946 153984 295014 154040
rect 295070 153984 295138 154040
rect 295194 153984 295228 154040
rect 293988 153916 295228 153984
rect 293988 153860 294022 153916
rect 294078 153860 294146 153916
rect 294202 153860 294270 153916
rect 294326 153860 294394 153916
rect 294450 153860 294518 153916
rect 294574 153860 294642 153916
rect 294698 153860 294766 153916
rect 294822 153860 294890 153916
rect 294946 153860 295014 153916
rect 295070 153860 295138 153916
rect 295194 153860 295228 153916
rect 293988 153826 295228 153860
rect 313988 154412 315228 154446
rect 313988 154356 314022 154412
rect 314078 154356 314146 154412
rect 314202 154356 314270 154412
rect 314326 154356 314394 154412
rect 314450 154356 314518 154412
rect 314574 154356 314642 154412
rect 314698 154356 314766 154412
rect 314822 154356 314890 154412
rect 314946 154356 315014 154412
rect 315070 154356 315138 154412
rect 315194 154356 315228 154412
rect 313988 154288 315228 154356
rect 313988 154232 314022 154288
rect 314078 154232 314146 154288
rect 314202 154232 314270 154288
rect 314326 154232 314394 154288
rect 314450 154232 314518 154288
rect 314574 154232 314642 154288
rect 314698 154232 314766 154288
rect 314822 154232 314890 154288
rect 314946 154232 315014 154288
rect 315070 154232 315138 154288
rect 315194 154232 315228 154288
rect 313988 154164 315228 154232
rect 313988 154108 314022 154164
rect 314078 154108 314146 154164
rect 314202 154108 314270 154164
rect 314326 154108 314394 154164
rect 314450 154108 314518 154164
rect 314574 154108 314642 154164
rect 314698 154108 314766 154164
rect 314822 154108 314890 154164
rect 314946 154108 315014 154164
rect 315070 154108 315138 154164
rect 315194 154108 315228 154164
rect 313988 154040 315228 154108
rect 313988 153984 314022 154040
rect 314078 153984 314146 154040
rect 314202 153984 314270 154040
rect 314326 153984 314394 154040
rect 314450 153984 314518 154040
rect 314574 153984 314642 154040
rect 314698 153984 314766 154040
rect 314822 153984 314890 154040
rect 314946 153984 315014 154040
rect 315070 153984 315138 154040
rect 315194 153984 315228 154040
rect 313988 153916 315228 153984
rect 313988 153860 314022 153916
rect 314078 153860 314146 153916
rect 314202 153860 314270 153916
rect 314326 153860 314394 153916
rect 314450 153860 314518 153916
rect 314574 153860 314642 153916
rect 314698 153860 314766 153916
rect 314822 153860 314890 153916
rect 314946 153860 315014 153916
rect 315070 153860 315138 153916
rect 315194 153860 315228 153916
rect 313988 153826 315228 153860
rect 283988 148412 285228 148446
rect 283988 148356 284022 148412
rect 284078 148356 284146 148412
rect 284202 148356 284270 148412
rect 284326 148356 284394 148412
rect 284450 148356 284518 148412
rect 284574 148356 284642 148412
rect 284698 148356 284766 148412
rect 284822 148356 284890 148412
rect 284946 148356 285014 148412
rect 285070 148356 285138 148412
rect 285194 148356 285228 148412
rect 283988 148288 285228 148356
rect 283988 148232 284022 148288
rect 284078 148232 284146 148288
rect 284202 148232 284270 148288
rect 284326 148232 284394 148288
rect 284450 148232 284518 148288
rect 284574 148232 284642 148288
rect 284698 148232 284766 148288
rect 284822 148232 284890 148288
rect 284946 148232 285014 148288
rect 285070 148232 285138 148288
rect 285194 148232 285228 148288
rect 283988 148164 285228 148232
rect 283988 148108 284022 148164
rect 284078 148108 284146 148164
rect 284202 148108 284270 148164
rect 284326 148108 284394 148164
rect 284450 148108 284518 148164
rect 284574 148108 284642 148164
rect 284698 148108 284766 148164
rect 284822 148108 284890 148164
rect 284946 148108 285014 148164
rect 285070 148108 285138 148164
rect 285194 148108 285228 148164
rect 283988 148040 285228 148108
rect 283988 147984 284022 148040
rect 284078 147984 284146 148040
rect 284202 147984 284270 148040
rect 284326 147984 284394 148040
rect 284450 147984 284518 148040
rect 284574 147984 284642 148040
rect 284698 147984 284766 148040
rect 284822 147984 284890 148040
rect 284946 147984 285014 148040
rect 285070 147984 285138 148040
rect 285194 147984 285228 148040
rect 283988 147916 285228 147984
rect 283988 147860 284022 147916
rect 284078 147860 284146 147916
rect 284202 147860 284270 147916
rect 284326 147860 284394 147916
rect 284450 147860 284518 147916
rect 284574 147860 284642 147916
rect 284698 147860 284766 147916
rect 284822 147860 284890 147916
rect 284946 147860 285014 147916
rect 285070 147860 285138 147916
rect 285194 147860 285228 147916
rect 283988 147826 285228 147860
rect 303988 148412 305228 148446
rect 303988 148356 304022 148412
rect 304078 148356 304146 148412
rect 304202 148356 304270 148412
rect 304326 148356 304394 148412
rect 304450 148356 304518 148412
rect 304574 148356 304642 148412
rect 304698 148356 304766 148412
rect 304822 148356 304890 148412
rect 304946 148356 305014 148412
rect 305070 148356 305138 148412
rect 305194 148356 305228 148412
rect 303988 148288 305228 148356
rect 303988 148232 304022 148288
rect 304078 148232 304146 148288
rect 304202 148232 304270 148288
rect 304326 148232 304394 148288
rect 304450 148232 304518 148288
rect 304574 148232 304642 148288
rect 304698 148232 304766 148288
rect 304822 148232 304890 148288
rect 304946 148232 305014 148288
rect 305070 148232 305138 148288
rect 305194 148232 305228 148288
rect 303988 148164 305228 148232
rect 303988 148108 304022 148164
rect 304078 148108 304146 148164
rect 304202 148108 304270 148164
rect 304326 148108 304394 148164
rect 304450 148108 304518 148164
rect 304574 148108 304642 148164
rect 304698 148108 304766 148164
rect 304822 148108 304890 148164
rect 304946 148108 305014 148164
rect 305070 148108 305138 148164
rect 305194 148108 305228 148164
rect 303988 148040 305228 148108
rect 303988 147984 304022 148040
rect 304078 147984 304146 148040
rect 304202 147984 304270 148040
rect 304326 147984 304394 148040
rect 304450 147984 304518 148040
rect 304574 147984 304642 148040
rect 304698 147984 304766 148040
rect 304822 147984 304890 148040
rect 304946 147984 305014 148040
rect 305070 147984 305138 148040
rect 305194 147984 305228 148040
rect 303988 147916 305228 147984
rect 303988 147860 304022 147916
rect 304078 147860 304146 147916
rect 304202 147860 304270 147916
rect 304326 147860 304394 147916
rect 304450 147860 304518 147916
rect 304574 147860 304642 147916
rect 304698 147860 304766 147916
rect 304822 147860 304890 147916
rect 304946 147860 305014 147916
rect 305070 147860 305138 147916
rect 305194 147860 305228 147916
rect 303988 147826 305228 147860
rect 327154 148350 327774 165922
rect 327154 148294 327250 148350
rect 327306 148294 327374 148350
rect 327430 148294 327498 148350
rect 327554 148294 327622 148350
rect 327678 148294 327774 148350
rect 327154 148226 327774 148294
rect 327154 148170 327250 148226
rect 327306 148170 327374 148226
rect 327430 148170 327498 148226
rect 327554 148170 327622 148226
rect 327678 148170 327774 148226
rect 327154 148102 327774 148170
rect 327154 148046 327250 148102
rect 327306 148046 327374 148102
rect 327430 148046 327498 148102
rect 327554 148046 327622 148102
rect 327678 148046 327774 148102
rect 327154 147978 327774 148046
rect 327154 147922 327250 147978
rect 327306 147922 327374 147978
rect 327430 147922 327498 147978
rect 327554 147922 327622 147978
rect 327678 147922 327774 147978
rect 276874 136294 276970 136350
rect 277026 136294 277094 136350
rect 277150 136294 277218 136350
rect 277274 136294 277342 136350
rect 277398 136294 277494 136350
rect 276874 136226 277494 136294
rect 276874 136170 276970 136226
rect 277026 136170 277094 136226
rect 277150 136170 277218 136226
rect 277274 136170 277342 136226
rect 277398 136170 277494 136226
rect 276874 136102 277494 136170
rect 276874 136046 276970 136102
rect 277026 136046 277094 136102
rect 277150 136046 277218 136102
rect 277274 136046 277342 136102
rect 277398 136046 277494 136102
rect 276874 135978 277494 136046
rect 276874 135922 276970 135978
rect 277026 135922 277094 135978
rect 277150 135922 277218 135978
rect 277274 135922 277342 135978
rect 277398 135922 277494 135978
rect 275548 131908 275604 131918
rect 275548 130564 275604 131852
rect 275548 130498 275604 130508
rect 274652 129378 274708 129388
rect 275548 121828 275604 121838
rect 275548 118244 275604 121772
rect 275548 118178 275604 118188
rect 276874 118350 277494 135922
rect 293988 136412 295228 136446
rect 293988 136356 294022 136412
rect 294078 136356 294146 136412
rect 294202 136356 294270 136412
rect 294326 136356 294394 136412
rect 294450 136356 294518 136412
rect 294574 136356 294642 136412
rect 294698 136356 294766 136412
rect 294822 136356 294890 136412
rect 294946 136356 295014 136412
rect 295070 136356 295138 136412
rect 295194 136356 295228 136412
rect 293988 136288 295228 136356
rect 293988 136232 294022 136288
rect 294078 136232 294146 136288
rect 294202 136232 294270 136288
rect 294326 136232 294394 136288
rect 294450 136232 294518 136288
rect 294574 136232 294642 136288
rect 294698 136232 294766 136288
rect 294822 136232 294890 136288
rect 294946 136232 295014 136288
rect 295070 136232 295138 136288
rect 295194 136232 295228 136288
rect 293988 136164 295228 136232
rect 293988 136108 294022 136164
rect 294078 136108 294146 136164
rect 294202 136108 294270 136164
rect 294326 136108 294394 136164
rect 294450 136108 294518 136164
rect 294574 136108 294642 136164
rect 294698 136108 294766 136164
rect 294822 136108 294890 136164
rect 294946 136108 295014 136164
rect 295070 136108 295138 136164
rect 295194 136108 295228 136164
rect 293988 136040 295228 136108
rect 293988 135984 294022 136040
rect 294078 135984 294146 136040
rect 294202 135984 294270 136040
rect 294326 135984 294394 136040
rect 294450 135984 294518 136040
rect 294574 135984 294642 136040
rect 294698 135984 294766 136040
rect 294822 135984 294890 136040
rect 294946 135984 295014 136040
rect 295070 135984 295138 136040
rect 295194 135984 295228 136040
rect 293988 135916 295228 135984
rect 293988 135860 294022 135916
rect 294078 135860 294146 135916
rect 294202 135860 294270 135916
rect 294326 135860 294394 135916
rect 294450 135860 294518 135916
rect 294574 135860 294642 135916
rect 294698 135860 294766 135916
rect 294822 135860 294890 135916
rect 294946 135860 295014 135916
rect 295070 135860 295138 135916
rect 295194 135860 295228 135916
rect 293988 135826 295228 135860
rect 313988 136412 315228 136446
rect 313988 136356 314022 136412
rect 314078 136356 314146 136412
rect 314202 136356 314270 136412
rect 314326 136356 314394 136412
rect 314450 136356 314518 136412
rect 314574 136356 314642 136412
rect 314698 136356 314766 136412
rect 314822 136356 314890 136412
rect 314946 136356 315014 136412
rect 315070 136356 315138 136412
rect 315194 136356 315228 136412
rect 313988 136288 315228 136356
rect 313988 136232 314022 136288
rect 314078 136232 314146 136288
rect 314202 136232 314270 136288
rect 314326 136232 314394 136288
rect 314450 136232 314518 136288
rect 314574 136232 314642 136288
rect 314698 136232 314766 136288
rect 314822 136232 314890 136288
rect 314946 136232 315014 136288
rect 315070 136232 315138 136288
rect 315194 136232 315228 136288
rect 313988 136164 315228 136232
rect 313988 136108 314022 136164
rect 314078 136108 314146 136164
rect 314202 136108 314270 136164
rect 314326 136108 314394 136164
rect 314450 136108 314518 136164
rect 314574 136108 314642 136164
rect 314698 136108 314766 136164
rect 314822 136108 314890 136164
rect 314946 136108 315014 136164
rect 315070 136108 315138 136164
rect 315194 136108 315228 136164
rect 313988 136040 315228 136108
rect 313988 135984 314022 136040
rect 314078 135984 314146 136040
rect 314202 135984 314270 136040
rect 314326 135984 314394 136040
rect 314450 135984 314518 136040
rect 314574 135984 314642 136040
rect 314698 135984 314766 136040
rect 314822 135984 314890 136040
rect 314946 135984 315014 136040
rect 315070 135984 315138 136040
rect 315194 135984 315228 136040
rect 313988 135916 315228 135984
rect 313988 135860 314022 135916
rect 314078 135860 314146 135916
rect 314202 135860 314270 135916
rect 314326 135860 314394 135916
rect 314450 135860 314518 135916
rect 314574 135860 314642 135916
rect 314698 135860 314766 135916
rect 314822 135860 314890 135916
rect 314946 135860 315014 135916
rect 315070 135860 315138 135916
rect 315194 135860 315228 135916
rect 313988 135826 315228 135860
rect 283988 130412 285228 130446
rect 283988 130356 284022 130412
rect 284078 130356 284146 130412
rect 284202 130356 284270 130412
rect 284326 130356 284394 130412
rect 284450 130356 284518 130412
rect 284574 130356 284642 130412
rect 284698 130356 284766 130412
rect 284822 130356 284890 130412
rect 284946 130356 285014 130412
rect 285070 130356 285138 130412
rect 285194 130356 285228 130412
rect 283988 130288 285228 130356
rect 283988 130232 284022 130288
rect 284078 130232 284146 130288
rect 284202 130232 284270 130288
rect 284326 130232 284394 130288
rect 284450 130232 284518 130288
rect 284574 130232 284642 130288
rect 284698 130232 284766 130288
rect 284822 130232 284890 130288
rect 284946 130232 285014 130288
rect 285070 130232 285138 130288
rect 285194 130232 285228 130288
rect 283988 130164 285228 130232
rect 283988 130108 284022 130164
rect 284078 130108 284146 130164
rect 284202 130108 284270 130164
rect 284326 130108 284394 130164
rect 284450 130108 284518 130164
rect 284574 130108 284642 130164
rect 284698 130108 284766 130164
rect 284822 130108 284890 130164
rect 284946 130108 285014 130164
rect 285070 130108 285138 130164
rect 285194 130108 285228 130164
rect 283988 130040 285228 130108
rect 283988 129984 284022 130040
rect 284078 129984 284146 130040
rect 284202 129984 284270 130040
rect 284326 129984 284394 130040
rect 284450 129984 284518 130040
rect 284574 129984 284642 130040
rect 284698 129984 284766 130040
rect 284822 129984 284890 130040
rect 284946 129984 285014 130040
rect 285070 129984 285138 130040
rect 285194 129984 285228 130040
rect 283988 129916 285228 129984
rect 283988 129860 284022 129916
rect 284078 129860 284146 129916
rect 284202 129860 284270 129916
rect 284326 129860 284394 129916
rect 284450 129860 284518 129916
rect 284574 129860 284642 129916
rect 284698 129860 284766 129916
rect 284822 129860 284890 129916
rect 284946 129860 285014 129916
rect 285070 129860 285138 129916
rect 285194 129860 285228 129916
rect 283988 129826 285228 129860
rect 303988 130412 305228 130446
rect 303988 130356 304022 130412
rect 304078 130356 304146 130412
rect 304202 130356 304270 130412
rect 304326 130356 304394 130412
rect 304450 130356 304518 130412
rect 304574 130356 304642 130412
rect 304698 130356 304766 130412
rect 304822 130356 304890 130412
rect 304946 130356 305014 130412
rect 305070 130356 305138 130412
rect 305194 130356 305228 130412
rect 303988 130288 305228 130356
rect 303988 130232 304022 130288
rect 304078 130232 304146 130288
rect 304202 130232 304270 130288
rect 304326 130232 304394 130288
rect 304450 130232 304518 130288
rect 304574 130232 304642 130288
rect 304698 130232 304766 130288
rect 304822 130232 304890 130288
rect 304946 130232 305014 130288
rect 305070 130232 305138 130288
rect 305194 130232 305228 130288
rect 303988 130164 305228 130232
rect 303988 130108 304022 130164
rect 304078 130108 304146 130164
rect 304202 130108 304270 130164
rect 304326 130108 304394 130164
rect 304450 130108 304518 130164
rect 304574 130108 304642 130164
rect 304698 130108 304766 130164
rect 304822 130108 304890 130164
rect 304946 130108 305014 130164
rect 305070 130108 305138 130164
rect 305194 130108 305228 130164
rect 303988 130040 305228 130108
rect 303988 129984 304022 130040
rect 304078 129984 304146 130040
rect 304202 129984 304270 130040
rect 304326 129984 304394 130040
rect 304450 129984 304518 130040
rect 304574 129984 304642 130040
rect 304698 129984 304766 130040
rect 304822 129984 304890 130040
rect 304946 129984 305014 130040
rect 305070 129984 305138 130040
rect 305194 129984 305228 130040
rect 303988 129916 305228 129984
rect 303988 129860 304022 129916
rect 304078 129860 304146 129916
rect 304202 129860 304270 129916
rect 304326 129860 304394 129916
rect 304450 129860 304518 129916
rect 304574 129860 304642 129916
rect 304698 129860 304766 129916
rect 304822 129860 304890 129916
rect 304946 129860 305014 129916
rect 305070 129860 305138 129916
rect 305194 129860 305228 129916
rect 303988 129826 305228 129860
rect 327154 130350 327774 147922
rect 327154 130294 327250 130350
rect 327306 130294 327374 130350
rect 327430 130294 327498 130350
rect 327554 130294 327622 130350
rect 327678 130294 327774 130350
rect 327154 130226 327774 130294
rect 327154 130170 327250 130226
rect 327306 130170 327374 130226
rect 327430 130170 327498 130226
rect 327554 130170 327622 130226
rect 327678 130170 327774 130226
rect 327154 130102 327774 130170
rect 327154 130046 327250 130102
rect 327306 130046 327374 130102
rect 327430 130046 327498 130102
rect 327554 130046 327622 130102
rect 327678 130046 327774 130102
rect 327154 129978 327774 130046
rect 327154 129922 327250 129978
rect 327306 129922 327374 129978
rect 327430 129922 327498 129978
rect 327554 129922 327622 129978
rect 327678 129922 327774 129978
rect 276874 118294 276970 118350
rect 277026 118294 277094 118350
rect 277150 118294 277218 118350
rect 277274 118294 277342 118350
rect 277398 118294 277494 118350
rect 276874 118226 277494 118294
rect 276874 118170 276970 118226
rect 277026 118170 277094 118226
rect 277150 118170 277218 118226
rect 277274 118170 277342 118226
rect 277398 118170 277494 118226
rect 276874 118102 277494 118170
rect 276874 118046 276970 118102
rect 277026 118046 277094 118102
rect 277150 118046 277218 118102
rect 277274 118046 277342 118102
rect 277398 118046 277494 118102
rect 276874 117978 277494 118046
rect 276874 117922 276970 117978
rect 277026 117922 277094 117978
rect 277150 117922 277218 117978
rect 277274 117922 277342 117978
rect 277398 117922 277494 117978
rect 273154 112294 273250 112350
rect 273306 112294 273374 112350
rect 273430 112294 273498 112350
rect 273554 112294 273622 112350
rect 273678 112294 273774 112350
rect 273154 112226 273774 112294
rect 273154 112170 273250 112226
rect 273306 112170 273374 112226
rect 273430 112170 273498 112226
rect 273554 112170 273622 112226
rect 273678 112170 273774 112226
rect 273154 112102 273774 112170
rect 273154 112046 273250 112102
rect 273306 112046 273374 112102
rect 273430 112046 273498 112102
rect 273554 112046 273622 112102
rect 273678 112046 273774 112102
rect 273154 111978 273774 112046
rect 273154 111922 273250 111978
rect 273306 111922 273374 111978
rect 273430 111922 273498 111978
rect 273554 111922 273622 111978
rect 273678 111922 273774 111978
rect 273154 94350 273774 111922
rect 275548 113428 275604 113438
rect 275548 111524 275604 113372
rect 275548 111458 275604 111468
rect 273868 101780 273924 101790
rect 273868 99204 273924 101724
rect 275548 101668 275604 101678
rect 275548 100324 275604 101612
rect 275548 100258 275604 100268
rect 276874 100350 277494 117922
rect 293988 118412 295228 118446
rect 293988 118356 294022 118412
rect 294078 118356 294146 118412
rect 294202 118356 294270 118412
rect 294326 118356 294394 118412
rect 294450 118356 294518 118412
rect 294574 118356 294642 118412
rect 294698 118356 294766 118412
rect 294822 118356 294890 118412
rect 294946 118356 295014 118412
rect 295070 118356 295138 118412
rect 295194 118356 295228 118412
rect 293988 118288 295228 118356
rect 293988 118232 294022 118288
rect 294078 118232 294146 118288
rect 294202 118232 294270 118288
rect 294326 118232 294394 118288
rect 294450 118232 294518 118288
rect 294574 118232 294642 118288
rect 294698 118232 294766 118288
rect 294822 118232 294890 118288
rect 294946 118232 295014 118288
rect 295070 118232 295138 118288
rect 295194 118232 295228 118288
rect 293988 118164 295228 118232
rect 293988 118108 294022 118164
rect 294078 118108 294146 118164
rect 294202 118108 294270 118164
rect 294326 118108 294394 118164
rect 294450 118108 294518 118164
rect 294574 118108 294642 118164
rect 294698 118108 294766 118164
rect 294822 118108 294890 118164
rect 294946 118108 295014 118164
rect 295070 118108 295138 118164
rect 295194 118108 295228 118164
rect 293988 118040 295228 118108
rect 293988 117984 294022 118040
rect 294078 117984 294146 118040
rect 294202 117984 294270 118040
rect 294326 117984 294394 118040
rect 294450 117984 294518 118040
rect 294574 117984 294642 118040
rect 294698 117984 294766 118040
rect 294822 117984 294890 118040
rect 294946 117984 295014 118040
rect 295070 117984 295138 118040
rect 295194 117984 295228 118040
rect 293988 117916 295228 117984
rect 293988 117860 294022 117916
rect 294078 117860 294146 117916
rect 294202 117860 294270 117916
rect 294326 117860 294394 117916
rect 294450 117860 294518 117916
rect 294574 117860 294642 117916
rect 294698 117860 294766 117916
rect 294822 117860 294890 117916
rect 294946 117860 295014 117916
rect 295070 117860 295138 117916
rect 295194 117860 295228 117916
rect 293988 117826 295228 117860
rect 313988 118412 315228 118446
rect 313988 118356 314022 118412
rect 314078 118356 314146 118412
rect 314202 118356 314270 118412
rect 314326 118356 314394 118412
rect 314450 118356 314518 118412
rect 314574 118356 314642 118412
rect 314698 118356 314766 118412
rect 314822 118356 314890 118412
rect 314946 118356 315014 118412
rect 315070 118356 315138 118412
rect 315194 118356 315228 118412
rect 313988 118288 315228 118356
rect 313988 118232 314022 118288
rect 314078 118232 314146 118288
rect 314202 118232 314270 118288
rect 314326 118232 314394 118288
rect 314450 118232 314518 118288
rect 314574 118232 314642 118288
rect 314698 118232 314766 118288
rect 314822 118232 314890 118288
rect 314946 118232 315014 118288
rect 315070 118232 315138 118288
rect 315194 118232 315228 118288
rect 313988 118164 315228 118232
rect 313988 118108 314022 118164
rect 314078 118108 314146 118164
rect 314202 118108 314270 118164
rect 314326 118108 314394 118164
rect 314450 118108 314518 118164
rect 314574 118108 314642 118164
rect 314698 118108 314766 118164
rect 314822 118108 314890 118164
rect 314946 118108 315014 118164
rect 315070 118108 315138 118164
rect 315194 118108 315228 118164
rect 313988 118040 315228 118108
rect 313988 117984 314022 118040
rect 314078 117984 314146 118040
rect 314202 117984 314270 118040
rect 314326 117984 314394 118040
rect 314450 117984 314518 118040
rect 314574 117984 314642 118040
rect 314698 117984 314766 118040
rect 314822 117984 314890 118040
rect 314946 117984 315014 118040
rect 315070 117984 315138 118040
rect 315194 117984 315228 118040
rect 313988 117916 315228 117984
rect 313988 117860 314022 117916
rect 314078 117860 314146 117916
rect 314202 117860 314270 117916
rect 314326 117860 314394 117916
rect 314450 117860 314518 117916
rect 314574 117860 314642 117916
rect 314698 117860 314766 117916
rect 314822 117860 314890 117916
rect 314946 117860 315014 117916
rect 315070 117860 315138 117916
rect 315194 117860 315228 117916
rect 313988 117826 315228 117860
rect 283988 112412 285228 112446
rect 283988 112356 284022 112412
rect 284078 112356 284146 112412
rect 284202 112356 284270 112412
rect 284326 112356 284394 112412
rect 284450 112356 284518 112412
rect 284574 112356 284642 112412
rect 284698 112356 284766 112412
rect 284822 112356 284890 112412
rect 284946 112356 285014 112412
rect 285070 112356 285138 112412
rect 285194 112356 285228 112412
rect 283988 112288 285228 112356
rect 283988 112232 284022 112288
rect 284078 112232 284146 112288
rect 284202 112232 284270 112288
rect 284326 112232 284394 112288
rect 284450 112232 284518 112288
rect 284574 112232 284642 112288
rect 284698 112232 284766 112288
rect 284822 112232 284890 112288
rect 284946 112232 285014 112288
rect 285070 112232 285138 112288
rect 285194 112232 285228 112288
rect 283988 112164 285228 112232
rect 283988 112108 284022 112164
rect 284078 112108 284146 112164
rect 284202 112108 284270 112164
rect 284326 112108 284394 112164
rect 284450 112108 284518 112164
rect 284574 112108 284642 112164
rect 284698 112108 284766 112164
rect 284822 112108 284890 112164
rect 284946 112108 285014 112164
rect 285070 112108 285138 112164
rect 285194 112108 285228 112164
rect 283988 112040 285228 112108
rect 283988 111984 284022 112040
rect 284078 111984 284146 112040
rect 284202 111984 284270 112040
rect 284326 111984 284394 112040
rect 284450 111984 284518 112040
rect 284574 111984 284642 112040
rect 284698 111984 284766 112040
rect 284822 111984 284890 112040
rect 284946 111984 285014 112040
rect 285070 111984 285138 112040
rect 285194 111984 285228 112040
rect 283988 111916 285228 111984
rect 283988 111860 284022 111916
rect 284078 111860 284146 111916
rect 284202 111860 284270 111916
rect 284326 111860 284394 111916
rect 284450 111860 284518 111916
rect 284574 111860 284642 111916
rect 284698 111860 284766 111916
rect 284822 111860 284890 111916
rect 284946 111860 285014 111916
rect 285070 111860 285138 111916
rect 285194 111860 285228 111916
rect 283988 111826 285228 111860
rect 303988 112412 305228 112446
rect 303988 112356 304022 112412
rect 304078 112356 304146 112412
rect 304202 112356 304270 112412
rect 304326 112356 304394 112412
rect 304450 112356 304518 112412
rect 304574 112356 304642 112412
rect 304698 112356 304766 112412
rect 304822 112356 304890 112412
rect 304946 112356 305014 112412
rect 305070 112356 305138 112412
rect 305194 112356 305228 112412
rect 303988 112288 305228 112356
rect 303988 112232 304022 112288
rect 304078 112232 304146 112288
rect 304202 112232 304270 112288
rect 304326 112232 304394 112288
rect 304450 112232 304518 112288
rect 304574 112232 304642 112288
rect 304698 112232 304766 112288
rect 304822 112232 304890 112288
rect 304946 112232 305014 112288
rect 305070 112232 305138 112288
rect 305194 112232 305228 112288
rect 303988 112164 305228 112232
rect 303988 112108 304022 112164
rect 304078 112108 304146 112164
rect 304202 112108 304270 112164
rect 304326 112108 304394 112164
rect 304450 112108 304518 112164
rect 304574 112108 304642 112164
rect 304698 112108 304766 112164
rect 304822 112108 304890 112164
rect 304946 112108 305014 112164
rect 305070 112108 305138 112164
rect 305194 112108 305228 112164
rect 303988 112040 305228 112108
rect 303988 111984 304022 112040
rect 304078 111984 304146 112040
rect 304202 111984 304270 112040
rect 304326 111984 304394 112040
rect 304450 111984 304518 112040
rect 304574 111984 304642 112040
rect 304698 111984 304766 112040
rect 304822 111984 304890 112040
rect 304946 111984 305014 112040
rect 305070 111984 305138 112040
rect 305194 111984 305228 112040
rect 303988 111916 305228 111984
rect 303988 111860 304022 111916
rect 304078 111860 304146 111916
rect 304202 111860 304270 111916
rect 304326 111860 304394 111916
rect 304450 111860 304518 111916
rect 304574 111860 304642 111916
rect 304698 111860 304766 111916
rect 304822 111860 304890 111916
rect 304946 111860 305014 111916
rect 305070 111860 305138 111916
rect 305194 111860 305228 111916
rect 303988 111826 305228 111860
rect 327154 112350 327774 129922
rect 327154 112294 327250 112350
rect 327306 112294 327374 112350
rect 327430 112294 327498 112350
rect 327554 112294 327622 112350
rect 327678 112294 327774 112350
rect 327154 112226 327774 112294
rect 327154 112170 327250 112226
rect 327306 112170 327374 112226
rect 327430 112170 327498 112226
rect 327554 112170 327622 112226
rect 327678 112170 327774 112226
rect 327154 112102 327774 112170
rect 327154 112046 327250 112102
rect 327306 112046 327374 112102
rect 327430 112046 327498 112102
rect 327554 112046 327622 112102
rect 327678 112046 327774 112102
rect 327154 111978 327774 112046
rect 327154 111922 327250 111978
rect 327306 111922 327374 111978
rect 327430 111922 327498 111978
rect 327554 111922 327622 111978
rect 327678 111922 327774 111978
rect 276874 100294 276970 100350
rect 277026 100294 277094 100350
rect 277150 100294 277218 100350
rect 277274 100294 277342 100350
rect 277398 100294 277494 100350
rect 273868 99138 273924 99148
rect 276874 100226 277494 100294
rect 276874 100170 276970 100226
rect 277026 100170 277094 100226
rect 277150 100170 277218 100226
rect 277274 100170 277342 100226
rect 277398 100170 277494 100226
rect 276874 100102 277494 100170
rect 276874 100046 276970 100102
rect 277026 100046 277094 100102
rect 277150 100046 277218 100102
rect 277274 100046 277342 100102
rect 277398 100046 277494 100102
rect 276874 99978 277494 100046
rect 276874 99922 276970 99978
rect 277026 99922 277094 99978
rect 277150 99922 277218 99978
rect 277274 99922 277342 99978
rect 277398 99922 277494 99978
rect 273154 94294 273250 94350
rect 273306 94294 273374 94350
rect 273430 94294 273498 94350
rect 273554 94294 273622 94350
rect 273678 94294 273774 94350
rect 273154 94226 273774 94294
rect 273154 94170 273250 94226
rect 273306 94170 273374 94226
rect 273430 94170 273498 94226
rect 273554 94170 273622 94226
rect 273678 94170 273774 94226
rect 273154 94102 273774 94170
rect 273154 94046 273250 94102
rect 273306 94046 273374 94102
rect 273430 94046 273498 94102
rect 273554 94046 273622 94102
rect 273678 94046 273774 94102
rect 273154 93978 273774 94046
rect 273154 93922 273250 93978
rect 273306 93922 273374 93978
rect 273430 93922 273498 93978
rect 273554 93922 273622 93978
rect 273678 93922 273774 93978
rect 273154 76350 273774 93922
rect 273154 76294 273250 76350
rect 273306 76294 273374 76350
rect 273430 76294 273498 76350
rect 273554 76294 273622 76350
rect 273678 76294 273774 76350
rect 273154 76226 273774 76294
rect 273154 76170 273250 76226
rect 273306 76170 273374 76226
rect 273430 76170 273498 76226
rect 273554 76170 273622 76226
rect 273678 76170 273774 76226
rect 273154 76102 273774 76170
rect 273154 76046 273250 76102
rect 273306 76046 273374 76102
rect 273430 76046 273498 76102
rect 273554 76046 273622 76102
rect 273678 76046 273774 76102
rect 273154 75978 273774 76046
rect 273154 75922 273250 75978
rect 273306 75922 273374 75978
rect 273430 75922 273498 75978
rect 273554 75922 273622 75978
rect 273678 75922 273774 75978
rect 273154 58350 273774 75922
rect 274764 83524 274820 83534
rect 274652 75684 274708 75694
rect 274652 59444 274708 75628
rect 274764 73556 274820 83468
rect 276874 82350 277494 99922
rect 293988 100412 295228 100446
rect 293988 100356 294022 100412
rect 294078 100356 294146 100412
rect 294202 100356 294270 100412
rect 294326 100356 294394 100412
rect 294450 100356 294518 100412
rect 294574 100356 294642 100412
rect 294698 100356 294766 100412
rect 294822 100356 294890 100412
rect 294946 100356 295014 100412
rect 295070 100356 295138 100412
rect 295194 100356 295228 100412
rect 293988 100288 295228 100356
rect 293988 100232 294022 100288
rect 294078 100232 294146 100288
rect 294202 100232 294270 100288
rect 294326 100232 294394 100288
rect 294450 100232 294518 100288
rect 294574 100232 294642 100288
rect 294698 100232 294766 100288
rect 294822 100232 294890 100288
rect 294946 100232 295014 100288
rect 295070 100232 295138 100288
rect 295194 100232 295228 100288
rect 293988 100164 295228 100232
rect 293988 100108 294022 100164
rect 294078 100108 294146 100164
rect 294202 100108 294270 100164
rect 294326 100108 294394 100164
rect 294450 100108 294518 100164
rect 294574 100108 294642 100164
rect 294698 100108 294766 100164
rect 294822 100108 294890 100164
rect 294946 100108 295014 100164
rect 295070 100108 295138 100164
rect 295194 100108 295228 100164
rect 293988 100040 295228 100108
rect 293988 99984 294022 100040
rect 294078 99984 294146 100040
rect 294202 99984 294270 100040
rect 294326 99984 294394 100040
rect 294450 99984 294518 100040
rect 294574 99984 294642 100040
rect 294698 99984 294766 100040
rect 294822 99984 294890 100040
rect 294946 99984 295014 100040
rect 295070 99984 295138 100040
rect 295194 99984 295228 100040
rect 293988 99916 295228 99984
rect 293988 99860 294022 99916
rect 294078 99860 294146 99916
rect 294202 99860 294270 99916
rect 294326 99860 294394 99916
rect 294450 99860 294518 99916
rect 294574 99860 294642 99916
rect 294698 99860 294766 99916
rect 294822 99860 294890 99916
rect 294946 99860 295014 99916
rect 295070 99860 295138 99916
rect 295194 99860 295228 99916
rect 293988 99826 295228 99860
rect 313988 100412 315228 100446
rect 313988 100356 314022 100412
rect 314078 100356 314146 100412
rect 314202 100356 314270 100412
rect 314326 100356 314394 100412
rect 314450 100356 314518 100412
rect 314574 100356 314642 100412
rect 314698 100356 314766 100412
rect 314822 100356 314890 100412
rect 314946 100356 315014 100412
rect 315070 100356 315138 100412
rect 315194 100356 315228 100412
rect 313988 100288 315228 100356
rect 313988 100232 314022 100288
rect 314078 100232 314146 100288
rect 314202 100232 314270 100288
rect 314326 100232 314394 100288
rect 314450 100232 314518 100288
rect 314574 100232 314642 100288
rect 314698 100232 314766 100288
rect 314822 100232 314890 100288
rect 314946 100232 315014 100288
rect 315070 100232 315138 100288
rect 315194 100232 315228 100288
rect 313988 100164 315228 100232
rect 313988 100108 314022 100164
rect 314078 100108 314146 100164
rect 314202 100108 314270 100164
rect 314326 100108 314394 100164
rect 314450 100108 314518 100164
rect 314574 100108 314642 100164
rect 314698 100108 314766 100164
rect 314822 100108 314890 100164
rect 314946 100108 315014 100164
rect 315070 100108 315138 100164
rect 315194 100108 315228 100164
rect 313988 100040 315228 100108
rect 313988 99984 314022 100040
rect 314078 99984 314146 100040
rect 314202 99984 314270 100040
rect 314326 99984 314394 100040
rect 314450 99984 314518 100040
rect 314574 99984 314642 100040
rect 314698 99984 314766 100040
rect 314822 99984 314890 100040
rect 314946 99984 315014 100040
rect 315070 99984 315138 100040
rect 315194 99984 315228 100040
rect 313988 99916 315228 99984
rect 313988 99860 314022 99916
rect 314078 99860 314146 99916
rect 314202 99860 314270 99916
rect 314326 99860 314394 99916
rect 314450 99860 314518 99916
rect 314574 99860 314642 99916
rect 314698 99860 314766 99916
rect 314822 99860 314890 99916
rect 314946 99860 315014 99916
rect 315070 99860 315138 99916
rect 315194 99860 315228 99916
rect 313988 99826 315228 99860
rect 283988 94412 285228 94446
rect 283988 94356 284022 94412
rect 284078 94356 284146 94412
rect 284202 94356 284270 94412
rect 284326 94356 284394 94412
rect 284450 94356 284518 94412
rect 284574 94356 284642 94412
rect 284698 94356 284766 94412
rect 284822 94356 284890 94412
rect 284946 94356 285014 94412
rect 285070 94356 285138 94412
rect 285194 94356 285228 94412
rect 283988 94288 285228 94356
rect 283988 94232 284022 94288
rect 284078 94232 284146 94288
rect 284202 94232 284270 94288
rect 284326 94232 284394 94288
rect 284450 94232 284518 94288
rect 284574 94232 284642 94288
rect 284698 94232 284766 94288
rect 284822 94232 284890 94288
rect 284946 94232 285014 94288
rect 285070 94232 285138 94288
rect 285194 94232 285228 94288
rect 283988 94164 285228 94232
rect 283988 94108 284022 94164
rect 284078 94108 284146 94164
rect 284202 94108 284270 94164
rect 284326 94108 284394 94164
rect 284450 94108 284518 94164
rect 284574 94108 284642 94164
rect 284698 94108 284766 94164
rect 284822 94108 284890 94164
rect 284946 94108 285014 94164
rect 285070 94108 285138 94164
rect 285194 94108 285228 94164
rect 283988 94040 285228 94108
rect 283988 93984 284022 94040
rect 284078 93984 284146 94040
rect 284202 93984 284270 94040
rect 284326 93984 284394 94040
rect 284450 93984 284518 94040
rect 284574 93984 284642 94040
rect 284698 93984 284766 94040
rect 284822 93984 284890 94040
rect 284946 93984 285014 94040
rect 285070 93984 285138 94040
rect 285194 93984 285228 94040
rect 283988 93916 285228 93984
rect 283988 93860 284022 93916
rect 284078 93860 284146 93916
rect 284202 93860 284270 93916
rect 284326 93860 284394 93916
rect 284450 93860 284518 93916
rect 284574 93860 284642 93916
rect 284698 93860 284766 93916
rect 284822 93860 284890 93916
rect 284946 93860 285014 93916
rect 285070 93860 285138 93916
rect 285194 93860 285228 93916
rect 283988 93826 285228 93860
rect 303988 94412 305228 94446
rect 303988 94356 304022 94412
rect 304078 94356 304146 94412
rect 304202 94356 304270 94412
rect 304326 94356 304394 94412
rect 304450 94356 304518 94412
rect 304574 94356 304642 94412
rect 304698 94356 304766 94412
rect 304822 94356 304890 94412
rect 304946 94356 305014 94412
rect 305070 94356 305138 94412
rect 305194 94356 305228 94412
rect 303988 94288 305228 94356
rect 303988 94232 304022 94288
rect 304078 94232 304146 94288
rect 304202 94232 304270 94288
rect 304326 94232 304394 94288
rect 304450 94232 304518 94288
rect 304574 94232 304642 94288
rect 304698 94232 304766 94288
rect 304822 94232 304890 94288
rect 304946 94232 305014 94288
rect 305070 94232 305138 94288
rect 305194 94232 305228 94288
rect 303988 94164 305228 94232
rect 303988 94108 304022 94164
rect 304078 94108 304146 94164
rect 304202 94108 304270 94164
rect 304326 94108 304394 94164
rect 304450 94108 304518 94164
rect 304574 94108 304642 94164
rect 304698 94108 304766 94164
rect 304822 94108 304890 94164
rect 304946 94108 305014 94164
rect 305070 94108 305138 94164
rect 305194 94108 305228 94164
rect 303988 94040 305228 94108
rect 303988 93984 304022 94040
rect 304078 93984 304146 94040
rect 304202 93984 304270 94040
rect 304326 93984 304394 94040
rect 304450 93984 304518 94040
rect 304574 93984 304642 94040
rect 304698 93984 304766 94040
rect 304822 93984 304890 94040
rect 304946 93984 305014 94040
rect 305070 93984 305138 94040
rect 305194 93984 305228 94040
rect 303988 93916 305228 93984
rect 303988 93860 304022 93916
rect 304078 93860 304146 93916
rect 304202 93860 304270 93916
rect 304326 93860 304394 93916
rect 304450 93860 304518 93916
rect 304574 93860 304642 93916
rect 304698 93860 304766 93916
rect 304822 93860 304890 93916
rect 304946 93860 305014 93916
rect 305070 93860 305138 93916
rect 305194 93860 305228 93916
rect 303988 93826 305228 93860
rect 327154 94350 327774 111922
rect 327154 94294 327250 94350
rect 327306 94294 327374 94350
rect 327430 94294 327498 94350
rect 327554 94294 327622 94350
rect 327678 94294 327774 94350
rect 327154 94226 327774 94294
rect 327154 94170 327250 94226
rect 327306 94170 327374 94226
rect 327430 94170 327498 94226
rect 327554 94170 327622 94226
rect 327678 94170 327774 94226
rect 327154 94102 327774 94170
rect 327154 94046 327250 94102
rect 327306 94046 327374 94102
rect 327430 94046 327498 94102
rect 327554 94046 327622 94102
rect 327678 94046 327774 94102
rect 327154 93978 327774 94046
rect 327154 93922 327250 93978
rect 327306 93922 327374 93978
rect 327430 93922 327498 93978
rect 327554 93922 327622 93978
rect 327678 93922 327774 93978
rect 276874 82294 276970 82350
rect 277026 82294 277094 82350
rect 277150 82294 277218 82350
rect 277274 82294 277342 82350
rect 277398 82294 277494 82350
rect 276874 82226 277494 82294
rect 276874 82170 276970 82226
rect 277026 82170 277094 82226
rect 277150 82170 277218 82226
rect 277274 82170 277342 82226
rect 277398 82170 277494 82226
rect 276874 82102 277494 82170
rect 276874 82046 276970 82102
rect 277026 82046 277094 82102
rect 277150 82046 277218 82102
rect 277274 82046 277342 82102
rect 277398 82046 277494 82102
rect 276874 81978 277494 82046
rect 276874 81922 276970 81978
rect 277026 81922 277094 81978
rect 277150 81922 277218 81978
rect 277274 81922 277342 81978
rect 277398 81922 277494 81978
rect 274764 73490 274820 73500
rect 275548 76804 275604 76814
rect 275548 73108 275604 76748
rect 275548 73042 275604 73052
rect 274652 59378 274708 59388
rect 276874 64350 277494 81922
rect 293988 82412 295228 82446
rect 293988 82356 294022 82412
rect 294078 82356 294146 82412
rect 294202 82356 294270 82412
rect 294326 82356 294394 82412
rect 294450 82356 294518 82412
rect 294574 82356 294642 82412
rect 294698 82356 294766 82412
rect 294822 82356 294890 82412
rect 294946 82356 295014 82412
rect 295070 82356 295138 82412
rect 295194 82356 295228 82412
rect 293988 82288 295228 82356
rect 293988 82232 294022 82288
rect 294078 82232 294146 82288
rect 294202 82232 294270 82288
rect 294326 82232 294394 82288
rect 294450 82232 294518 82288
rect 294574 82232 294642 82288
rect 294698 82232 294766 82288
rect 294822 82232 294890 82288
rect 294946 82232 295014 82288
rect 295070 82232 295138 82288
rect 295194 82232 295228 82288
rect 293988 82164 295228 82232
rect 293988 82108 294022 82164
rect 294078 82108 294146 82164
rect 294202 82108 294270 82164
rect 294326 82108 294394 82164
rect 294450 82108 294518 82164
rect 294574 82108 294642 82164
rect 294698 82108 294766 82164
rect 294822 82108 294890 82164
rect 294946 82108 295014 82164
rect 295070 82108 295138 82164
rect 295194 82108 295228 82164
rect 293988 82040 295228 82108
rect 293988 81984 294022 82040
rect 294078 81984 294146 82040
rect 294202 81984 294270 82040
rect 294326 81984 294394 82040
rect 294450 81984 294518 82040
rect 294574 81984 294642 82040
rect 294698 81984 294766 82040
rect 294822 81984 294890 82040
rect 294946 81984 295014 82040
rect 295070 81984 295138 82040
rect 295194 81984 295228 82040
rect 293988 81916 295228 81984
rect 293988 81860 294022 81916
rect 294078 81860 294146 81916
rect 294202 81860 294270 81916
rect 294326 81860 294394 81916
rect 294450 81860 294518 81916
rect 294574 81860 294642 81916
rect 294698 81860 294766 81916
rect 294822 81860 294890 81916
rect 294946 81860 295014 81916
rect 295070 81860 295138 81916
rect 295194 81860 295228 81916
rect 293988 81826 295228 81860
rect 313988 82412 315228 82446
rect 313988 82356 314022 82412
rect 314078 82356 314146 82412
rect 314202 82356 314270 82412
rect 314326 82356 314394 82412
rect 314450 82356 314518 82412
rect 314574 82356 314642 82412
rect 314698 82356 314766 82412
rect 314822 82356 314890 82412
rect 314946 82356 315014 82412
rect 315070 82356 315138 82412
rect 315194 82356 315228 82412
rect 313988 82288 315228 82356
rect 313988 82232 314022 82288
rect 314078 82232 314146 82288
rect 314202 82232 314270 82288
rect 314326 82232 314394 82288
rect 314450 82232 314518 82288
rect 314574 82232 314642 82288
rect 314698 82232 314766 82288
rect 314822 82232 314890 82288
rect 314946 82232 315014 82288
rect 315070 82232 315138 82288
rect 315194 82232 315228 82288
rect 313988 82164 315228 82232
rect 313988 82108 314022 82164
rect 314078 82108 314146 82164
rect 314202 82108 314270 82164
rect 314326 82108 314394 82164
rect 314450 82108 314518 82164
rect 314574 82108 314642 82164
rect 314698 82108 314766 82164
rect 314822 82108 314890 82164
rect 314946 82108 315014 82164
rect 315070 82108 315138 82164
rect 315194 82108 315228 82164
rect 313988 82040 315228 82108
rect 313988 81984 314022 82040
rect 314078 81984 314146 82040
rect 314202 81984 314270 82040
rect 314326 81984 314394 82040
rect 314450 81984 314518 82040
rect 314574 81984 314642 82040
rect 314698 81984 314766 82040
rect 314822 81984 314890 82040
rect 314946 81984 315014 82040
rect 315070 81984 315138 82040
rect 315194 81984 315228 82040
rect 313988 81916 315228 81984
rect 313988 81860 314022 81916
rect 314078 81860 314146 81916
rect 314202 81860 314270 81916
rect 314326 81860 314394 81916
rect 314450 81860 314518 81916
rect 314574 81860 314642 81916
rect 314698 81860 314766 81916
rect 314822 81860 314890 81916
rect 314946 81860 315014 81916
rect 315070 81860 315138 81916
rect 315194 81860 315228 81916
rect 313988 81826 315228 81860
rect 283988 76412 285228 76446
rect 283988 76356 284022 76412
rect 284078 76356 284146 76412
rect 284202 76356 284270 76412
rect 284326 76356 284394 76412
rect 284450 76356 284518 76412
rect 284574 76356 284642 76412
rect 284698 76356 284766 76412
rect 284822 76356 284890 76412
rect 284946 76356 285014 76412
rect 285070 76356 285138 76412
rect 285194 76356 285228 76412
rect 283988 76288 285228 76356
rect 283988 76232 284022 76288
rect 284078 76232 284146 76288
rect 284202 76232 284270 76288
rect 284326 76232 284394 76288
rect 284450 76232 284518 76288
rect 284574 76232 284642 76288
rect 284698 76232 284766 76288
rect 284822 76232 284890 76288
rect 284946 76232 285014 76288
rect 285070 76232 285138 76288
rect 285194 76232 285228 76288
rect 283988 76164 285228 76232
rect 283988 76108 284022 76164
rect 284078 76108 284146 76164
rect 284202 76108 284270 76164
rect 284326 76108 284394 76164
rect 284450 76108 284518 76164
rect 284574 76108 284642 76164
rect 284698 76108 284766 76164
rect 284822 76108 284890 76164
rect 284946 76108 285014 76164
rect 285070 76108 285138 76164
rect 285194 76108 285228 76164
rect 283988 76040 285228 76108
rect 283988 75984 284022 76040
rect 284078 75984 284146 76040
rect 284202 75984 284270 76040
rect 284326 75984 284394 76040
rect 284450 75984 284518 76040
rect 284574 75984 284642 76040
rect 284698 75984 284766 76040
rect 284822 75984 284890 76040
rect 284946 75984 285014 76040
rect 285070 75984 285138 76040
rect 285194 75984 285228 76040
rect 283988 75916 285228 75984
rect 283988 75860 284022 75916
rect 284078 75860 284146 75916
rect 284202 75860 284270 75916
rect 284326 75860 284394 75916
rect 284450 75860 284518 75916
rect 284574 75860 284642 75916
rect 284698 75860 284766 75916
rect 284822 75860 284890 75916
rect 284946 75860 285014 75916
rect 285070 75860 285138 75916
rect 285194 75860 285228 75916
rect 283988 75826 285228 75860
rect 291154 76350 291774 79330
rect 291154 76294 291250 76350
rect 291306 76294 291374 76350
rect 291430 76294 291498 76350
rect 291554 76294 291622 76350
rect 291678 76294 291774 76350
rect 291154 76226 291774 76294
rect 291154 76170 291250 76226
rect 291306 76170 291374 76226
rect 291430 76170 291498 76226
rect 291554 76170 291622 76226
rect 291678 76170 291774 76226
rect 291154 76102 291774 76170
rect 291154 76046 291250 76102
rect 291306 76046 291374 76102
rect 291430 76046 291498 76102
rect 291554 76046 291622 76102
rect 291678 76046 291774 76102
rect 291154 75978 291774 76046
rect 291154 75922 291250 75978
rect 291306 75922 291374 75978
rect 291430 75922 291498 75978
rect 291554 75922 291622 75978
rect 291678 75922 291774 75978
rect 276874 64294 276970 64350
rect 277026 64294 277094 64350
rect 277150 64294 277218 64350
rect 277274 64294 277342 64350
rect 277398 64294 277494 64350
rect 276874 64226 277494 64294
rect 276874 64170 276970 64226
rect 277026 64170 277094 64226
rect 277150 64170 277218 64226
rect 277274 64170 277342 64226
rect 277398 64170 277494 64226
rect 276874 64102 277494 64170
rect 276874 64046 276970 64102
rect 277026 64046 277094 64102
rect 277150 64046 277218 64102
rect 277274 64046 277342 64102
rect 277398 64046 277494 64102
rect 276874 63978 277494 64046
rect 276874 63922 276970 63978
rect 277026 63922 277094 63978
rect 277150 63922 277218 63978
rect 277274 63922 277342 63978
rect 277398 63922 277494 63978
rect 273154 58294 273250 58350
rect 273306 58294 273374 58350
rect 273430 58294 273498 58350
rect 273554 58294 273622 58350
rect 273678 58294 273774 58350
rect 273154 58226 273774 58294
rect 273154 58170 273250 58226
rect 273306 58170 273374 58226
rect 273430 58170 273498 58226
rect 273554 58170 273622 58226
rect 273678 58170 273774 58226
rect 273154 58102 273774 58170
rect 273154 58046 273250 58102
rect 273306 58046 273374 58102
rect 273430 58046 273498 58102
rect 273554 58046 273622 58102
rect 273678 58046 273774 58102
rect 273154 57978 273774 58046
rect 273154 57922 273250 57978
rect 273306 57922 273374 57978
rect 273430 57922 273498 57978
rect 273554 57922 273622 57978
rect 273678 57922 273774 57978
rect 273154 40350 273774 57922
rect 273154 40294 273250 40350
rect 273306 40294 273374 40350
rect 273430 40294 273498 40350
rect 273554 40294 273622 40350
rect 273678 40294 273774 40350
rect 273154 40226 273774 40294
rect 273154 40170 273250 40226
rect 273306 40170 273374 40226
rect 273430 40170 273498 40226
rect 273554 40170 273622 40226
rect 273678 40170 273774 40226
rect 273154 40102 273774 40170
rect 273154 40046 273250 40102
rect 273306 40046 273374 40102
rect 273430 40046 273498 40102
rect 273554 40046 273622 40102
rect 273678 40046 273774 40102
rect 273154 39978 273774 40046
rect 273154 39922 273250 39978
rect 273306 39922 273374 39978
rect 273430 39922 273498 39978
rect 273554 39922 273622 39978
rect 273678 39922 273774 39978
rect 273154 22350 273774 39922
rect 273154 22294 273250 22350
rect 273306 22294 273374 22350
rect 273430 22294 273498 22350
rect 273554 22294 273622 22350
rect 273678 22294 273774 22350
rect 273154 22226 273774 22294
rect 273154 22170 273250 22226
rect 273306 22170 273374 22226
rect 273430 22170 273498 22226
rect 273554 22170 273622 22226
rect 273678 22170 273774 22226
rect 273154 22102 273774 22170
rect 273154 22046 273250 22102
rect 273306 22046 273374 22102
rect 273430 22046 273498 22102
rect 273554 22046 273622 22102
rect 273678 22046 273774 22102
rect 273154 21978 273774 22046
rect 273154 21922 273250 21978
rect 273306 21922 273374 21978
rect 273430 21922 273498 21978
rect 273554 21922 273622 21978
rect 273678 21922 273774 21978
rect 273154 4350 273774 21922
rect 273154 4294 273250 4350
rect 273306 4294 273374 4350
rect 273430 4294 273498 4350
rect 273554 4294 273622 4350
rect 273678 4294 273774 4350
rect 273154 4226 273774 4294
rect 273154 4170 273250 4226
rect 273306 4170 273374 4226
rect 273430 4170 273498 4226
rect 273554 4170 273622 4226
rect 273678 4170 273774 4226
rect 273154 4102 273774 4170
rect 273154 4046 273250 4102
rect 273306 4046 273374 4102
rect 273430 4046 273498 4102
rect 273554 4046 273622 4102
rect 273678 4046 273774 4102
rect 273154 3978 273774 4046
rect 273154 3922 273250 3978
rect 273306 3922 273374 3978
rect 273430 3922 273498 3978
rect 273554 3922 273622 3978
rect 273678 3922 273774 3978
rect 273154 -160 273774 3922
rect 273154 -216 273250 -160
rect 273306 -216 273374 -160
rect 273430 -216 273498 -160
rect 273554 -216 273622 -160
rect 273678 -216 273774 -160
rect 273154 -284 273774 -216
rect 273154 -340 273250 -284
rect 273306 -340 273374 -284
rect 273430 -340 273498 -284
rect 273554 -340 273622 -284
rect 273678 -340 273774 -284
rect 273154 -408 273774 -340
rect 273154 -464 273250 -408
rect 273306 -464 273374 -408
rect 273430 -464 273498 -408
rect 273554 -464 273622 -408
rect 273678 -464 273774 -408
rect 273154 -532 273774 -464
rect 273154 -588 273250 -532
rect 273306 -588 273374 -532
rect 273430 -588 273498 -532
rect 273554 -588 273622 -532
rect 273678 -588 273774 -532
rect 273154 -1644 273774 -588
rect 276874 46350 277494 63922
rect 276874 46294 276970 46350
rect 277026 46294 277094 46350
rect 277150 46294 277218 46350
rect 277274 46294 277342 46350
rect 277398 46294 277494 46350
rect 276874 46226 277494 46294
rect 276874 46170 276970 46226
rect 277026 46170 277094 46226
rect 277150 46170 277218 46226
rect 277274 46170 277342 46226
rect 277398 46170 277494 46226
rect 276874 46102 277494 46170
rect 276874 46046 276970 46102
rect 277026 46046 277094 46102
rect 277150 46046 277218 46102
rect 277274 46046 277342 46102
rect 277398 46046 277494 46102
rect 276874 45978 277494 46046
rect 276874 45922 276970 45978
rect 277026 45922 277094 45978
rect 277150 45922 277218 45978
rect 277274 45922 277342 45978
rect 277398 45922 277494 45978
rect 276874 28350 277494 45922
rect 276874 28294 276970 28350
rect 277026 28294 277094 28350
rect 277150 28294 277218 28350
rect 277274 28294 277342 28350
rect 277398 28294 277494 28350
rect 276874 28226 277494 28294
rect 276874 28170 276970 28226
rect 277026 28170 277094 28226
rect 277150 28170 277218 28226
rect 277274 28170 277342 28226
rect 277398 28170 277494 28226
rect 276874 28102 277494 28170
rect 276874 28046 276970 28102
rect 277026 28046 277094 28102
rect 277150 28046 277218 28102
rect 277274 28046 277342 28102
rect 277398 28046 277494 28102
rect 276874 27978 277494 28046
rect 276874 27922 276970 27978
rect 277026 27922 277094 27978
rect 277150 27922 277218 27978
rect 277274 27922 277342 27978
rect 277398 27922 277494 27978
rect 276874 10350 277494 27922
rect 276874 10294 276970 10350
rect 277026 10294 277094 10350
rect 277150 10294 277218 10350
rect 277274 10294 277342 10350
rect 277398 10294 277494 10350
rect 276874 10226 277494 10294
rect 276874 10170 276970 10226
rect 277026 10170 277094 10226
rect 277150 10170 277218 10226
rect 277274 10170 277342 10226
rect 277398 10170 277494 10226
rect 276874 10102 277494 10170
rect 276874 10046 276970 10102
rect 277026 10046 277094 10102
rect 277150 10046 277218 10102
rect 277274 10046 277342 10102
rect 277398 10046 277494 10102
rect 276874 9978 277494 10046
rect 276874 9922 276970 9978
rect 277026 9922 277094 9978
rect 277150 9922 277218 9978
rect 277274 9922 277342 9978
rect 277398 9922 277494 9978
rect 276874 -1120 277494 9922
rect 276874 -1176 276970 -1120
rect 277026 -1176 277094 -1120
rect 277150 -1176 277218 -1120
rect 277274 -1176 277342 -1120
rect 277398 -1176 277494 -1120
rect 276874 -1244 277494 -1176
rect 276874 -1300 276970 -1244
rect 277026 -1300 277094 -1244
rect 277150 -1300 277218 -1244
rect 277274 -1300 277342 -1244
rect 277398 -1300 277494 -1244
rect 276874 -1368 277494 -1300
rect 276874 -1424 276970 -1368
rect 277026 -1424 277094 -1368
rect 277150 -1424 277218 -1368
rect 277274 -1424 277342 -1368
rect 277398 -1424 277494 -1368
rect 276874 -1492 277494 -1424
rect 276874 -1548 276970 -1492
rect 277026 -1548 277094 -1492
rect 277150 -1548 277218 -1492
rect 277274 -1548 277342 -1492
rect 277398 -1548 277494 -1492
rect 276874 -1644 277494 -1548
rect 291154 58350 291774 75922
rect 303988 76412 305228 76446
rect 303988 76356 304022 76412
rect 304078 76356 304146 76412
rect 304202 76356 304270 76412
rect 304326 76356 304394 76412
rect 304450 76356 304518 76412
rect 304574 76356 304642 76412
rect 304698 76356 304766 76412
rect 304822 76356 304890 76412
rect 304946 76356 305014 76412
rect 305070 76356 305138 76412
rect 305194 76356 305228 76412
rect 303988 76288 305228 76356
rect 303988 76232 304022 76288
rect 304078 76232 304146 76288
rect 304202 76232 304270 76288
rect 304326 76232 304394 76288
rect 304450 76232 304518 76288
rect 304574 76232 304642 76288
rect 304698 76232 304766 76288
rect 304822 76232 304890 76288
rect 304946 76232 305014 76288
rect 305070 76232 305138 76288
rect 305194 76232 305228 76288
rect 303988 76164 305228 76232
rect 303988 76108 304022 76164
rect 304078 76108 304146 76164
rect 304202 76108 304270 76164
rect 304326 76108 304394 76164
rect 304450 76108 304518 76164
rect 304574 76108 304642 76164
rect 304698 76108 304766 76164
rect 304822 76108 304890 76164
rect 304946 76108 305014 76164
rect 305070 76108 305138 76164
rect 305194 76108 305228 76164
rect 303988 76040 305228 76108
rect 303988 75984 304022 76040
rect 304078 75984 304146 76040
rect 304202 75984 304270 76040
rect 304326 75984 304394 76040
rect 304450 75984 304518 76040
rect 304574 75984 304642 76040
rect 304698 75984 304766 76040
rect 304822 75984 304890 76040
rect 304946 75984 305014 76040
rect 305070 75984 305138 76040
rect 305194 75984 305228 76040
rect 303988 75916 305228 75984
rect 303988 75860 304022 75916
rect 304078 75860 304146 75916
rect 304202 75860 304270 75916
rect 304326 75860 304394 75916
rect 304450 75860 304518 75916
rect 304574 75860 304642 75916
rect 304698 75860 304766 75916
rect 304822 75860 304890 75916
rect 304946 75860 305014 75916
rect 305070 75860 305138 75916
rect 305194 75860 305228 75916
rect 303988 75826 305228 75860
rect 309154 76350 309774 79330
rect 309154 76294 309250 76350
rect 309306 76294 309374 76350
rect 309430 76294 309498 76350
rect 309554 76294 309622 76350
rect 309678 76294 309774 76350
rect 309154 76226 309774 76294
rect 309154 76170 309250 76226
rect 309306 76170 309374 76226
rect 309430 76170 309498 76226
rect 309554 76170 309622 76226
rect 309678 76170 309774 76226
rect 309154 76102 309774 76170
rect 309154 76046 309250 76102
rect 309306 76046 309374 76102
rect 309430 76046 309498 76102
rect 309554 76046 309622 76102
rect 309678 76046 309774 76102
rect 309154 75978 309774 76046
rect 309154 75922 309250 75978
rect 309306 75922 309374 75978
rect 309430 75922 309498 75978
rect 309554 75922 309622 75978
rect 309678 75922 309774 75978
rect 291154 58294 291250 58350
rect 291306 58294 291374 58350
rect 291430 58294 291498 58350
rect 291554 58294 291622 58350
rect 291678 58294 291774 58350
rect 291154 58226 291774 58294
rect 291154 58170 291250 58226
rect 291306 58170 291374 58226
rect 291430 58170 291498 58226
rect 291554 58170 291622 58226
rect 291678 58170 291774 58226
rect 291154 58102 291774 58170
rect 291154 58046 291250 58102
rect 291306 58046 291374 58102
rect 291430 58046 291498 58102
rect 291554 58046 291622 58102
rect 291678 58046 291774 58102
rect 291154 57978 291774 58046
rect 291154 57922 291250 57978
rect 291306 57922 291374 57978
rect 291430 57922 291498 57978
rect 291554 57922 291622 57978
rect 291678 57922 291774 57978
rect 291154 40350 291774 57922
rect 291154 40294 291250 40350
rect 291306 40294 291374 40350
rect 291430 40294 291498 40350
rect 291554 40294 291622 40350
rect 291678 40294 291774 40350
rect 291154 40226 291774 40294
rect 291154 40170 291250 40226
rect 291306 40170 291374 40226
rect 291430 40170 291498 40226
rect 291554 40170 291622 40226
rect 291678 40170 291774 40226
rect 291154 40102 291774 40170
rect 291154 40046 291250 40102
rect 291306 40046 291374 40102
rect 291430 40046 291498 40102
rect 291554 40046 291622 40102
rect 291678 40046 291774 40102
rect 291154 39978 291774 40046
rect 291154 39922 291250 39978
rect 291306 39922 291374 39978
rect 291430 39922 291498 39978
rect 291554 39922 291622 39978
rect 291678 39922 291774 39978
rect 291154 22350 291774 39922
rect 291154 22294 291250 22350
rect 291306 22294 291374 22350
rect 291430 22294 291498 22350
rect 291554 22294 291622 22350
rect 291678 22294 291774 22350
rect 291154 22226 291774 22294
rect 291154 22170 291250 22226
rect 291306 22170 291374 22226
rect 291430 22170 291498 22226
rect 291554 22170 291622 22226
rect 291678 22170 291774 22226
rect 291154 22102 291774 22170
rect 291154 22046 291250 22102
rect 291306 22046 291374 22102
rect 291430 22046 291498 22102
rect 291554 22046 291622 22102
rect 291678 22046 291774 22102
rect 291154 21978 291774 22046
rect 291154 21922 291250 21978
rect 291306 21922 291374 21978
rect 291430 21922 291498 21978
rect 291554 21922 291622 21978
rect 291678 21922 291774 21978
rect 291154 4350 291774 21922
rect 291154 4294 291250 4350
rect 291306 4294 291374 4350
rect 291430 4294 291498 4350
rect 291554 4294 291622 4350
rect 291678 4294 291774 4350
rect 291154 4226 291774 4294
rect 291154 4170 291250 4226
rect 291306 4170 291374 4226
rect 291430 4170 291498 4226
rect 291554 4170 291622 4226
rect 291678 4170 291774 4226
rect 291154 4102 291774 4170
rect 291154 4046 291250 4102
rect 291306 4046 291374 4102
rect 291430 4046 291498 4102
rect 291554 4046 291622 4102
rect 291678 4046 291774 4102
rect 291154 3978 291774 4046
rect 291154 3922 291250 3978
rect 291306 3922 291374 3978
rect 291430 3922 291498 3978
rect 291554 3922 291622 3978
rect 291678 3922 291774 3978
rect 291154 -160 291774 3922
rect 291154 -216 291250 -160
rect 291306 -216 291374 -160
rect 291430 -216 291498 -160
rect 291554 -216 291622 -160
rect 291678 -216 291774 -160
rect 291154 -284 291774 -216
rect 291154 -340 291250 -284
rect 291306 -340 291374 -284
rect 291430 -340 291498 -284
rect 291554 -340 291622 -284
rect 291678 -340 291774 -284
rect 291154 -408 291774 -340
rect 291154 -464 291250 -408
rect 291306 -464 291374 -408
rect 291430 -464 291498 -408
rect 291554 -464 291622 -408
rect 291678 -464 291774 -408
rect 291154 -532 291774 -464
rect 291154 -588 291250 -532
rect 291306 -588 291374 -532
rect 291430 -588 291498 -532
rect 291554 -588 291622 -532
rect 291678 -588 291774 -532
rect 291154 -1644 291774 -588
rect 294874 64350 295494 70964
rect 294874 64294 294970 64350
rect 295026 64294 295094 64350
rect 295150 64294 295218 64350
rect 295274 64294 295342 64350
rect 295398 64294 295494 64350
rect 294874 64226 295494 64294
rect 294874 64170 294970 64226
rect 295026 64170 295094 64226
rect 295150 64170 295218 64226
rect 295274 64170 295342 64226
rect 295398 64170 295494 64226
rect 294874 64102 295494 64170
rect 294874 64046 294970 64102
rect 295026 64046 295094 64102
rect 295150 64046 295218 64102
rect 295274 64046 295342 64102
rect 295398 64046 295494 64102
rect 294874 63978 295494 64046
rect 294874 63922 294970 63978
rect 295026 63922 295094 63978
rect 295150 63922 295218 63978
rect 295274 63922 295342 63978
rect 295398 63922 295494 63978
rect 294874 46350 295494 63922
rect 294874 46294 294970 46350
rect 295026 46294 295094 46350
rect 295150 46294 295218 46350
rect 295274 46294 295342 46350
rect 295398 46294 295494 46350
rect 294874 46226 295494 46294
rect 294874 46170 294970 46226
rect 295026 46170 295094 46226
rect 295150 46170 295218 46226
rect 295274 46170 295342 46226
rect 295398 46170 295494 46226
rect 294874 46102 295494 46170
rect 294874 46046 294970 46102
rect 295026 46046 295094 46102
rect 295150 46046 295218 46102
rect 295274 46046 295342 46102
rect 295398 46046 295494 46102
rect 294874 45978 295494 46046
rect 294874 45922 294970 45978
rect 295026 45922 295094 45978
rect 295150 45922 295218 45978
rect 295274 45922 295342 45978
rect 295398 45922 295494 45978
rect 294874 28350 295494 45922
rect 294874 28294 294970 28350
rect 295026 28294 295094 28350
rect 295150 28294 295218 28350
rect 295274 28294 295342 28350
rect 295398 28294 295494 28350
rect 294874 28226 295494 28294
rect 294874 28170 294970 28226
rect 295026 28170 295094 28226
rect 295150 28170 295218 28226
rect 295274 28170 295342 28226
rect 295398 28170 295494 28226
rect 294874 28102 295494 28170
rect 294874 28046 294970 28102
rect 295026 28046 295094 28102
rect 295150 28046 295218 28102
rect 295274 28046 295342 28102
rect 295398 28046 295494 28102
rect 294874 27978 295494 28046
rect 294874 27922 294970 27978
rect 295026 27922 295094 27978
rect 295150 27922 295218 27978
rect 295274 27922 295342 27978
rect 295398 27922 295494 27978
rect 294874 10350 295494 27922
rect 294874 10294 294970 10350
rect 295026 10294 295094 10350
rect 295150 10294 295218 10350
rect 295274 10294 295342 10350
rect 295398 10294 295494 10350
rect 294874 10226 295494 10294
rect 294874 10170 294970 10226
rect 295026 10170 295094 10226
rect 295150 10170 295218 10226
rect 295274 10170 295342 10226
rect 295398 10170 295494 10226
rect 294874 10102 295494 10170
rect 294874 10046 294970 10102
rect 295026 10046 295094 10102
rect 295150 10046 295218 10102
rect 295274 10046 295342 10102
rect 295398 10046 295494 10102
rect 294874 9978 295494 10046
rect 294874 9922 294970 9978
rect 295026 9922 295094 9978
rect 295150 9922 295218 9978
rect 295274 9922 295342 9978
rect 295398 9922 295494 9978
rect 294874 -1120 295494 9922
rect 294874 -1176 294970 -1120
rect 295026 -1176 295094 -1120
rect 295150 -1176 295218 -1120
rect 295274 -1176 295342 -1120
rect 295398 -1176 295494 -1120
rect 294874 -1244 295494 -1176
rect 294874 -1300 294970 -1244
rect 295026 -1300 295094 -1244
rect 295150 -1300 295218 -1244
rect 295274 -1300 295342 -1244
rect 295398 -1300 295494 -1244
rect 294874 -1368 295494 -1300
rect 294874 -1424 294970 -1368
rect 295026 -1424 295094 -1368
rect 295150 -1424 295218 -1368
rect 295274 -1424 295342 -1368
rect 295398 -1424 295494 -1368
rect 294874 -1492 295494 -1424
rect 294874 -1548 294970 -1492
rect 295026 -1548 295094 -1492
rect 295150 -1548 295218 -1492
rect 295274 -1548 295342 -1492
rect 295398 -1548 295494 -1492
rect 294874 -1644 295494 -1548
rect 309154 58350 309774 75922
rect 309154 58294 309250 58350
rect 309306 58294 309374 58350
rect 309430 58294 309498 58350
rect 309554 58294 309622 58350
rect 309678 58294 309774 58350
rect 309154 58226 309774 58294
rect 309154 58170 309250 58226
rect 309306 58170 309374 58226
rect 309430 58170 309498 58226
rect 309554 58170 309622 58226
rect 309678 58170 309774 58226
rect 309154 58102 309774 58170
rect 309154 58046 309250 58102
rect 309306 58046 309374 58102
rect 309430 58046 309498 58102
rect 309554 58046 309622 58102
rect 309678 58046 309774 58102
rect 309154 57978 309774 58046
rect 309154 57922 309250 57978
rect 309306 57922 309374 57978
rect 309430 57922 309498 57978
rect 309554 57922 309622 57978
rect 309678 57922 309774 57978
rect 309154 40350 309774 57922
rect 309154 40294 309250 40350
rect 309306 40294 309374 40350
rect 309430 40294 309498 40350
rect 309554 40294 309622 40350
rect 309678 40294 309774 40350
rect 309154 40226 309774 40294
rect 309154 40170 309250 40226
rect 309306 40170 309374 40226
rect 309430 40170 309498 40226
rect 309554 40170 309622 40226
rect 309678 40170 309774 40226
rect 309154 40102 309774 40170
rect 309154 40046 309250 40102
rect 309306 40046 309374 40102
rect 309430 40046 309498 40102
rect 309554 40046 309622 40102
rect 309678 40046 309774 40102
rect 309154 39978 309774 40046
rect 309154 39922 309250 39978
rect 309306 39922 309374 39978
rect 309430 39922 309498 39978
rect 309554 39922 309622 39978
rect 309678 39922 309774 39978
rect 309154 22350 309774 39922
rect 309154 22294 309250 22350
rect 309306 22294 309374 22350
rect 309430 22294 309498 22350
rect 309554 22294 309622 22350
rect 309678 22294 309774 22350
rect 309154 22226 309774 22294
rect 309154 22170 309250 22226
rect 309306 22170 309374 22226
rect 309430 22170 309498 22226
rect 309554 22170 309622 22226
rect 309678 22170 309774 22226
rect 309154 22102 309774 22170
rect 309154 22046 309250 22102
rect 309306 22046 309374 22102
rect 309430 22046 309498 22102
rect 309554 22046 309622 22102
rect 309678 22046 309774 22102
rect 309154 21978 309774 22046
rect 309154 21922 309250 21978
rect 309306 21922 309374 21978
rect 309430 21922 309498 21978
rect 309554 21922 309622 21978
rect 309678 21922 309774 21978
rect 309154 4350 309774 21922
rect 309154 4294 309250 4350
rect 309306 4294 309374 4350
rect 309430 4294 309498 4350
rect 309554 4294 309622 4350
rect 309678 4294 309774 4350
rect 309154 4226 309774 4294
rect 309154 4170 309250 4226
rect 309306 4170 309374 4226
rect 309430 4170 309498 4226
rect 309554 4170 309622 4226
rect 309678 4170 309774 4226
rect 309154 4102 309774 4170
rect 309154 4046 309250 4102
rect 309306 4046 309374 4102
rect 309430 4046 309498 4102
rect 309554 4046 309622 4102
rect 309678 4046 309774 4102
rect 309154 3978 309774 4046
rect 309154 3922 309250 3978
rect 309306 3922 309374 3978
rect 309430 3922 309498 3978
rect 309554 3922 309622 3978
rect 309678 3922 309774 3978
rect 309154 -160 309774 3922
rect 309154 -216 309250 -160
rect 309306 -216 309374 -160
rect 309430 -216 309498 -160
rect 309554 -216 309622 -160
rect 309678 -216 309774 -160
rect 309154 -284 309774 -216
rect 309154 -340 309250 -284
rect 309306 -340 309374 -284
rect 309430 -340 309498 -284
rect 309554 -340 309622 -284
rect 309678 -340 309774 -284
rect 309154 -408 309774 -340
rect 309154 -464 309250 -408
rect 309306 -464 309374 -408
rect 309430 -464 309498 -408
rect 309554 -464 309622 -408
rect 309678 -464 309774 -408
rect 309154 -532 309774 -464
rect 309154 -588 309250 -532
rect 309306 -588 309374 -532
rect 309430 -588 309498 -532
rect 309554 -588 309622 -532
rect 309678 -588 309774 -532
rect 309154 -1644 309774 -588
rect 312874 64350 313494 79330
rect 312874 64294 312970 64350
rect 313026 64294 313094 64350
rect 313150 64294 313218 64350
rect 313274 64294 313342 64350
rect 313398 64294 313494 64350
rect 312874 64226 313494 64294
rect 312874 64170 312970 64226
rect 313026 64170 313094 64226
rect 313150 64170 313218 64226
rect 313274 64170 313342 64226
rect 313398 64170 313494 64226
rect 312874 64102 313494 64170
rect 312874 64046 312970 64102
rect 313026 64046 313094 64102
rect 313150 64046 313218 64102
rect 313274 64046 313342 64102
rect 313398 64046 313494 64102
rect 312874 63978 313494 64046
rect 312874 63922 312970 63978
rect 313026 63922 313094 63978
rect 313150 63922 313218 63978
rect 313274 63922 313342 63978
rect 313398 63922 313494 63978
rect 312874 46350 313494 63922
rect 312874 46294 312970 46350
rect 313026 46294 313094 46350
rect 313150 46294 313218 46350
rect 313274 46294 313342 46350
rect 313398 46294 313494 46350
rect 312874 46226 313494 46294
rect 312874 46170 312970 46226
rect 313026 46170 313094 46226
rect 313150 46170 313218 46226
rect 313274 46170 313342 46226
rect 313398 46170 313494 46226
rect 312874 46102 313494 46170
rect 312874 46046 312970 46102
rect 313026 46046 313094 46102
rect 313150 46046 313218 46102
rect 313274 46046 313342 46102
rect 313398 46046 313494 46102
rect 312874 45978 313494 46046
rect 312874 45922 312970 45978
rect 313026 45922 313094 45978
rect 313150 45922 313218 45978
rect 313274 45922 313342 45978
rect 313398 45922 313494 45978
rect 312874 28350 313494 45922
rect 312874 28294 312970 28350
rect 313026 28294 313094 28350
rect 313150 28294 313218 28350
rect 313274 28294 313342 28350
rect 313398 28294 313494 28350
rect 312874 28226 313494 28294
rect 312874 28170 312970 28226
rect 313026 28170 313094 28226
rect 313150 28170 313218 28226
rect 313274 28170 313342 28226
rect 313398 28170 313494 28226
rect 312874 28102 313494 28170
rect 312874 28046 312970 28102
rect 313026 28046 313094 28102
rect 313150 28046 313218 28102
rect 313274 28046 313342 28102
rect 313398 28046 313494 28102
rect 312874 27978 313494 28046
rect 312874 27922 312970 27978
rect 313026 27922 313094 27978
rect 313150 27922 313218 27978
rect 313274 27922 313342 27978
rect 313398 27922 313494 27978
rect 312874 10350 313494 27922
rect 312874 10294 312970 10350
rect 313026 10294 313094 10350
rect 313150 10294 313218 10350
rect 313274 10294 313342 10350
rect 313398 10294 313494 10350
rect 312874 10226 313494 10294
rect 312874 10170 312970 10226
rect 313026 10170 313094 10226
rect 313150 10170 313218 10226
rect 313274 10170 313342 10226
rect 313398 10170 313494 10226
rect 312874 10102 313494 10170
rect 312874 10046 312970 10102
rect 313026 10046 313094 10102
rect 313150 10046 313218 10102
rect 313274 10046 313342 10102
rect 313398 10046 313494 10102
rect 312874 9978 313494 10046
rect 312874 9922 312970 9978
rect 313026 9922 313094 9978
rect 313150 9922 313218 9978
rect 313274 9922 313342 9978
rect 313398 9922 313494 9978
rect 312874 -1120 313494 9922
rect 312874 -1176 312970 -1120
rect 313026 -1176 313094 -1120
rect 313150 -1176 313218 -1120
rect 313274 -1176 313342 -1120
rect 313398 -1176 313494 -1120
rect 312874 -1244 313494 -1176
rect 312874 -1300 312970 -1244
rect 313026 -1300 313094 -1244
rect 313150 -1300 313218 -1244
rect 313274 -1300 313342 -1244
rect 313398 -1300 313494 -1244
rect 312874 -1368 313494 -1300
rect 312874 -1424 312970 -1368
rect 313026 -1424 313094 -1368
rect 313150 -1424 313218 -1368
rect 313274 -1424 313342 -1368
rect 313398 -1424 313494 -1368
rect 312874 -1492 313494 -1424
rect 312874 -1548 312970 -1492
rect 313026 -1548 313094 -1492
rect 313150 -1548 313218 -1492
rect 313274 -1548 313342 -1492
rect 313398 -1548 313494 -1492
rect 312874 -1644 313494 -1548
rect 327154 76350 327774 93922
rect 327154 76294 327250 76350
rect 327306 76294 327374 76350
rect 327430 76294 327498 76350
rect 327554 76294 327622 76350
rect 327678 76294 327774 76350
rect 327154 76226 327774 76294
rect 327154 76170 327250 76226
rect 327306 76170 327374 76226
rect 327430 76170 327498 76226
rect 327554 76170 327622 76226
rect 327678 76170 327774 76226
rect 327154 76102 327774 76170
rect 327154 76046 327250 76102
rect 327306 76046 327374 76102
rect 327430 76046 327498 76102
rect 327554 76046 327622 76102
rect 327678 76046 327774 76102
rect 327154 75978 327774 76046
rect 327154 75922 327250 75978
rect 327306 75922 327374 75978
rect 327430 75922 327498 75978
rect 327554 75922 327622 75978
rect 327678 75922 327774 75978
rect 327154 58350 327774 75922
rect 327154 58294 327250 58350
rect 327306 58294 327374 58350
rect 327430 58294 327498 58350
rect 327554 58294 327622 58350
rect 327678 58294 327774 58350
rect 327154 58226 327774 58294
rect 327154 58170 327250 58226
rect 327306 58170 327374 58226
rect 327430 58170 327498 58226
rect 327554 58170 327622 58226
rect 327678 58170 327774 58226
rect 327154 58102 327774 58170
rect 327154 58046 327250 58102
rect 327306 58046 327374 58102
rect 327430 58046 327498 58102
rect 327554 58046 327622 58102
rect 327678 58046 327774 58102
rect 327154 57978 327774 58046
rect 327154 57922 327250 57978
rect 327306 57922 327374 57978
rect 327430 57922 327498 57978
rect 327554 57922 327622 57978
rect 327678 57922 327774 57978
rect 327154 40350 327774 57922
rect 327154 40294 327250 40350
rect 327306 40294 327374 40350
rect 327430 40294 327498 40350
rect 327554 40294 327622 40350
rect 327678 40294 327774 40350
rect 327154 40226 327774 40294
rect 327154 40170 327250 40226
rect 327306 40170 327374 40226
rect 327430 40170 327498 40226
rect 327554 40170 327622 40226
rect 327678 40170 327774 40226
rect 327154 40102 327774 40170
rect 327154 40046 327250 40102
rect 327306 40046 327374 40102
rect 327430 40046 327498 40102
rect 327554 40046 327622 40102
rect 327678 40046 327774 40102
rect 327154 39978 327774 40046
rect 327154 39922 327250 39978
rect 327306 39922 327374 39978
rect 327430 39922 327498 39978
rect 327554 39922 327622 39978
rect 327678 39922 327774 39978
rect 327154 22350 327774 39922
rect 327154 22294 327250 22350
rect 327306 22294 327374 22350
rect 327430 22294 327498 22350
rect 327554 22294 327622 22350
rect 327678 22294 327774 22350
rect 327154 22226 327774 22294
rect 327154 22170 327250 22226
rect 327306 22170 327374 22226
rect 327430 22170 327498 22226
rect 327554 22170 327622 22226
rect 327678 22170 327774 22226
rect 327154 22102 327774 22170
rect 327154 22046 327250 22102
rect 327306 22046 327374 22102
rect 327430 22046 327498 22102
rect 327554 22046 327622 22102
rect 327678 22046 327774 22102
rect 327154 21978 327774 22046
rect 327154 21922 327250 21978
rect 327306 21922 327374 21978
rect 327430 21922 327498 21978
rect 327554 21922 327622 21978
rect 327678 21922 327774 21978
rect 327154 4350 327774 21922
rect 327154 4294 327250 4350
rect 327306 4294 327374 4350
rect 327430 4294 327498 4350
rect 327554 4294 327622 4350
rect 327678 4294 327774 4350
rect 327154 4226 327774 4294
rect 327154 4170 327250 4226
rect 327306 4170 327374 4226
rect 327430 4170 327498 4226
rect 327554 4170 327622 4226
rect 327678 4170 327774 4226
rect 327154 4102 327774 4170
rect 327154 4046 327250 4102
rect 327306 4046 327374 4102
rect 327430 4046 327498 4102
rect 327554 4046 327622 4102
rect 327678 4046 327774 4102
rect 327154 3978 327774 4046
rect 327154 3922 327250 3978
rect 327306 3922 327374 3978
rect 327430 3922 327498 3978
rect 327554 3922 327622 3978
rect 327678 3922 327774 3978
rect 327154 -160 327774 3922
rect 327154 -216 327250 -160
rect 327306 -216 327374 -160
rect 327430 -216 327498 -160
rect 327554 -216 327622 -160
rect 327678 -216 327774 -160
rect 327154 -284 327774 -216
rect 327154 -340 327250 -284
rect 327306 -340 327374 -284
rect 327430 -340 327498 -284
rect 327554 -340 327622 -284
rect 327678 -340 327774 -284
rect 327154 -408 327774 -340
rect 327154 -464 327250 -408
rect 327306 -464 327374 -408
rect 327430 -464 327498 -408
rect 327554 -464 327622 -408
rect 327678 -464 327774 -408
rect 327154 -532 327774 -464
rect 327154 -588 327250 -532
rect 327306 -588 327374 -532
rect 327430 -588 327498 -532
rect 327554 -588 327622 -532
rect 327678 -588 327774 -532
rect 327154 -1644 327774 -588
rect 330874 598172 331494 598268
rect 330874 598116 330970 598172
rect 331026 598116 331094 598172
rect 331150 598116 331218 598172
rect 331274 598116 331342 598172
rect 331398 598116 331494 598172
rect 330874 598048 331494 598116
rect 330874 597992 330970 598048
rect 331026 597992 331094 598048
rect 331150 597992 331218 598048
rect 331274 597992 331342 598048
rect 331398 597992 331494 598048
rect 330874 597924 331494 597992
rect 330874 597868 330970 597924
rect 331026 597868 331094 597924
rect 331150 597868 331218 597924
rect 331274 597868 331342 597924
rect 331398 597868 331494 597924
rect 330874 597800 331494 597868
rect 330874 597744 330970 597800
rect 331026 597744 331094 597800
rect 331150 597744 331218 597800
rect 331274 597744 331342 597800
rect 331398 597744 331494 597800
rect 330874 586350 331494 597744
rect 330874 586294 330970 586350
rect 331026 586294 331094 586350
rect 331150 586294 331218 586350
rect 331274 586294 331342 586350
rect 331398 586294 331494 586350
rect 330874 586226 331494 586294
rect 330874 586170 330970 586226
rect 331026 586170 331094 586226
rect 331150 586170 331218 586226
rect 331274 586170 331342 586226
rect 331398 586170 331494 586226
rect 330874 586102 331494 586170
rect 330874 586046 330970 586102
rect 331026 586046 331094 586102
rect 331150 586046 331218 586102
rect 331274 586046 331342 586102
rect 331398 586046 331494 586102
rect 330874 585978 331494 586046
rect 330874 585922 330970 585978
rect 331026 585922 331094 585978
rect 331150 585922 331218 585978
rect 331274 585922 331342 585978
rect 331398 585922 331494 585978
rect 330874 568350 331494 585922
rect 330874 568294 330970 568350
rect 331026 568294 331094 568350
rect 331150 568294 331218 568350
rect 331274 568294 331342 568350
rect 331398 568294 331494 568350
rect 330874 568226 331494 568294
rect 330874 568170 330970 568226
rect 331026 568170 331094 568226
rect 331150 568170 331218 568226
rect 331274 568170 331342 568226
rect 331398 568170 331494 568226
rect 330874 568102 331494 568170
rect 330874 568046 330970 568102
rect 331026 568046 331094 568102
rect 331150 568046 331218 568102
rect 331274 568046 331342 568102
rect 331398 568046 331494 568102
rect 330874 567978 331494 568046
rect 330874 567922 330970 567978
rect 331026 567922 331094 567978
rect 331150 567922 331218 567978
rect 331274 567922 331342 567978
rect 331398 567922 331494 567978
rect 330874 550350 331494 567922
rect 330874 550294 330970 550350
rect 331026 550294 331094 550350
rect 331150 550294 331218 550350
rect 331274 550294 331342 550350
rect 331398 550294 331494 550350
rect 330874 550226 331494 550294
rect 330874 550170 330970 550226
rect 331026 550170 331094 550226
rect 331150 550170 331218 550226
rect 331274 550170 331342 550226
rect 331398 550170 331494 550226
rect 330874 550102 331494 550170
rect 330874 550046 330970 550102
rect 331026 550046 331094 550102
rect 331150 550046 331218 550102
rect 331274 550046 331342 550102
rect 331398 550046 331494 550102
rect 330874 549978 331494 550046
rect 330874 549922 330970 549978
rect 331026 549922 331094 549978
rect 331150 549922 331218 549978
rect 331274 549922 331342 549978
rect 331398 549922 331494 549978
rect 330874 532350 331494 549922
rect 330874 532294 330970 532350
rect 331026 532294 331094 532350
rect 331150 532294 331218 532350
rect 331274 532294 331342 532350
rect 331398 532294 331494 532350
rect 330874 532226 331494 532294
rect 330874 532170 330970 532226
rect 331026 532170 331094 532226
rect 331150 532170 331218 532226
rect 331274 532170 331342 532226
rect 331398 532170 331494 532226
rect 330874 532102 331494 532170
rect 330874 532046 330970 532102
rect 331026 532046 331094 532102
rect 331150 532046 331218 532102
rect 331274 532046 331342 532102
rect 331398 532046 331494 532102
rect 330874 531978 331494 532046
rect 330874 531922 330970 531978
rect 331026 531922 331094 531978
rect 331150 531922 331218 531978
rect 331274 531922 331342 531978
rect 331398 531922 331494 531978
rect 330874 514350 331494 531922
rect 330874 514294 330970 514350
rect 331026 514294 331094 514350
rect 331150 514294 331218 514350
rect 331274 514294 331342 514350
rect 331398 514294 331494 514350
rect 330874 514226 331494 514294
rect 330874 514170 330970 514226
rect 331026 514170 331094 514226
rect 331150 514170 331218 514226
rect 331274 514170 331342 514226
rect 331398 514170 331494 514226
rect 330874 514102 331494 514170
rect 330874 514046 330970 514102
rect 331026 514046 331094 514102
rect 331150 514046 331218 514102
rect 331274 514046 331342 514102
rect 331398 514046 331494 514102
rect 330874 513978 331494 514046
rect 330874 513922 330970 513978
rect 331026 513922 331094 513978
rect 331150 513922 331218 513978
rect 331274 513922 331342 513978
rect 331398 513922 331494 513978
rect 330874 496350 331494 513922
rect 330874 496294 330970 496350
rect 331026 496294 331094 496350
rect 331150 496294 331218 496350
rect 331274 496294 331342 496350
rect 331398 496294 331494 496350
rect 330874 496226 331494 496294
rect 330874 496170 330970 496226
rect 331026 496170 331094 496226
rect 331150 496170 331218 496226
rect 331274 496170 331342 496226
rect 331398 496170 331494 496226
rect 330874 496102 331494 496170
rect 330874 496046 330970 496102
rect 331026 496046 331094 496102
rect 331150 496046 331218 496102
rect 331274 496046 331342 496102
rect 331398 496046 331494 496102
rect 330874 495978 331494 496046
rect 330874 495922 330970 495978
rect 331026 495922 331094 495978
rect 331150 495922 331218 495978
rect 331274 495922 331342 495978
rect 331398 495922 331494 495978
rect 330874 478350 331494 495922
rect 330874 478294 330970 478350
rect 331026 478294 331094 478350
rect 331150 478294 331218 478350
rect 331274 478294 331342 478350
rect 331398 478294 331494 478350
rect 330874 478226 331494 478294
rect 330874 478170 330970 478226
rect 331026 478170 331094 478226
rect 331150 478170 331218 478226
rect 331274 478170 331342 478226
rect 331398 478170 331494 478226
rect 330874 478102 331494 478170
rect 330874 478046 330970 478102
rect 331026 478046 331094 478102
rect 331150 478046 331218 478102
rect 331274 478046 331342 478102
rect 331398 478046 331494 478102
rect 330874 477978 331494 478046
rect 330874 477922 330970 477978
rect 331026 477922 331094 477978
rect 331150 477922 331218 477978
rect 331274 477922 331342 477978
rect 331398 477922 331494 477978
rect 330874 460350 331494 477922
rect 330874 460294 330970 460350
rect 331026 460294 331094 460350
rect 331150 460294 331218 460350
rect 331274 460294 331342 460350
rect 331398 460294 331494 460350
rect 330874 460226 331494 460294
rect 330874 460170 330970 460226
rect 331026 460170 331094 460226
rect 331150 460170 331218 460226
rect 331274 460170 331342 460226
rect 331398 460170 331494 460226
rect 330874 460102 331494 460170
rect 330874 460046 330970 460102
rect 331026 460046 331094 460102
rect 331150 460046 331218 460102
rect 331274 460046 331342 460102
rect 331398 460046 331494 460102
rect 330874 459978 331494 460046
rect 330874 459922 330970 459978
rect 331026 459922 331094 459978
rect 331150 459922 331218 459978
rect 331274 459922 331342 459978
rect 331398 459922 331494 459978
rect 330874 442350 331494 459922
rect 330874 442294 330970 442350
rect 331026 442294 331094 442350
rect 331150 442294 331218 442350
rect 331274 442294 331342 442350
rect 331398 442294 331494 442350
rect 330874 442226 331494 442294
rect 330874 442170 330970 442226
rect 331026 442170 331094 442226
rect 331150 442170 331218 442226
rect 331274 442170 331342 442226
rect 331398 442170 331494 442226
rect 330874 442102 331494 442170
rect 330874 442046 330970 442102
rect 331026 442046 331094 442102
rect 331150 442046 331218 442102
rect 331274 442046 331342 442102
rect 331398 442046 331494 442102
rect 330874 441978 331494 442046
rect 330874 441922 330970 441978
rect 331026 441922 331094 441978
rect 331150 441922 331218 441978
rect 331274 441922 331342 441978
rect 331398 441922 331494 441978
rect 330874 424350 331494 441922
rect 330874 424294 330970 424350
rect 331026 424294 331094 424350
rect 331150 424294 331218 424350
rect 331274 424294 331342 424350
rect 331398 424294 331494 424350
rect 330874 424226 331494 424294
rect 330874 424170 330970 424226
rect 331026 424170 331094 424226
rect 331150 424170 331218 424226
rect 331274 424170 331342 424226
rect 331398 424170 331494 424226
rect 330874 424102 331494 424170
rect 330874 424046 330970 424102
rect 331026 424046 331094 424102
rect 331150 424046 331218 424102
rect 331274 424046 331342 424102
rect 331398 424046 331494 424102
rect 330874 423978 331494 424046
rect 330874 423922 330970 423978
rect 331026 423922 331094 423978
rect 331150 423922 331218 423978
rect 331274 423922 331342 423978
rect 331398 423922 331494 423978
rect 330874 406350 331494 423922
rect 330874 406294 330970 406350
rect 331026 406294 331094 406350
rect 331150 406294 331218 406350
rect 331274 406294 331342 406350
rect 331398 406294 331494 406350
rect 330874 406226 331494 406294
rect 330874 406170 330970 406226
rect 331026 406170 331094 406226
rect 331150 406170 331218 406226
rect 331274 406170 331342 406226
rect 331398 406170 331494 406226
rect 330874 406102 331494 406170
rect 330874 406046 330970 406102
rect 331026 406046 331094 406102
rect 331150 406046 331218 406102
rect 331274 406046 331342 406102
rect 331398 406046 331494 406102
rect 330874 405978 331494 406046
rect 330874 405922 330970 405978
rect 331026 405922 331094 405978
rect 331150 405922 331218 405978
rect 331274 405922 331342 405978
rect 331398 405922 331494 405978
rect 330874 388350 331494 405922
rect 330874 388294 330970 388350
rect 331026 388294 331094 388350
rect 331150 388294 331218 388350
rect 331274 388294 331342 388350
rect 331398 388294 331494 388350
rect 330874 388226 331494 388294
rect 330874 388170 330970 388226
rect 331026 388170 331094 388226
rect 331150 388170 331218 388226
rect 331274 388170 331342 388226
rect 331398 388170 331494 388226
rect 330874 388102 331494 388170
rect 330874 388046 330970 388102
rect 331026 388046 331094 388102
rect 331150 388046 331218 388102
rect 331274 388046 331342 388102
rect 331398 388046 331494 388102
rect 330874 387978 331494 388046
rect 330874 387922 330970 387978
rect 331026 387922 331094 387978
rect 331150 387922 331218 387978
rect 331274 387922 331342 387978
rect 331398 387922 331494 387978
rect 330874 370350 331494 387922
rect 330874 370294 330970 370350
rect 331026 370294 331094 370350
rect 331150 370294 331218 370350
rect 331274 370294 331342 370350
rect 331398 370294 331494 370350
rect 330874 370226 331494 370294
rect 330874 370170 330970 370226
rect 331026 370170 331094 370226
rect 331150 370170 331218 370226
rect 331274 370170 331342 370226
rect 331398 370170 331494 370226
rect 330874 370102 331494 370170
rect 330874 370046 330970 370102
rect 331026 370046 331094 370102
rect 331150 370046 331218 370102
rect 331274 370046 331342 370102
rect 331398 370046 331494 370102
rect 330874 369978 331494 370046
rect 330874 369922 330970 369978
rect 331026 369922 331094 369978
rect 331150 369922 331218 369978
rect 331274 369922 331342 369978
rect 331398 369922 331494 369978
rect 330874 352350 331494 369922
rect 330874 352294 330970 352350
rect 331026 352294 331094 352350
rect 331150 352294 331218 352350
rect 331274 352294 331342 352350
rect 331398 352294 331494 352350
rect 330874 352226 331494 352294
rect 330874 352170 330970 352226
rect 331026 352170 331094 352226
rect 331150 352170 331218 352226
rect 331274 352170 331342 352226
rect 331398 352170 331494 352226
rect 330874 352102 331494 352170
rect 330874 352046 330970 352102
rect 331026 352046 331094 352102
rect 331150 352046 331218 352102
rect 331274 352046 331342 352102
rect 331398 352046 331494 352102
rect 330874 351978 331494 352046
rect 330874 351922 330970 351978
rect 331026 351922 331094 351978
rect 331150 351922 331218 351978
rect 331274 351922 331342 351978
rect 331398 351922 331494 351978
rect 330874 334350 331494 351922
rect 330874 334294 330970 334350
rect 331026 334294 331094 334350
rect 331150 334294 331218 334350
rect 331274 334294 331342 334350
rect 331398 334294 331494 334350
rect 330874 334226 331494 334294
rect 330874 334170 330970 334226
rect 331026 334170 331094 334226
rect 331150 334170 331218 334226
rect 331274 334170 331342 334226
rect 331398 334170 331494 334226
rect 330874 334102 331494 334170
rect 330874 334046 330970 334102
rect 331026 334046 331094 334102
rect 331150 334046 331218 334102
rect 331274 334046 331342 334102
rect 331398 334046 331494 334102
rect 330874 333978 331494 334046
rect 330874 333922 330970 333978
rect 331026 333922 331094 333978
rect 331150 333922 331218 333978
rect 331274 333922 331342 333978
rect 331398 333922 331494 333978
rect 330874 316350 331494 333922
rect 330874 316294 330970 316350
rect 331026 316294 331094 316350
rect 331150 316294 331218 316350
rect 331274 316294 331342 316350
rect 331398 316294 331494 316350
rect 330874 316226 331494 316294
rect 330874 316170 330970 316226
rect 331026 316170 331094 316226
rect 331150 316170 331218 316226
rect 331274 316170 331342 316226
rect 331398 316170 331494 316226
rect 330874 316102 331494 316170
rect 330874 316046 330970 316102
rect 331026 316046 331094 316102
rect 331150 316046 331218 316102
rect 331274 316046 331342 316102
rect 331398 316046 331494 316102
rect 330874 315978 331494 316046
rect 330874 315922 330970 315978
rect 331026 315922 331094 315978
rect 331150 315922 331218 315978
rect 331274 315922 331342 315978
rect 331398 315922 331494 315978
rect 330874 298350 331494 315922
rect 330874 298294 330970 298350
rect 331026 298294 331094 298350
rect 331150 298294 331218 298350
rect 331274 298294 331342 298350
rect 331398 298294 331494 298350
rect 330874 298226 331494 298294
rect 330874 298170 330970 298226
rect 331026 298170 331094 298226
rect 331150 298170 331218 298226
rect 331274 298170 331342 298226
rect 331398 298170 331494 298226
rect 330874 298102 331494 298170
rect 330874 298046 330970 298102
rect 331026 298046 331094 298102
rect 331150 298046 331218 298102
rect 331274 298046 331342 298102
rect 331398 298046 331494 298102
rect 330874 297978 331494 298046
rect 330874 297922 330970 297978
rect 331026 297922 331094 297978
rect 331150 297922 331218 297978
rect 331274 297922 331342 297978
rect 331398 297922 331494 297978
rect 330874 280350 331494 297922
rect 330874 280294 330970 280350
rect 331026 280294 331094 280350
rect 331150 280294 331218 280350
rect 331274 280294 331342 280350
rect 331398 280294 331494 280350
rect 330874 280226 331494 280294
rect 330874 280170 330970 280226
rect 331026 280170 331094 280226
rect 331150 280170 331218 280226
rect 331274 280170 331342 280226
rect 331398 280170 331494 280226
rect 330874 280102 331494 280170
rect 330874 280046 330970 280102
rect 331026 280046 331094 280102
rect 331150 280046 331218 280102
rect 331274 280046 331342 280102
rect 331398 280046 331494 280102
rect 330874 279978 331494 280046
rect 330874 279922 330970 279978
rect 331026 279922 331094 279978
rect 331150 279922 331218 279978
rect 331274 279922 331342 279978
rect 331398 279922 331494 279978
rect 330874 262350 331494 279922
rect 330874 262294 330970 262350
rect 331026 262294 331094 262350
rect 331150 262294 331218 262350
rect 331274 262294 331342 262350
rect 331398 262294 331494 262350
rect 330874 262226 331494 262294
rect 330874 262170 330970 262226
rect 331026 262170 331094 262226
rect 331150 262170 331218 262226
rect 331274 262170 331342 262226
rect 331398 262170 331494 262226
rect 330874 262102 331494 262170
rect 330874 262046 330970 262102
rect 331026 262046 331094 262102
rect 331150 262046 331218 262102
rect 331274 262046 331342 262102
rect 331398 262046 331494 262102
rect 330874 261978 331494 262046
rect 330874 261922 330970 261978
rect 331026 261922 331094 261978
rect 331150 261922 331218 261978
rect 331274 261922 331342 261978
rect 331398 261922 331494 261978
rect 330874 244350 331494 261922
rect 330874 244294 330970 244350
rect 331026 244294 331094 244350
rect 331150 244294 331218 244350
rect 331274 244294 331342 244350
rect 331398 244294 331494 244350
rect 330874 244226 331494 244294
rect 330874 244170 330970 244226
rect 331026 244170 331094 244226
rect 331150 244170 331218 244226
rect 331274 244170 331342 244226
rect 331398 244170 331494 244226
rect 330874 244102 331494 244170
rect 330874 244046 330970 244102
rect 331026 244046 331094 244102
rect 331150 244046 331218 244102
rect 331274 244046 331342 244102
rect 331398 244046 331494 244102
rect 330874 243978 331494 244046
rect 330874 243922 330970 243978
rect 331026 243922 331094 243978
rect 331150 243922 331218 243978
rect 331274 243922 331342 243978
rect 331398 243922 331494 243978
rect 330874 226350 331494 243922
rect 348874 598172 349494 598268
rect 348874 598116 348970 598172
rect 349026 598116 349094 598172
rect 349150 598116 349218 598172
rect 349274 598116 349342 598172
rect 349398 598116 349494 598172
rect 348874 598048 349494 598116
rect 348874 597992 348970 598048
rect 349026 597992 349094 598048
rect 349150 597992 349218 598048
rect 349274 597992 349342 598048
rect 349398 597992 349494 598048
rect 348874 597924 349494 597992
rect 348874 597868 348970 597924
rect 349026 597868 349094 597924
rect 349150 597868 349218 597924
rect 349274 597868 349342 597924
rect 349398 597868 349494 597924
rect 348874 597800 349494 597868
rect 348874 597744 348970 597800
rect 349026 597744 349094 597800
rect 349150 597744 349218 597800
rect 349274 597744 349342 597800
rect 349398 597744 349494 597800
rect 348874 586350 349494 597744
rect 348874 586294 348970 586350
rect 349026 586294 349094 586350
rect 349150 586294 349218 586350
rect 349274 586294 349342 586350
rect 349398 586294 349494 586350
rect 348874 586226 349494 586294
rect 348874 586170 348970 586226
rect 349026 586170 349094 586226
rect 349150 586170 349218 586226
rect 349274 586170 349342 586226
rect 349398 586170 349494 586226
rect 348874 586102 349494 586170
rect 348874 586046 348970 586102
rect 349026 586046 349094 586102
rect 349150 586046 349218 586102
rect 349274 586046 349342 586102
rect 349398 586046 349494 586102
rect 348874 585978 349494 586046
rect 348874 585922 348970 585978
rect 349026 585922 349094 585978
rect 349150 585922 349218 585978
rect 349274 585922 349342 585978
rect 349398 585922 349494 585978
rect 348874 568350 349494 585922
rect 348874 568294 348970 568350
rect 349026 568294 349094 568350
rect 349150 568294 349218 568350
rect 349274 568294 349342 568350
rect 349398 568294 349494 568350
rect 348874 568226 349494 568294
rect 348874 568170 348970 568226
rect 349026 568170 349094 568226
rect 349150 568170 349218 568226
rect 349274 568170 349342 568226
rect 349398 568170 349494 568226
rect 348874 568102 349494 568170
rect 348874 568046 348970 568102
rect 349026 568046 349094 568102
rect 349150 568046 349218 568102
rect 349274 568046 349342 568102
rect 349398 568046 349494 568102
rect 348874 567978 349494 568046
rect 348874 567922 348970 567978
rect 349026 567922 349094 567978
rect 349150 567922 349218 567978
rect 349274 567922 349342 567978
rect 349398 567922 349494 567978
rect 348874 550350 349494 567922
rect 348874 550294 348970 550350
rect 349026 550294 349094 550350
rect 349150 550294 349218 550350
rect 349274 550294 349342 550350
rect 349398 550294 349494 550350
rect 348874 550226 349494 550294
rect 348874 550170 348970 550226
rect 349026 550170 349094 550226
rect 349150 550170 349218 550226
rect 349274 550170 349342 550226
rect 349398 550170 349494 550226
rect 348874 550102 349494 550170
rect 348874 550046 348970 550102
rect 349026 550046 349094 550102
rect 349150 550046 349218 550102
rect 349274 550046 349342 550102
rect 349398 550046 349494 550102
rect 348874 549978 349494 550046
rect 348874 549922 348970 549978
rect 349026 549922 349094 549978
rect 349150 549922 349218 549978
rect 349274 549922 349342 549978
rect 349398 549922 349494 549978
rect 348874 532350 349494 549922
rect 348874 532294 348970 532350
rect 349026 532294 349094 532350
rect 349150 532294 349218 532350
rect 349274 532294 349342 532350
rect 349398 532294 349494 532350
rect 348874 532226 349494 532294
rect 348874 532170 348970 532226
rect 349026 532170 349094 532226
rect 349150 532170 349218 532226
rect 349274 532170 349342 532226
rect 349398 532170 349494 532226
rect 348874 532102 349494 532170
rect 348874 532046 348970 532102
rect 349026 532046 349094 532102
rect 349150 532046 349218 532102
rect 349274 532046 349342 532102
rect 349398 532046 349494 532102
rect 348874 531978 349494 532046
rect 348874 531922 348970 531978
rect 349026 531922 349094 531978
rect 349150 531922 349218 531978
rect 349274 531922 349342 531978
rect 349398 531922 349494 531978
rect 348874 514350 349494 531922
rect 348874 514294 348970 514350
rect 349026 514294 349094 514350
rect 349150 514294 349218 514350
rect 349274 514294 349342 514350
rect 349398 514294 349494 514350
rect 348874 514226 349494 514294
rect 348874 514170 348970 514226
rect 349026 514170 349094 514226
rect 349150 514170 349218 514226
rect 349274 514170 349342 514226
rect 349398 514170 349494 514226
rect 348874 514102 349494 514170
rect 348874 514046 348970 514102
rect 349026 514046 349094 514102
rect 349150 514046 349218 514102
rect 349274 514046 349342 514102
rect 349398 514046 349494 514102
rect 348874 513978 349494 514046
rect 348874 513922 348970 513978
rect 349026 513922 349094 513978
rect 349150 513922 349218 513978
rect 349274 513922 349342 513978
rect 349398 513922 349494 513978
rect 348874 496350 349494 513922
rect 348874 496294 348970 496350
rect 349026 496294 349094 496350
rect 349150 496294 349218 496350
rect 349274 496294 349342 496350
rect 349398 496294 349494 496350
rect 348874 496226 349494 496294
rect 348874 496170 348970 496226
rect 349026 496170 349094 496226
rect 349150 496170 349218 496226
rect 349274 496170 349342 496226
rect 349398 496170 349494 496226
rect 348874 496102 349494 496170
rect 348874 496046 348970 496102
rect 349026 496046 349094 496102
rect 349150 496046 349218 496102
rect 349274 496046 349342 496102
rect 349398 496046 349494 496102
rect 348874 495978 349494 496046
rect 348874 495922 348970 495978
rect 349026 495922 349094 495978
rect 349150 495922 349218 495978
rect 349274 495922 349342 495978
rect 349398 495922 349494 495978
rect 348874 478350 349494 495922
rect 348874 478294 348970 478350
rect 349026 478294 349094 478350
rect 349150 478294 349218 478350
rect 349274 478294 349342 478350
rect 349398 478294 349494 478350
rect 348874 478226 349494 478294
rect 348874 478170 348970 478226
rect 349026 478170 349094 478226
rect 349150 478170 349218 478226
rect 349274 478170 349342 478226
rect 349398 478170 349494 478226
rect 348874 478102 349494 478170
rect 348874 478046 348970 478102
rect 349026 478046 349094 478102
rect 349150 478046 349218 478102
rect 349274 478046 349342 478102
rect 349398 478046 349494 478102
rect 348874 477978 349494 478046
rect 348874 477922 348970 477978
rect 349026 477922 349094 477978
rect 349150 477922 349218 477978
rect 349274 477922 349342 477978
rect 349398 477922 349494 477978
rect 348874 460350 349494 477922
rect 348874 460294 348970 460350
rect 349026 460294 349094 460350
rect 349150 460294 349218 460350
rect 349274 460294 349342 460350
rect 349398 460294 349494 460350
rect 348874 460226 349494 460294
rect 348874 460170 348970 460226
rect 349026 460170 349094 460226
rect 349150 460170 349218 460226
rect 349274 460170 349342 460226
rect 349398 460170 349494 460226
rect 348874 460102 349494 460170
rect 348874 460046 348970 460102
rect 349026 460046 349094 460102
rect 349150 460046 349218 460102
rect 349274 460046 349342 460102
rect 349398 460046 349494 460102
rect 348874 459978 349494 460046
rect 348874 459922 348970 459978
rect 349026 459922 349094 459978
rect 349150 459922 349218 459978
rect 349274 459922 349342 459978
rect 349398 459922 349494 459978
rect 348874 442350 349494 459922
rect 348874 442294 348970 442350
rect 349026 442294 349094 442350
rect 349150 442294 349218 442350
rect 349274 442294 349342 442350
rect 349398 442294 349494 442350
rect 348874 442226 349494 442294
rect 348874 442170 348970 442226
rect 349026 442170 349094 442226
rect 349150 442170 349218 442226
rect 349274 442170 349342 442226
rect 349398 442170 349494 442226
rect 348874 442102 349494 442170
rect 348874 442046 348970 442102
rect 349026 442046 349094 442102
rect 349150 442046 349218 442102
rect 349274 442046 349342 442102
rect 349398 442046 349494 442102
rect 348874 441978 349494 442046
rect 348874 441922 348970 441978
rect 349026 441922 349094 441978
rect 349150 441922 349218 441978
rect 349274 441922 349342 441978
rect 349398 441922 349494 441978
rect 348874 424350 349494 441922
rect 348874 424294 348970 424350
rect 349026 424294 349094 424350
rect 349150 424294 349218 424350
rect 349274 424294 349342 424350
rect 349398 424294 349494 424350
rect 348874 424226 349494 424294
rect 348874 424170 348970 424226
rect 349026 424170 349094 424226
rect 349150 424170 349218 424226
rect 349274 424170 349342 424226
rect 349398 424170 349494 424226
rect 348874 424102 349494 424170
rect 348874 424046 348970 424102
rect 349026 424046 349094 424102
rect 349150 424046 349218 424102
rect 349274 424046 349342 424102
rect 349398 424046 349494 424102
rect 348874 423978 349494 424046
rect 348874 423922 348970 423978
rect 349026 423922 349094 423978
rect 349150 423922 349218 423978
rect 349274 423922 349342 423978
rect 349398 423922 349494 423978
rect 348874 406350 349494 423922
rect 348874 406294 348970 406350
rect 349026 406294 349094 406350
rect 349150 406294 349218 406350
rect 349274 406294 349342 406350
rect 349398 406294 349494 406350
rect 348874 406226 349494 406294
rect 348874 406170 348970 406226
rect 349026 406170 349094 406226
rect 349150 406170 349218 406226
rect 349274 406170 349342 406226
rect 349398 406170 349494 406226
rect 348874 406102 349494 406170
rect 348874 406046 348970 406102
rect 349026 406046 349094 406102
rect 349150 406046 349218 406102
rect 349274 406046 349342 406102
rect 349398 406046 349494 406102
rect 348874 405978 349494 406046
rect 348874 405922 348970 405978
rect 349026 405922 349094 405978
rect 349150 405922 349218 405978
rect 349274 405922 349342 405978
rect 349398 405922 349494 405978
rect 348874 388350 349494 405922
rect 348874 388294 348970 388350
rect 349026 388294 349094 388350
rect 349150 388294 349218 388350
rect 349274 388294 349342 388350
rect 349398 388294 349494 388350
rect 348874 388226 349494 388294
rect 348874 388170 348970 388226
rect 349026 388170 349094 388226
rect 349150 388170 349218 388226
rect 349274 388170 349342 388226
rect 349398 388170 349494 388226
rect 348874 388102 349494 388170
rect 348874 388046 348970 388102
rect 349026 388046 349094 388102
rect 349150 388046 349218 388102
rect 349274 388046 349342 388102
rect 349398 388046 349494 388102
rect 348874 387978 349494 388046
rect 348874 387922 348970 387978
rect 349026 387922 349094 387978
rect 349150 387922 349218 387978
rect 349274 387922 349342 387978
rect 349398 387922 349494 387978
rect 348874 370350 349494 387922
rect 348874 370294 348970 370350
rect 349026 370294 349094 370350
rect 349150 370294 349218 370350
rect 349274 370294 349342 370350
rect 349398 370294 349494 370350
rect 348874 370226 349494 370294
rect 348874 370170 348970 370226
rect 349026 370170 349094 370226
rect 349150 370170 349218 370226
rect 349274 370170 349342 370226
rect 349398 370170 349494 370226
rect 348874 370102 349494 370170
rect 348874 370046 348970 370102
rect 349026 370046 349094 370102
rect 349150 370046 349218 370102
rect 349274 370046 349342 370102
rect 349398 370046 349494 370102
rect 348874 369978 349494 370046
rect 348874 369922 348970 369978
rect 349026 369922 349094 369978
rect 349150 369922 349218 369978
rect 349274 369922 349342 369978
rect 349398 369922 349494 369978
rect 348874 352350 349494 369922
rect 348874 352294 348970 352350
rect 349026 352294 349094 352350
rect 349150 352294 349218 352350
rect 349274 352294 349342 352350
rect 349398 352294 349494 352350
rect 348874 352226 349494 352294
rect 348874 352170 348970 352226
rect 349026 352170 349094 352226
rect 349150 352170 349218 352226
rect 349274 352170 349342 352226
rect 349398 352170 349494 352226
rect 348874 352102 349494 352170
rect 348874 352046 348970 352102
rect 349026 352046 349094 352102
rect 349150 352046 349218 352102
rect 349274 352046 349342 352102
rect 349398 352046 349494 352102
rect 348874 351978 349494 352046
rect 348874 351922 348970 351978
rect 349026 351922 349094 351978
rect 349150 351922 349218 351978
rect 349274 351922 349342 351978
rect 349398 351922 349494 351978
rect 348874 334350 349494 351922
rect 348874 334294 348970 334350
rect 349026 334294 349094 334350
rect 349150 334294 349218 334350
rect 349274 334294 349342 334350
rect 349398 334294 349494 334350
rect 348874 334226 349494 334294
rect 348874 334170 348970 334226
rect 349026 334170 349094 334226
rect 349150 334170 349218 334226
rect 349274 334170 349342 334226
rect 349398 334170 349494 334226
rect 348874 334102 349494 334170
rect 348874 334046 348970 334102
rect 349026 334046 349094 334102
rect 349150 334046 349218 334102
rect 349274 334046 349342 334102
rect 349398 334046 349494 334102
rect 348874 333978 349494 334046
rect 348874 333922 348970 333978
rect 349026 333922 349094 333978
rect 349150 333922 349218 333978
rect 349274 333922 349342 333978
rect 349398 333922 349494 333978
rect 348874 316350 349494 333922
rect 348874 316294 348970 316350
rect 349026 316294 349094 316350
rect 349150 316294 349218 316350
rect 349274 316294 349342 316350
rect 349398 316294 349494 316350
rect 348874 316226 349494 316294
rect 348874 316170 348970 316226
rect 349026 316170 349094 316226
rect 349150 316170 349218 316226
rect 349274 316170 349342 316226
rect 349398 316170 349494 316226
rect 348874 316102 349494 316170
rect 348874 316046 348970 316102
rect 349026 316046 349094 316102
rect 349150 316046 349218 316102
rect 349274 316046 349342 316102
rect 349398 316046 349494 316102
rect 348874 315978 349494 316046
rect 348874 315922 348970 315978
rect 349026 315922 349094 315978
rect 349150 315922 349218 315978
rect 349274 315922 349342 315978
rect 349398 315922 349494 315978
rect 348874 298350 349494 315922
rect 348874 298294 348970 298350
rect 349026 298294 349094 298350
rect 349150 298294 349218 298350
rect 349274 298294 349342 298350
rect 349398 298294 349494 298350
rect 348874 298226 349494 298294
rect 348874 298170 348970 298226
rect 349026 298170 349094 298226
rect 349150 298170 349218 298226
rect 349274 298170 349342 298226
rect 349398 298170 349494 298226
rect 348874 298102 349494 298170
rect 348874 298046 348970 298102
rect 349026 298046 349094 298102
rect 349150 298046 349218 298102
rect 349274 298046 349342 298102
rect 349398 298046 349494 298102
rect 348874 297978 349494 298046
rect 348874 297922 348970 297978
rect 349026 297922 349094 297978
rect 349150 297922 349218 297978
rect 349274 297922 349342 297978
rect 349398 297922 349494 297978
rect 348874 280350 349494 297922
rect 348874 280294 348970 280350
rect 349026 280294 349094 280350
rect 349150 280294 349218 280350
rect 349274 280294 349342 280350
rect 349398 280294 349494 280350
rect 348874 280226 349494 280294
rect 348874 280170 348970 280226
rect 349026 280170 349094 280226
rect 349150 280170 349218 280226
rect 349274 280170 349342 280226
rect 349398 280170 349494 280226
rect 348874 280102 349494 280170
rect 348874 280046 348970 280102
rect 349026 280046 349094 280102
rect 349150 280046 349218 280102
rect 349274 280046 349342 280102
rect 349398 280046 349494 280102
rect 348874 279978 349494 280046
rect 348874 279922 348970 279978
rect 349026 279922 349094 279978
rect 349150 279922 349218 279978
rect 349274 279922 349342 279978
rect 349398 279922 349494 279978
rect 348874 262350 349494 279922
rect 348874 262294 348970 262350
rect 349026 262294 349094 262350
rect 349150 262294 349218 262350
rect 349274 262294 349342 262350
rect 349398 262294 349494 262350
rect 348874 262226 349494 262294
rect 348874 262170 348970 262226
rect 349026 262170 349094 262226
rect 349150 262170 349218 262226
rect 349274 262170 349342 262226
rect 349398 262170 349494 262226
rect 348874 262102 349494 262170
rect 348874 262046 348970 262102
rect 349026 262046 349094 262102
rect 349150 262046 349218 262102
rect 349274 262046 349342 262102
rect 349398 262046 349494 262102
rect 348874 261978 349494 262046
rect 348874 261922 348970 261978
rect 349026 261922 349094 261978
rect 349150 261922 349218 261978
rect 349274 261922 349342 261978
rect 349398 261922 349494 261978
rect 348874 244350 349494 261922
rect 348874 244294 348970 244350
rect 349026 244294 349094 244350
rect 349150 244294 349218 244350
rect 349274 244294 349342 244350
rect 349398 244294 349494 244350
rect 348874 244226 349494 244294
rect 348874 244170 348970 244226
rect 349026 244170 349094 244226
rect 349150 244170 349218 244226
rect 349274 244170 349342 244226
rect 349398 244170 349494 244226
rect 348874 244102 349494 244170
rect 348874 244046 348970 244102
rect 349026 244046 349094 244102
rect 349150 244046 349218 244102
rect 349274 244046 349342 244102
rect 349398 244046 349494 244102
rect 348874 243978 349494 244046
rect 348874 243922 348970 243978
rect 349026 243922 349094 243978
rect 349150 243922 349218 243978
rect 349274 243922 349342 243978
rect 349398 243922 349494 243978
rect 330874 226294 330970 226350
rect 331026 226294 331094 226350
rect 331150 226294 331218 226350
rect 331274 226294 331342 226350
rect 331398 226294 331494 226350
rect 330874 226226 331494 226294
rect 330874 226170 330970 226226
rect 331026 226170 331094 226226
rect 331150 226170 331218 226226
rect 331274 226170 331342 226226
rect 331398 226170 331494 226226
rect 330874 226102 331494 226170
rect 330874 226046 330970 226102
rect 331026 226046 331094 226102
rect 331150 226046 331218 226102
rect 331274 226046 331342 226102
rect 331398 226046 331494 226102
rect 330874 225978 331494 226046
rect 330874 225922 330970 225978
rect 331026 225922 331094 225978
rect 331150 225922 331218 225978
rect 331274 225922 331342 225978
rect 331398 225922 331494 225978
rect 330874 208350 331494 225922
rect 330874 208294 330970 208350
rect 331026 208294 331094 208350
rect 331150 208294 331218 208350
rect 331274 208294 331342 208350
rect 331398 208294 331494 208350
rect 330874 208226 331494 208294
rect 330874 208170 330970 208226
rect 331026 208170 331094 208226
rect 331150 208170 331218 208226
rect 331274 208170 331342 208226
rect 331398 208170 331494 208226
rect 330874 208102 331494 208170
rect 330874 208046 330970 208102
rect 331026 208046 331094 208102
rect 331150 208046 331218 208102
rect 331274 208046 331342 208102
rect 331398 208046 331494 208102
rect 330874 207978 331494 208046
rect 330874 207922 330970 207978
rect 331026 207922 331094 207978
rect 331150 207922 331218 207978
rect 331274 207922 331342 207978
rect 331398 207922 331494 207978
rect 330874 190350 331494 207922
rect 330874 190294 330970 190350
rect 331026 190294 331094 190350
rect 331150 190294 331218 190350
rect 331274 190294 331342 190350
rect 331398 190294 331494 190350
rect 330874 190226 331494 190294
rect 330874 190170 330970 190226
rect 331026 190170 331094 190226
rect 331150 190170 331218 190226
rect 331274 190170 331342 190226
rect 331398 190170 331494 190226
rect 330874 190102 331494 190170
rect 330874 190046 330970 190102
rect 331026 190046 331094 190102
rect 331150 190046 331218 190102
rect 331274 190046 331342 190102
rect 331398 190046 331494 190102
rect 330874 189978 331494 190046
rect 330874 189922 330970 189978
rect 331026 189922 331094 189978
rect 331150 189922 331218 189978
rect 331274 189922 331342 189978
rect 331398 189922 331494 189978
rect 330874 172350 331494 189922
rect 330874 172294 330970 172350
rect 331026 172294 331094 172350
rect 331150 172294 331218 172350
rect 331274 172294 331342 172350
rect 331398 172294 331494 172350
rect 330874 172226 331494 172294
rect 330874 172170 330970 172226
rect 331026 172170 331094 172226
rect 331150 172170 331218 172226
rect 331274 172170 331342 172226
rect 331398 172170 331494 172226
rect 330874 172102 331494 172170
rect 330874 172046 330970 172102
rect 331026 172046 331094 172102
rect 331150 172046 331218 172102
rect 331274 172046 331342 172102
rect 331398 172046 331494 172102
rect 330874 171978 331494 172046
rect 330874 171922 330970 171978
rect 331026 171922 331094 171978
rect 331150 171922 331218 171978
rect 331274 171922 331342 171978
rect 331398 171922 331494 171978
rect 330874 154350 331494 171922
rect 330874 154294 330970 154350
rect 331026 154294 331094 154350
rect 331150 154294 331218 154350
rect 331274 154294 331342 154350
rect 331398 154294 331494 154350
rect 330874 154226 331494 154294
rect 330874 154170 330970 154226
rect 331026 154170 331094 154226
rect 331150 154170 331218 154226
rect 331274 154170 331342 154226
rect 331398 154170 331494 154226
rect 330874 154102 331494 154170
rect 330874 154046 330970 154102
rect 331026 154046 331094 154102
rect 331150 154046 331218 154102
rect 331274 154046 331342 154102
rect 331398 154046 331494 154102
rect 330874 153978 331494 154046
rect 330874 153922 330970 153978
rect 331026 153922 331094 153978
rect 331150 153922 331218 153978
rect 331274 153922 331342 153978
rect 331398 153922 331494 153978
rect 330874 136350 331494 153922
rect 330874 136294 330970 136350
rect 331026 136294 331094 136350
rect 331150 136294 331218 136350
rect 331274 136294 331342 136350
rect 331398 136294 331494 136350
rect 330874 136226 331494 136294
rect 330874 136170 330970 136226
rect 331026 136170 331094 136226
rect 331150 136170 331218 136226
rect 331274 136170 331342 136226
rect 331398 136170 331494 136226
rect 330874 136102 331494 136170
rect 330874 136046 330970 136102
rect 331026 136046 331094 136102
rect 331150 136046 331218 136102
rect 331274 136046 331342 136102
rect 331398 136046 331494 136102
rect 330874 135978 331494 136046
rect 330874 135922 330970 135978
rect 331026 135922 331094 135978
rect 331150 135922 331218 135978
rect 331274 135922 331342 135978
rect 331398 135922 331494 135978
rect 330874 118350 331494 135922
rect 330874 118294 330970 118350
rect 331026 118294 331094 118350
rect 331150 118294 331218 118350
rect 331274 118294 331342 118350
rect 331398 118294 331494 118350
rect 330874 118226 331494 118294
rect 330874 118170 330970 118226
rect 331026 118170 331094 118226
rect 331150 118170 331218 118226
rect 331274 118170 331342 118226
rect 331398 118170 331494 118226
rect 330874 118102 331494 118170
rect 330874 118046 330970 118102
rect 331026 118046 331094 118102
rect 331150 118046 331218 118102
rect 331274 118046 331342 118102
rect 331398 118046 331494 118102
rect 330874 117978 331494 118046
rect 330874 117922 330970 117978
rect 331026 117922 331094 117978
rect 331150 117922 331218 117978
rect 331274 117922 331342 117978
rect 331398 117922 331494 117978
rect 330874 100350 331494 117922
rect 330874 100294 330970 100350
rect 331026 100294 331094 100350
rect 331150 100294 331218 100350
rect 331274 100294 331342 100350
rect 331398 100294 331494 100350
rect 330874 100226 331494 100294
rect 330874 100170 330970 100226
rect 331026 100170 331094 100226
rect 331150 100170 331218 100226
rect 331274 100170 331342 100226
rect 331398 100170 331494 100226
rect 330874 100102 331494 100170
rect 330874 100046 330970 100102
rect 331026 100046 331094 100102
rect 331150 100046 331218 100102
rect 331274 100046 331342 100102
rect 331398 100046 331494 100102
rect 330874 99978 331494 100046
rect 330874 99922 330970 99978
rect 331026 99922 331094 99978
rect 331150 99922 331218 99978
rect 331274 99922 331342 99978
rect 331398 99922 331494 99978
rect 330874 82350 331494 99922
rect 330874 82294 330970 82350
rect 331026 82294 331094 82350
rect 331150 82294 331218 82350
rect 331274 82294 331342 82350
rect 331398 82294 331494 82350
rect 330874 82226 331494 82294
rect 330874 82170 330970 82226
rect 331026 82170 331094 82226
rect 331150 82170 331218 82226
rect 331274 82170 331342 82226
rect 331398 82170 331494 82226
rect 330874 82102 331494 82170
rect 330874 82046 330970 82102
rect 331026 82046 331094 82102
rect 331150 82046 331218 82102
rect 331274 82046 331342 82102
rect 331398 82046 331494 82102
rect 330874 81978 331494 82046
rect 330874 81922 330970 81978
rect 331026 81922 331094 81978
rect 331150 81922 331218 81978
rect 331274 81922 331342 81978
rect 331398 81922 331494 81978
rect 330874 64350 331494 81922
rect 330874 64294 330970 64350
rect 331026 64294 331094 64350
rect 331150 64294 331218 64350
rect 331274 64294 331342 64350
rect 331398 64294 331494 64350
rect 330874 64226 331494 64294
rect 330874 64170 330970 64226
rect 331026 64170 331094 64226
rect 331150 64170 331218 64226
rect 331274 64170 331342 64226
rect 331398 64170 331494 64226
rect 330874 64102 331494 64170
rect 330874 64046 330970 64102
rect 331026 64046 331094 64102
rect 331150 64046 331218 64102
rect 331274 64046 331342 64102
rect 331398 64046 331494 64102
rect 330874 63978 331494 64046
rect 330874 63922 330970 63978
rect 331026 63922 331094 63978
rect 331150 63922 331218 63978
rect 331274 63922 331342 63978
rect 331398 63922 331494 63978
rect 330874 46350 331494 63922
rect 345154 238350 345774 242964
rect 345154 238294 345250 238350
rect 345306 238294 345374 238350
rect 345430 238294 345498 238350
rect 345554 238294 345622 238350
rect 345678 238294 345774 238350
rect 345154 238226 345774 238294
rect 345154 238170 345250 238226
rect 345306 238170 345374 238226
rect 345430 238170 345498 238226
rect 345554 238170 345622 238226
rect 345678 238170 345774 238226
rect 345154 238102 345774 238170
rect 345154 238046 345250 238102
rect 345306 238046 345374 238102
rect 345430 238046 345498 238102
rect 345554 238046 345622 238102
rect 345678 238046 345774 238102
rect 345154 237978 345774 238046
rect 345154 237922 345250 237978
rect 345306 237922 345374 237978
rect 345430 237922 345498 237978
rect 345554 237922 345622 237978
rect 345678 237922 345774 237978
rect 345154 220350 345774 237922
rect 345154 220294 345250 220350
rect 345306 220294 345374 220350
rect 345430 220294 345498 220350
rect 345554 220294 345622 220350
rect 345678 220294 345774 220350
rect 345154 220226 345774 220294
rect 345154 220170 345250 220226
rect 345306 220170 345374 220226
rect 345430 220170 345498 220226
rect 345554 220170 345622 220226
rect 345678 220170 345774 220226
rect 345154 220102 345774 220170
rect 345154 220046 345250 220102
rect 345306 220046 345374 220102
rect 345430 220046 345498 220102
rect 345554 220046 345622 220102
rect 345678 220046 345774 220102
rect 345154 219978 345774 220046
rect 345154 219922 345250 219978
rect 345306 219922 345374 219978
rect 345430 219922 345498 219978
rect 345554 219922 345622 219978
rect 345678 219922 345774 219978
rect 345154 202350 345774 219922
rect 345154 202294 345250 202350
rect 345306 202294 345374 202350
rect 345430 202294 345498 202350
rect 345554 202294 345622 202350
rect 345678 202294 345774 202350
rect 345154 202226 345774 202294
rect 345154 202170 345250 202226
rect 345306 202170 345374 202226
rect 345430 202170 345498 202226
rect 345554 202170 345622 202226
rect 345678 202170 345774 202226
rect 345154 202102 345774 202170
rect 345154 202046 345250 202102
rect 345306 202046 345374 202102
rect 345430 202046 345498 202102
rect 345554 202046 345622 202102
rect 345678 202046 345774 202102
rect 345154 201978 345774 202046
rect 345154 201922 345250 201978
rect 345306 201922 345374 201978
rect 345430 201922 345498 201978
rect 345554 201922 345622 201978
rect 345678 201922 345774 201978
rect 345154 184350 345774 201922
rect 345154 184294 345250 184350
rect 345306 184294 345374 184350
rect 345430 184294 345498 184350
rect 345554 184294 345622 184350
rect 345678 184294 345774 184350
rect 345154 184226 345774 184294
rect 345154 184170 345250 184226
rect 345306 184170 345374 184226
rect 345430 184170 345498 184226
rect 345554 184170 345622 184226
rect 345678 184170 345774 184226
rect 345154 184102 345774 184170
rect 345154 184046 345250 184102
rect 345306 184046 345374 184102
rect 345430 184046 345498 184102
rect 345554 184046 345622 184102
rect 345678 184046 345774 184102
rect 345154 183978 345774 184046
rect 345154 183922 345250 183978
rect 345306 183922 345374 183978
rect 345430 183922 345498 183978
rect 345554 183922 345622 183978
rect 345678 183922 345774 183978
rect 345154 166350 345774 183922
rect 348874 226350 349494 243922
rect 348874 226294 348970 226350
rect 349026 226294 349094 226350
rect 349150 226294 349218 226350
rect 349274 226294 349342 226350
rect 349398 226294 349494 226350
rect 348874 226226 349494 226294
rect 348874 226170 348970 226226
rect 349026 226170 349094 226226
rect 349150 226170 349218 226226
rect 349274 226170 349342 226226
rect 349398 226170 349494 226226
rect 348874 226102 349494 226170
rect 348874 226046 348970 226102
rect 349026 226046 349094 226102
rect 349150 226046 349218 226102
rect 349274 226046 349342 226102
rect 349398 226046 349494 226102
rect 348874 225978 349494 226046
rect 348874 225922 348970 225978
rect 349026 225922 349094 225978
rect 349150 225922 349218 225978
rect 349274 225922 349342 225978
rect 349398 225922 349494 225978
rect 348874 208350 349494 225922
rect 363154 597212 363774 598268
rect 363154 597156 363250 597212
rect 363306 597156 363374 597212
rect 363430 597156 363498 597212
rect 363554 597156 363622 597212
rect 363678 597156 363774 597212
rect 363154 597088 363774 597156
rect 363154 597032 363250 597088
rect 363306 597032 363374 597088
rect 363430 597032 363498 597088
rect 363554 597032 363622 597088
rect 363678 597032 363774 597088
rect 363154 596964 363774 597032
rect 363154 596908 363250 596964
rect 363306 596908 363374 596964
rect 363430 596908 363498 596964
rect 363554 596908 363622 596964
rect 363678 596908 363774 596964
rect 363154 596840 363774 596908
rect 363154 596784 363250 596840
rect 363306 596784 363374 596840
rect 363430 596784 363498 596840
rect 363554 596784 363622 596840
rect 363678 596784 363774 596840
rect 363154 580350 363774 596784
rect 363154 580294 363250 580350
rect 363306 580294 363374 580350
rect 363430 580294 363498 580350
rect 363554 580294 363622 580350
rect 363678 580294 363774 580350
rect 363154 580226 363774 580294
rect 363154 580170 363250 580226
rect 363306 580170 363374 580226
rect 363430 580170 363498 580226
rect 363554 580170 363622 580226
rect 363678 580170 363774 580226
rect 363154 580102 363774 580170
rect 363154 580046 363250 580102
rect 363306 580046 363374 580102
rect 363430 580046 363498 580102
rect 363554 580046 363622 580102
rect 363678 580046 363774 580102
rect 363154 579978 363774 580046
rect 363154 579922 363250 579978
rect 363306 579922 363374 579978
rect 363430 579922 363498 579978
rect 363554 579922 363622 579978
rect 363678 579922 363774 579978
rect 363154 562350 363774 579922
rect 363154 562294 363250 562350
rect 363306 562294 363374 562350
rect 363430 562294 363498 562350
rect 363554 562294 363622 562350
rect 363678 562294 363774 562350
rect 363154 562226 363774 562294
rect 363154 562170 363250 562226
rect 363306 562170 363374 562226
rect 363430 562170 363498 562226
rect 363554 562170 363622 562226
rect 363678 562170 363774 562226
rect 363154 562102 363774 562170
rect 363154 562046 363250 562102
rect 363306 562046 363374 562102
rect 363430 562046 363498 562102
rect 363554 562046 363622 562102
rect 363678 562046 363774 562102
rect 363154 561978 363774 562046
rect 363154 561922 363250 561978
rect 363306 561922 363374 561978
rect 363430 561922 363498 561978
rect 363554 561922 363622 561978
rect 363678 561922 363774 561978
rect 363154 544350 363774 561922
rect 363154 544294 363250 544350
rect 363306 544294 363374 544350
rect 363430 544294 363498 544350
rect 363554 544294 363622 544350
rect 363678 544294 363774 544350
rect 363154 544226 363774 544294
rect 363154 544170 363250 544226
rect 363306 544170 363374 544226
rect 363430 544170 363498 544226
rect 363554 544170 363622 544226
rect 363678 544170 363774 544226
rect 363154 544102 363774 544170
rect 363154 544046 363250 544102
rect 363306 544046 363374 544102
rect 363430 544046 363498 544102
rect 363554 544046 363622 544102
rect 363678 544046 363774 544102
rect 363154 543978 363774 544046
rect 363154 543922 363250 543978
rect 363306 543922 363374 543978
rect 363430 543922 363498 543978
rect 363554 543922 363622 543978
rect 363678 543922 363774 543978
rect 363154 526350 363774 543922
rect 363154 526294 363250 526350
rect 363306 526294 363374 526350
rect 363430 526294 363498 526350
rect 363554 526294 363622 526350
rect 363678 526294 363774 526350
rect 363154 526226 363774 526294
rect 363154 526170 363250 526226
rect 363306 526170 363374 526226
rect 363430 526170 363498 526226
rect 363554 526170 363622 526226
rect 363678 526170 363774 526226
rect 363154 526102 363774 526170
rect 363154 526046 363250 526102
rect 363306 526046 363374 526102
rect 363430 526046 363498 526102
rect 363554 526046 363622 526102
rect 363678 526046 363774 526102
rect 363154 525978 363774 526046
rect 363154 525922 363250 525978
rect 363306 525922 363374 525978
rect 363430 525922 363498 525978
rect 363554 525922 363622 525978
rect 363678 525922 363774 525978
rect 363154 508350 363774 525922
rect 363154 508294 363250 508350
rect 363306 508294 363374 508350
rect 363430 508294 363498 508350
rect 363554 508294 363622 508350
rect 363678 508294 363774 508350
rect 363154 508226 363774 508294
rect 363154 508170 363250 508226
rect 363306 508170 363374 508226
rect 363430 508170 363498 508226
rect 363554 508170 363622 508226
rect 363678 508170 363774 508226
rect 363154 508102 363774 508170
rect 363154 508046 363250 508102
rect 363306 508046 363374 508102
rect 363430 508046 363498 508102
rect 363554 508046 363622 508102
rect 363678 508046 363774 508102
rect 363154 507978 363774 508046
rect 363154 507922 363250 507978
rect 363306 507922 363374 507978
rect 363430 507922 363498 507978
rect 363554 507922 363622 507978
rect 363678 507922 363774 507978
rect 363154 490350 363774 507922
rect 363154 490294 363250 490350
rect 363306 490294 363374 490350
rect 363430 490294 363498 490350
rect 363554 490294 363622 490350
rect 363678 490294 363774 490350
rect 363154 490226 363774 490294
rect 363154 490170 363250 490226
rect 363306 490170 363374 490226
rect 363430 490170 363498 490226
rect 363554 490170 363622 490226
rect 363678 490170 363774 490226
rect 363154 490102 363774 490170
rect 363154 490046 363250 490102
rect 363306 490046 363374 490102
rect 363430 490046 363498 490102
rect 363554 490046 363622 490102
rect 363678 490046 363774 490102
rect 363154 489978 363774 490046
rect 363154 489922 363250 489978
rect 363306 489922 363374 489978
rect 363430 489922 363498 489978
rect 363554 489922 363622 489978
rect 363678 489922 363774 489978
rect 363154 472350 363774 489922
rect 363154 472294 363250 472350
rect 363306 472294 363374 472350
rect 363430 472294 363498 472350
rect 363554 472294 363622 472350
rect 363678 472294 363774 472350
rect 363154 472226 363774 472294
rect 363154 472170 363250 472226
rect 363306 472170 363374 472226
rect 363430 472170 363498 472226
rect 363554 472170 363622 472226
rect 363678 472170 363774 472226
rect 363154 472102 363774 472170
rect 363154 472046 363250 472102
rect 363306 472046 363374 472102
rect 363430 472046 363498 472102
rect 363554 472046 363622 472102
rect 363678 472046 363774 472102
rect 363154 471978 363774 472046
rect 363154 471922 363250 471978
rect 363306 471922 363374 471978
rect 363430 471922 363498 471978
rect 363554 471922 363622 471978
rect 363678 471922 363774 471978
rect 363154 454350 363774 471922
rect 363154 454294 363250 454350
rect 363306 454294 363374 454350
rect 363430 454294 363498 454350
rect 363554 454294 363622 454350
rect 363678 454294 363774 454350
rect 363154 454226 363774 454294
rect 363154 454170 363250 454226
rect 363306 454170 363374 454226
rect 363430 454170 363498 454226
rect 363554 454170 363622 454226
rect 363678 454170 363774 454226
rect 363154 454102 363774 454170
rect 363154 454046 363250 454102
rect 363306 454046 363374 454102
rect 363430 454046 363498 454102
rect 363554 454046 363622 454102
rect 363678 454046 363774 454102
rect 363154 453978 363774 454046
rect 363154 453922 363250 453978
rect 363306 453922 363374 453978
rect 363430 453922 363498 453978
rect 363554 453922 363622 453978
rect 363678 453922 363774 453978
rect 363154 436350 363774 453922
rect 363154 436294 363250 436350
rect 363306 436294 363374 436350
rect 363430 436294 363498 436350
rect 363554 436294 363622 436350
rect 363678 436294 363774 436350
rect 363154 436226 363774 436294
rect 363154 436170 363250 436226
rect 363306 436170 363374 436226
rect 363430 436170 363498 436226
rect 363554 436170 363622 436226
rect 363678 436170 363774 436226
rect 363154 436102 363774 436170
rect 363154 436046 363250 436102
rect 363306 436046 363374 436102
rect 363430 436046 363498 436102
rect 363554 436046 363622 436102
rect 363678 436046 363774 436102
rect 363154 435978 363774 436046
rect 363154 435922 363250 435978
rect 363306 435922 363374 435978
rect 363430 435922 363498 435978
rect 363554 435922 363622 435978
rect 363678 435922 363774 435978
rect 363154 418350 363774 435922
rect 363154 418294 363250 418350
rect 363306 418294 363374 418350
rect 363430 418294 363498 418350
rect 363554 418294 363622 418350
rect 363678 418294 363774 418350
rect 363154 418226 363774 418294
rect 363154 418170 363250 418226
rect 363306 418170 363374 418226
rect 363430 418170 363498 418226
rect 363554 418170 363622 418226
rect 363678 418170 363774 418226
rect 363154 418102 363774 418170
rect 363154 418046 363250 418102
rect 363306 418046 363374 418102
rect 363430 418046 363498 418102
rect 363554 418046 363622 418102
rect 363678 418046 363774 418102
rect 363154 417978 363774 418046
rect 363154 417922 363250 417978
rect 363306 417922 363374 417978
rect 363430 417922 363498 417978
rect 363554 417922 363622 417978
rect 363678 417922 363774 417978
rect 363154 400350 363774 417922
rect 363154 400294 363250 400350
rect 363306 400294 363374 400350
rect 363430 400294 363498 400350
rect 363554 400294 363622 400350
rect 363678 400294 363774 400350
rect 363154 400226 363774 400294
rect 363154 400170 363250 400226
rect 363306 400170 363374 400226
rect 363430 400170 363498 400226
rect 363554 400170 363622 400226
rect 363678 400170 363774 400226
rect 363154 400102 363774 400170
rect 363154 400046 363250 400102
rect 363306 400046 363374 400102
rect 363430 400046 363498 400102
rect 363554 400046 363622 400102
rect 363678 400046 363774 400102
rect 363154 399978 363774 400046
rect 363154 399922 363250 399978
rect 363306 399922 363374 399978
rect 363430 399922 363498 399978
rect 363554 399922 363622 399978
rect 363678 399922 363774 399978
rect 363154 382350 363774 399922
rect 363154 382294 363250 382350
rect 363306 382294 363374 382350
rect 363430 382294 363498 382350
rect 363554 382294 363622 382350
rect 363678 382294 363774 382350
rect 363154 382226 363774 382294
rect 363154 382170 363250 382226
rect 363306 382170 363374 382226
rect 363430 382170 363498 382226
rect 363554 382170 363622 382226
rect 363678 382170 363774 382226
rect 363154 382102 363774 382170
rect 363154 382046 363250 382102
rect 363306 382046 363374 382102
rect 363430 382046 363498 382102
rect 363554 382046 363622 382102
rect 363678 382046 363774 382102
rect 363154 381978 363774 382046
rect 363154 381922 363250 381978
rect 363306 381922 363374 381978
rect 363430 381922 363498 381978
rect 363554 381922 363622 381978
rect 363678 381922 363774 381978
rect 363154 364350 363774 381922
rect 363154 364294 363250 364350
rect 363306 364294 363374 364350
rect 363430 364294 363498 364350
rect 363554 364294 363622 364350
rect 363678 364294 363774 364350
rect 363154 364226 363774 364294
rect 363154 364170 363250 364226
rect 363306 364170 363374 364226
rect 363430 364170 363498 364226
rect 363554 364170 363622 364226
rect 363678 364170 363774 364226
rect 363154 364102 363774 364170
rect 363154 364046 363250 364102
rect 363306 364046 363374 364102
rect 363430 364046 363498 364102
rect 363554 364046 363622 364102
rect 363678 364046 363774 364102
rect 363154 363978 363774 364046
rect 363154 363922 363250 363978
rect 363306 363922 363374 363978
rect 363430 363922 363498 363978
rect 363554 363922 363622 363978
rect 363678 363922 363774 363978
rect 363154 346350 363774 363922
rect 363154 346294 363250 346350
rect 363306 346294 363374 346350
rect 363430 346294 363498 346350
rect 363554 346294 363622 346350
rect 363678 346294 363774 346350
rect 363154 346226 363774 346294
rect 363154 346170 363250 346226
rect 363306 346170 363374 346226
rect 363430 346170 363498 346226
rect 363554 346170 363622 346226
rect 363678 346170 363774 346226
rect 363154 346102 363774 346170
rect 363154 346046 363250 346102
rect 363306 346046 363374 346102
rect 363430 346046 363498 346102
rect 363554 346046 363622 346102
rect 363678 346046 363774 346102
rect 363154 345978 363774 346046
rect 363154 345922 363250 345978
rect 363306 345922 363374 345978
rect 363430 345922 363498 345978
rect 363554 345922 363622 345978
rect 363678 345922 363774 345978
rect 363154 328350 363774 345922
rect 363154 328294 363250 328350
rect 363306 328294 363374 328350
rect 363430 328294 363498 328350
rect 363554 328294 363622 328350
rect 363678 328294 363774 328350
rect 363154 328226 363774 328294
rect 363154 328170 363250 328226
rect 363306 328170 363374 328226
rect 363430 328170 363498 328226
rect 363554 328170 363622 328226
rect 363678 328170 363774 328226
rect 363154 328102 363774 328170
rect 363154 328046 363250 328102
rect 363306 328046 363374 328102
rect 363430 328046 363498 328102
rect 363554 328046 363622 328102
rect 363678 328046 363774 328102
rect 363154 327978 363774 328046
rect 363154 327922 363250 327978
rect 363306 327922 363374 327978
rect 363430 327922 363498 327978
rect 363554 327922 363622 327978
rect 363678 327922 363774 327978
rect 363154 310350 363774 327922
rect 363154 310294 363250 310350
rect 363306 310294 363374 310350
rect 363430 310294 363498 310350
rect 363554 310294 363622 310350
rect 363678 310294 363774 310350
rect 363154 310226 363774 310294
rect 363154 310170 363250 310226
rect 363306 310170 363374 310226
rect 363430 310170 363498 310226
rect 363554 310170 363622 310226
rect 363678 310170 363774 310226
rect 363154 310102 363774 310170
rect 363154 310046 363250 310102
rect 363306 310046 363374 310102
rect 363430 310046 363498 310102
rect 363554 310046 363622 310102
rect 363678 310046 363774 310102
rect 363154 309978 363774 310046
rect 363154 309922 363250 309978
rect 363306 309922 363374 309978
rect 363430 309922 363498 309978
rect 363554 309922 363622 309978
rect 363678 309922 363774 309978
rect 363154 292350 363774 309922
rect 363154 292294 363250 292350
rect 363306 292294 363374 292350
rect 363430 292294 363498 292350
rect 363554 292294 363622 292350
rect 363678 292294 363774 292350
rect 363154 292226 363774 292294
rect 363154 292170 363250 292226
rect 363306 292170 363374 292226
rect 363430 292170 363498 292226
rect 363554 292170 363622 292226
rect 363678 292170 363774 292226
rect 363154 292102 363774 292170
rect 363154 292046 363250 292102
rect 363306 292046 363374 292102
rect 363430 292046 363498 292102
rect 363554 292046 363622 292102
rect 363678 292046 363774 292102
rect 363154 291978 363774 292046
rect 363154 291922 363250 291978
rect 363306 291922 363374 291978
rect 363430 291922 363498 291978
rect 363554 291922 363622 291978
rect 363678 291922 363774 291978
rect 363154 274350 363774 291922
rect 363154 274294 363250 274350
rect 363306 274294 363374 274350
rect 363430 274294 363498 274350
rect 363554 274294 363622 274350
rect 363678 274294 363774 274350
rect 363154 274226 363774 274294
rect 363154 274170 363250 274226
rect 363306 274170 363374 274226
rect 363430 274170 363498 274226
rect 363554 274170 363622 274226
rect 363678 274170 363774 274226
rect 363154 274102 363774 274170
rect 363154 274046 363250 274102
rect 363306 274046 363374 274102
rect 363430 274046 363498 274102
rect 363554 274046 363622 274102
rect 363678 274046 363774 274102
rect 363154 273978 363774 274046
rect 363154 273922 363250 273978
rect 363306 273922 363374 273978
rect 363430 273922 363498 273978
rect 363554 273922 363622 273978
rect 363678 273922 363774 273978
rect 363154 256350 363774 273922
rect 363154 256294 363250 256350
rect 363306 256294 363374 256350
rect 363430 256294 363498 256350
rect 363554 256294 363622 256350
rect 363678 256294 363774 256350
rect 363154 256226 363774 256294
rect 363154 256170 363250 256226
rect 363306 256170 363374 256226
rect 363430 256170 363498 256226
rect 363554 256170 363622 256226
rect 363678 256170 363774 256226
rect 363154 256102 363774 256170
rect 363154 256046 363250 256102
rect 363306 256046 363374 256102
rect 363430 256046 363498 256102
rect 363554 256046 363622 256102
rect 363678 256046 363774 256102
rect 363154 255978 363774 256046
rect 363154 255922 363250 255978
rect 363306 255922 363374 255978
rect 363430 255922 363498 255978
rect 363554 255922 363622 255978
rect 363678 255922 363774 255978
rect 363154 238350 363774 255922
rect 363154 238294 363250 238350
rect 363306 238294 363374 238350
rect 363430 238294 363498 238350
rect 363554 238294 363622 238350
rect 363678 238294 363774 238350
rect 363154 238226 363774 238294
rect 363154 238170 363250 238226
rect 363306 238170 363374 238226
rect 363430 238170 363498 238226
rect 363554 238170 363622 238226
rect 363678 238170 363774 238226
rect 363154 238102 363774 238170
rect 363154 238046 363250 238102
rect 363306 238046 363374 238102
rect 363430 238046 363498 238102
rect 363554 238046 363622 238102
rect 363678 238046 363774 238102
rect 363154 237978 363774 238046
rect 363154 237922 363250 237978
rect 363306 237922 363374 237978
rect 363430 237922 363498 237978
rect 363554 237922 363622 237978
rect 363678 237922 363774 237978
rect 363154 220350 363774 237922
rect 363154 220294 363250 220350
rect 363306 220294 363374 220350
rect 363430 220294 363498 220350
rect 363554 220294 363622 220350
rect 363678 220294 363774 220350
rect 363154 220226 363774 220294
rect 363154 220170 363250 220226
rect 363306 220170 363374 220226
rect 363430 220170 363498 220226
rect 363554 220170 363622 220226
rect 363678 220170 363774 220226
rect 363154 220102 363774 220170
rect 363154 220046 363250 220102
rect 363306 220046 363374 220102
rect 363430 220046 363498 220102
rect 363554 220046 363622 220102
rect 363678 220046 363774 220102
rect 363154 219978 363774 220046
rect 363154 219922 363250 219978
rect 363306 219922 363374 219978
rect 363430 219922 363498 219978
rect 363554 219922 363622 219978
rect 363678 219922 363774 219978
rect 363154 217934 363774 219922
rect 366874 598172 367494 598268
rect 366874 598116 366970 598172
rect 367026 598116 367094 598172
rect 367150 598116 367218 598172
rect 367274 598116 367342 598172
rect 367398 598116 367494 598172
rect 366874 598048 367494 598116
rect 366874 597992 366970 598048
rect 367026 597992 367094 598048
rect 367150 597992 367218 598048
rect 367274 597992 367342 598048
rect 367398 597992 367494 598048
rect 366874 597924 367494 597992
rect 366874 597868 366970 597924
rect 367026 597868 367094 597924
rect 367150 597868 367218 597924
rect 367274 597868 367342 597924
rect 367398 597868 367494 597924
rect 366874 597800 367494 597868
rect 366874 597744 366970 597800
rect 367026 597744 367094 597800
rect 367150 597744 367218 597800
rect 367274 597744 367342 597800
rect 367398 597744 367494 597800
rect 366874 586350 367494 597744
rect 366874 586294 366970 586350
rect 367026 586294 367094 586350
rect 367150 586294 367218 586350
rect 367274 586294 367342 586350
rect 367398 586294 367494 586350
rect 366874 586226 367494 586294
rect 366874 586170 366970 586226
rect 367026 586170 367094 586226
rect 367150 586170 367218 586226
rect 367274 586170 367342 586226
rect 367398 586170 367494 586226
rect 366874 586102 367494 586170
rect 366874 586046 366970 586102
rect 367026 586046 367094 586102
rect 367150 586046 367218 586102
rect 367274 586046 367342 586102
rect 367398 586046 367494 586102
rect 366874 585978 367494 586046
rect 366874 585922 366970 585978
rect 367026 585922 367094 585978
rect 367150 585922 367218 585978
rect 367274 585922 367342 585978
rect 367398 585922 367494 585978
rect 366874 568350 367494 585922
rect 366874 568294 366970 568350
rect 367026 568294 367094 568350
rect 367150 568294 367218 568350
rect 367274 568294 367342 568350
rect 367398 568294 367494 568350
rect 366874 568226 367494 568294
rect 366874 568170 366970 568226
rect 367026 568170 367094 568226
rect 367150 568170 367218 568226
rect 367274 568170 367342 568226
rect 367398 568170 367494 568226
rect 366874 568102 367494 568170
rect 366874 568046 366970 568102
rect 367026 568046 367094 568102
rect 367150 568046 367218 568102
rect 367274 568046 367342 568102
rect 367398 568046 367494 568102
rect 366874 567978 367494 568046
rect 366874 567922 366970 567978
rect 367026 567922 367094 567978
rect 367150 567922 367218 567978
rect 367274 567922 367342 567978
rect 367398 567922 367494 567978
rect 366874 550350 367494 567922
rect 366874 550294 366970 550350
rect 367026 550294 367094 550350
rect 367150 550294 367218 550350
rect 367274 550294 367342 550350
rect 367398 550294 367494 550350
rect 366874 550226 367494 550294
rect 366874 550170 366970 550226
rect 367026 550170 367094 550226
rect 367150 550170 367218 550226
rect 367274 550170 367342 550226
rect 367398 550170 367494 550226
rect 366874 550102 367494 550170
rect 366874 550046 366970 550102
rect 367026 550046 367094 550102
rect 367150 550046 367218 550102
rect 367274 550046 367342 550102
rect 367398 550046 367494 550102
rect 366874 549978 367494 550046
rect 366874 549922 366970 549978
rect 367026 549922 367094 549978
rect 367150 549922 367218 549978
rect 367274 549922 367342 549978
rect 367398 549922 367494 549978
rect 366874 532350 367494 549922
rect 366874 532294 366970 532350
rect 367026 532294 367094 532350
rect 367150 532294 367218 532350
rect 367274 532294 367342 532350
rect 367398 532294 367494 532350
rect 366874 532226 367494 532294
rect 366874 532170 366970 532226
rect 367026 532170 367094 532226
rect 367150 532170 367218 532226
rect 367274 532170 367342 532226
rect 367398 532170 367494 532226
rect 366874 532102 367494 532170
rect 366874 532046 366970 532102
rect 367026 532046 367094 532102
rect 367150 532046 367218 532102
rect 367274 532046 367342 532102
rect 367398 532046 367494 532102
rect 366874 531978 367494 532046
rect 366874 531922 366970 531978
rect 367026 531922 367094 531978
rect 367150 531922 367218 531978
rect 367274 531922 367342 531978
rect 367398 531922 367494 531978
rect 366874 514350 367494 531922
rect 366874 514294 366970 514350
rect 367026 514294 367094 514350
rect 367150 514294 367218 514350
rect 367274 514294 367342 514350
rect 367398 514294 367494 514350
rect 366874 514226 367494 514294
rect 366874 514170 366970 514226
rect 367026 514170 367094 514226
rect 367150 514170 367218 514226
rect 367274 514170 367342 514226
rect 367398 514170 367494 514226
rect 366874 514102 367494 514170
rect 366874 514046 366970 514102
rect 367026 514046 367094 514102
rect 367150 514046 367218 514102
rect 367274 514046 367342 514102
rect 367398 514046 367494 514102
rect 366874 513978 367494 514046
rect 366874 513922 366970 513978
rect 367026 513922 367094 513978
rect 367150 513922 367218 513978
rect 367274 513922 367342 513978
rect 367398 513922 367494 513978
rect 366874 496350 367494 513922
rect 366874 496294 366970 496350
rect 367026 496294 367094 496350
rect 367150 496294 367218 496350
rect 367274 496294 367342 496350
rect 367398 496294 367494 496350
rect 366874 496226 367494 496294
rect 366874 496170 366970 496226
rect 367026 496170 367094 496226
rect 367150 496170 367218 496226
rect 367274 496170 367342 496226
rect 367398 496170 367494 496226
rect 366874 496102 367494 496170
rect 366874 496046 366970 496102
rect 367026 496046 367094 496102
rect 367150 496046 367218 496102
rect 367274 496046 367342 496102
rect 367398 496046 367494 496102
rect 366874 495978 367494 496046
rect 366874 495922 366970 495978
rect 367026 495922 367094 495978
rect 367150 495922 367218 495978
rect 367274 495922 367342 495978
rect 367398 495922 367494 495978
rect 366874 478350 367494 495922
rect 366874 478294 366970 478350
rect 367026 478294 367094 478350
rect 367150 478294 367218 478350
rect 367274 478294 367342 478350
rect 367398 478294 367494 478350
rect 366874 478226 367494 478294
rect 366874 478170 366970 478226
rect 367026 478170 367094 478226
rect 367150 478170 367218 478226
rect 367274 478170 367342 478226
rect 367398 478170 367494 478226
rect 366874 478102 367494 478170
rect 366874 478046 366970 478102
rect 367026 478046 367094 478102
rect 367150 478046 367218 478102
rect 367274 478046 367342 478102
rect 367398 478046 367494 478102
rect 366874 477978 367494 478046
rect 366874 477922 366970 477978
rect 367026 477922 367094 477978
rect 367150 477922 367218 477978
rect 367274 477922 367342 477978
rect 367398 477922 367494 477978
rect 366874 460350 367494 477922
rect 366874 460294 366970 460350
rect 367026 460294 367094 460350
rect 367150 460294 367218 460350
rect 367274 460294 367342 460350
rect 367398 460294 367494 460350
rect 366874 460226 367494 460294
rect 366874 460170 366970 460226
rect 367026 460170 367094 460226
rect 367150 460170 367218 460226
rect 367274 460170 367342 460226
rect 367398 460170 367494 460226
rect 366874 460102 367494 460170
rect 366874 460046 366970 460102
rect 367026 460046 367094 460102
rect 367150 460046 367218 460102
rect 367274 460046 367342 460102
rect 367398 460046 367494 460102
rect 366874 459978 367494 460046
rect 366874 459922 366970 459978
rect 367026 459922 367094 459978
rect 367150 459922 367218 459978
rect 367274 459922 367342 459978
rect 367398 459922 367494 459978
rect 366874 442350 367494 459922
rect 366874 442294 366970 442350
rect 367026 442294 367094 442350
rect 367150 442294 367218 442350
rect 367274 442294 367342 442350
rect 367398 442294 367494 442350
rect 366874 442226 367494 442294
rect 366874 442170 366970 442226
rect 367026 442170 367094 442226
rect 367150 442170 367218 442226
rect 367274 442170 367342 442226
rect 367398 442170 367494 442226
rect 366874 442102 367494 442170
rect 366874 442046 366970 442102
rect 367026 442046 367094 442102
rect 367150 442046 367218 442102
rect 367274 442046 367342 442102
rect 367398 442046 367494 442102
rect 366874 441978 367494 442046
rect 366874 441922 366970 441978
rect 367026 441922 367094 441978
rect 367150 441922 367218 441978
rect 367274 441922 367342 441978
rect 367398 441922 367494 441978
rect 366874 424350 367494 441922
rect 366874 424294 366970 424350
rect 367026 424294 367094 424350
rect 367150 424294 367218 424350
rect 367274 424294 367342 424350
rect 367398 424294 367494 424350
rect 366874 424226 367494 424294
rect 366874 424170 366970 424226
rect 367026 424170 367094 424226
rect 367150 424170 367218 424226
rect 367274 424170 367342 424226
rect 367398 424170 367494 424226
rect 366874 424102 367494 424170
rect 366874 424046 366970 424102
rect 367026 424046 367094 424102
rect 367150 424046 367218 424102
rect 367274 424046 367342 424102
rect 367398 424046 367494 424102
rect 366874 423978 367494 424046
rect 366874 423922 366970 423978
rect 367026 423922 367094 423978
rect 367150 423922 367218 423978
rect 367274 423922 367342 423978
rect 367398 423922 367494 423978
rect 366874 406350 367494 423922
rect 366874 406294 366970 406350
rect 367026 406294 367094 406350
rect 367150 406294 367218 406350
rect 367274 406294 367342 406350
rect 367398 406294 367494 406350
rect 366874 406226 367494 406294
rect 366874 406170 366970 406226
rect 367026 406170 367094 406226
rect 367150 406170 367218 406226
rect 367274 406170 367342 406226
rect 367398 406170 367494 406226
rect 366874 406102 367494 406170
rect 366874 406046 366970 406102
rect 367026 406046 367094 406102
rect 367150 406046 367218 406102
rect 367274 406046 367342 406102
rect 367398 406046 367494 406102
rect 366874 405978 367494 406046
rect 366874 405922 366970 405978
rect 367026 405922 367094 405978
rect 367150 405922 367218 405978
rect 367274 405922 367342 405978
rect 367398 405922 367494 405978
rect 366874 388350 367494 405922
rect 366874 388294 366970 388350
rect 367026 388294 367094 388350
rect 367150 388294 367218 388350
rect 367274 388294 367342 388350
rect 367398 388294 367494 388350
rect 366874 388226 367494 388294
rect 366874 388170 366970 388226
rect 367026 388170 367094 388226
rect 367150 388170 367218 388226
rect 367274 388170 367342 388226
rect 367398 388170 367494 388226
rect 366874 388102 367494 388170
rect 366874 388046 366970 388102
rect 367026 388046 367094 388102
rect 367150 388046 367218 388102
rect 367274 388046 367342 388102
rect 367398 388046 367494 388102
rect 366874 387978 367494 388046
rect 366874 387922 366970 387978
rect 367026 387922 367094 387978
rect 367150 387922 367218 387978
rect 367274 387922 367342 387978
rect 367398 387922 367494 387978
rect 366874 370350 367494 387922
rect 366874 370294 366970 370350
rect 367026 370294 367094 370350
rect 367150 370294 367218 370350
rect 367274 370294 367342 370350
rect 367398 370294 367494 370350
rect 366874 370226 367494 370294
rect 366874 370170 366970 370226
rect 367026 370170 367094 370226
rect 367150 370170 367218 370226
rect 367274 370170 367342 370226
rect 367398 370170 367494 370226
rect 366874 370102 367494 370170
rect 366874 370046 366970 370102
rect 367026 370046 367094 370102
rect 367150 370046 367218 370102
rect 367274 370046 367342 370102
rect 367398 370046 367494 370102
rect 366874 369978 367494 370046
rect 366874 369922 366970 369978
rect 367026 369922 367094 369978
rect 367150 369922 367218 369978
rect 367274 369922 367342 369978
rect 367398 369922 367494 369978
rect 366874 352350 367494 369922
rect 366874 352294 366970 352350
rect 367026 352294 367094 352350
rect 367150 352294 367218 352350
rect 367274 352294 367342 352350
rect 367398 352294 367494 352350
rect 366874 352226 367494 352294
rect 366874 352170 366970 352226
rect 367026 352170 367094 352226
rect 367150 352170 367218 352226
rect 367274 352170 367342 352226
rect 367398 352170 367494 352226
rect 366874 352102 367494 352170
rect 366874 352046 366970 352102
rect 367026 352046 367094 352102
rect 367150 352046 367218 352102
rect 367274 352046 367342 352102
rect 367398 352046 367494 352102
rect 366874 351978 367494 352046
rect 366874 351922 366970 351978
rect 367026 351922 367094 351978
rect 367150 351922 367218 351978
rect 367274 351922 367342 351978
rect 367398 351922 367494 351978
rect 366874 334350 367494 351922
rect 366874 334294 366970 334350
rect 367026 334294 367094 334350
rect 367150 334294 367218 334350
rect 367274 334294 367342 334350
rect 367398 334294 367494 334350
rect 366874 334226 367494 334294
rect 366874 334170 366970 334226
rect 367026 334170 367094 334226
rect 367150 334170 367218 334226
rect 367274 334170 367342 334226
rect 367398 334170 367494 334226
rect 366874 334102 367494 334170
rect 366874 334046 366970 334102
rect 367026 334046 367094 334102
rect 367150 334046 367218 334102
rect 367274 334046 367342 334102
rect 367398 334046 367494 334102
rect 366874 333978 367494 334046
rect 366874 333922 366970 333978
rect 367026 333922 367094 333978
rect 367150 333922 367218 333978
rect 367274 333922 367342 333978
rect 367398 333922 367494 333978
rect 366874 316350 367494 333922
rect 366874 316294 366970 316350
rect 367026 316294 367094 316350
rect 367150 316294 367218 316350
rect 367274 316294 367342 316350
rect 367398 316294 367494 316350
rect 366874 316226 367494 316294
rect 366874 316170 366970 316226
rect 367026 316170 367094 316226
rect 367150 316170 367218 316226
rect 367274 316170 367342 316226
rect 367398 316170 367494 316226
rect 366874 316102 367494 316170
rect 366874 316046 366970 316102
rect 367026 316046 367094 316102
rect 367150 316046 367218 316102
rect 367274 316046 367342 316102
rect 367398 316046 367494 316102
rect 366874 315978 367494 316046
rect 366874 315922 366970 315978
rect 367026 315922 367094 315978
rect 367150 315922 367218 315978
rect 367274 315922 367342 315978
rect 367398 315922 367494 315978
rect 366874 298350 367494 315922
rect 366874 298294 366970 298350
rect 367026 298294 367094 298350
rect 367150 298294 367218 298350
rect 367274 298294 367342 298350
rect 367398 298294 367494 298350
rect 366874 298226 367494 298294
rect 366874 298170 366970 298226
rect 367026 298170 367094 298226
rect 367150 298170 367218 298226
rect 367274 298170 367342 298226
rect 367398 298170 367494 298226
rect 366874 298102 367494 298170
rect 366874 298046 366970 298102
rect 367026 298046 367094 298102
rect 367150 298046 367218 298102
rect 367274 298046 367342 298102
rect 367398 298046 367494 298102
rect 366874 297978 367494 298046
rect 366874 297922 366970 297978
rect 367026 297922 367094 297978
rect 367150 297922 367218 297978
rect 367274 297922 367342 297978
rect 367398 297922 367494 297978
rect 366874 280350 367494 297922
rect 366874 280294 366970 280350
rect 367026 280294 367094 280350
rect 367150 280294 367218 280350
rect 367274 280294 367342 280350
rect 367398 280294 367494 280350
rect 366874 280226 367494 280294
rect 366874 280170 366970 280226
rect 367026 280170 367094 280226
rect 367150 280170 367218 280226
rect 367274 280170 367342 280226
rect 367398 280170 367494 280226
rect 366874 280102 367494 280170
rect 366874 280046 366970 280102
rect 367026 280046 367094 280102
rect 367150 280046 367218 280102
rect 367274 280046 367342 280102
rect 367398 280046 367494 280102
rect 366874 279978 367494 280046
rect 366874 279922 366970 279978
rect 367026 279922 367094 279978
rect 367150 279922 367218 279978
rect 367274 279922 367342 279978
rect 367398 279922 367494 279978
rect 366874 262350 367494 279922
rect 366874 262294 366970 262350
rect 367026 262294 367094 262350
rect 367150 262294 367218 262350
rect 367274 262294 367342 262350
rect 367398 262294 367494 262350
rect 366874 262226 367494 262294
rect 366874 262170 366970 262226
rect 367026 262170 367094 262226
rect 367150 262170 367218 262226
rect 367274 262170 367342 262226
rect 367398 262170 367494 262226
rect 366874 262102 367494 262170
rect 366874 262046 366970 262102
rect 367026 262046 367094 262102
rect 367150 262046 367218 262102
rect 367274 262046 367342 262102
rect 367398 262046 367494 262102
rect 366874 261978 367494 262046
rect 366874 261922 366970 261978
rect 367026 261922 367094 261978
rect 367150 261922 367218 261978
rect 367274 261922 367342 261978
rect 367398 261922 367494 261978
rect 366874 244350 367494 261922
rect 366874 244294 366970 244350
rect 367026 244294 367094 244350
rect 367150 244294 367218 244350
rect 367274 244294 367342 244350
rect 367398 244294 367494 244350
rect 366874 244226 367494 244294
rect 366874 244170 366970 244226
rect 367026 244170 367094 244226
rect 367150 244170 367218 244226
rect 367274 244170 367342 244226
rect 367398 244170 367494 244226
rect 366874 244102 367494 244170
rect 366874 244046 366970 244102
rect 367026 244046 367094 244102
rect 367150 244046 367218 244102
rect 367274 244046 367342 244102
rect 367398 244046 367494 244102
rect 366874 243978 367494 244046
rect 366874 243922 366970 243978
rect 367026 243922 367094 243978
rect 367150 243922 367218 243978
rect 367274 243922 367342 243978
rect 367398 243922 367494 243978
rect 366874 226350 367494 243922
rect 366874 226294 366970 226350
rect 367026 226294 367094 226350
rect 367150 226294 367218 226350
rect 367274 226294 367342 226350
rect 367398 226294 367494 226350
rect 366874 226226 367494 226294
rect 366874 226170 366970 226226
rect 367026 226170 367094 226226
rect 367150 226170 367218 226226
rect 367274 226170 367342 226226
rect 367398 226170 367494 226226
rect 366874 226102 367494 226170
rect 366874 226046 366970 226102
rect 367026 226046 367094 226102
rect 367150 226046 367218 226102
rect 367274 226046 367342 226102
rect 367398 226046 367494 226102
rect 366874 225978 367494 226046
rect 366874 225922 366970 225978
rect 367026 225922 367094 225978
rect 367150 225922 367218 225978
rect 367274 225922 367342 225978
rect 367398 225922 367494 225978
rect 366874 217934 367494 225922
rect 381154 597212 381774 598268
rect 381154 597156 381250 597212
rect 381306 597156 381374 597212
rect 381430 597156 381498 597212
rect 381554 597156 381622 597212
rect 381678 597156 381774 597212
rect 381154 597088 381774 597156
rect 381154 597032 381250 597088
rect 381306 597032 381374 597088
rect 381430 597032 381498 597088
rect 381554 597032 381622 597088
rect 381678 597032 381774 597088
rect 381154 596964 381774 597032
rect 381154 596908 381250 596964
rect 381306 596908 381374 596964
rect 381430 596908 381498 596964
rect 381554 596908 381622 596964
rect 381678 596908 381774 596964
rect 381154 596840 381774 596908
rect 381154 596784 381250 596840
rect 381306 596784 381374 596840
rect 381430 596784 381498 596840
rect 381554 596784 381622 596840
rect 381678 596784 381774 596840
rect 381154 580350 381774 596784
rect 381154 580294 381250 580350
rect 381306 580294 381374 580350
rect 381430 580294 381498 580350
rect 381554 580294 381622 580350
rect 381678 580294 381774 580350
rect 381154 580226 381774 580294
rect 381154 580170 381250 580226
rect 381306 580170 381374 580226
rect 381430 580170 381498 580226
rect 381554 580170 381622 580226
rect 381678 580170 381774 580226
rect 381154 580102 381774 580170
rect 381154 580046 381250 580102
rect 381306 580046 381374 580102
rect 381430 580046 381498 580102
rect 381554 580046 381622 580102
rect 381678 580046 381774 580102
rect 381154 579978 381774 580046
rect 381154 579922 381250 579978
rect 381306 579922 381374 579978
rect 381430 579922 381498 579978
rect 381554 579922 381622 579978
rect 381678 579922 381774 579978
rect 381154 562350 381774 579922
rect 381154 562294 381250 562350
rect 381306 562294 381374 562350
rect 381430 562294 381498 562350
rect 381554 562294 381622 562350
rect 381678 562294 381774 562350
rect 381154 562226 381774 562294
rect 381154 562170 381250 562226
rect 381306 562170 381374 562226
rect 381430 562170 381498 562226
rect 381554 562170 381622 562226
rect 381678 562170 381774 562226
rect 381154 562102 381774 562170
rect 381154 562046 381250 562102
rect 381306 562046 381374 562102
rect 381430 562046 381498 562102
rect 381554 562046 381622 562102
rect 381678 562046 381774 562102
rect 381154 561978 381774 562046
rect 381154 561922 381250 561978
rect 381306 561922 381374 561978
rect 381430 561922 381498 561978
rect 381554 561922 381622 561978
rect 381678 561922 381774 561978
rect 381154 544350 381774 561922
rect 381154 544294 381250 544350
rect 381306 544294 381374 544350
rect 381430 544294 381498 544350
rect 381554 544294 381622 544350
rect 381678 544294 381774 544350
rect 381154 544226 381774 544294
rect 381154 544170 381250 544226
rect 381306 544170 381374 544226
rect 381430 544170 381498 544226
rect 381554 544170 381622 544226
rect 381678 544170 381774 544226
rect 381154 544102 381774 544170
rect 381154 544046 381250 544102
rect 381306 544046 381374 544102
rect 381430 544046 381498 544102
rect 381554 544046 381622 544102
rect 381678 544046 381774 544102
rect 381154 543978 381774 544046
rect 381154 543922 381250 543978
rect 381306 543922 381374 543978
rect 381430 543922 381498 543978
rect 381554 543922 381622 543978
rect 381678 543922 381774 543978
rect 381154 526350 381774 543922
rect 381154 526294 381250 526350
rect 381306 526294 381374 526350
rect 381430 526294 381498 526350
rect 381554 526294 381622 526350
rect 381678 526294 381774 526350
rect 381154 526226 381774 526294
rect 381154 526170 381250 526226
rect 381306 526170 381374 526226
rect 381430 526170 381498 526226
rect 381554 526170 381622 526226
rect 381678 526170 381774 526226
rect 381154 526102 381774 526170
rect 381154 526046 381250 526102
rect 381306 526046 381374 526102
rect 381430 526046 381498 526102
rect 381554 526046 381622 526102
rect 381678 526046 381774 526102
rect 381154 525978 381774 526046
rect 381154 525922 381250 525978
rect 381306 525922 381374 525978
rect 381430 525922 381498 525978
rect 381554 525922 381622 525978
rect 381678 525922 381774 525978
rect 381154 508350 381774 525922
rect 381154 508294 381250 508350
rect 381306 508294 381374 508350
rect 381430 508294 381498 508350
rect 381554 508294 381622 508350
rect 381678 508294 381774 508350
rect 381154 508226 381774 508294
rect 381154 508170 381250 508226
rect 381306 508170 381374 508226
rect 381430 508170 381498 508226
rect 381554 508170 381622 508226
rect 381678 508170 381774 508226
rect 381154 508102 381774 508170
rect 381154 508046 381250 508102
rect 381306 508046 381374 508102
rect 381430 508046 381498 508102
rect 381554 508046 381622 508102
rect 381678 508046 381774 508102
rect 381154 507978 381774 508046
rect 381154 507922 381250 507978
rect 381306 507922 381374 507978
rect 381430 507922 381498 507978
rect 381554 507922 381622 507978
rect 381678 507922 381774 507978
rect 381154 490350 381774 507922
rect 381154 490294 381250 490350
rect 381306 490294 381374 490350
rect 381430 490294 381498 490350
rect 381554 490294 381622 490350
rect 381678 490294 381774 490350
rect 381154 490226 381774 490294
rect 381154 490170 381250 490226
rect 381306 490170 381374 490226
rect 381430 490170 381498 490226
rect 381554 490170 381622 490226
rect 381678 490170 381774 490226
rect 381154 490102 381774 490170
rect 381154 490046 381250 490102
rect 381306 490046 381374 490102
rect 381430 490046 381498 490102
rect 381554 490046 381622 490102
rect 381678 490046 381774 490102
rect 381154 489978 381774 490046
rect 381154 489922 381250 489978
rect 381306 489922 381374 489978
rect 381430 489922 381498 489978
rect 381554 489922 381622 489978
rect 381678 489922 381774 489978
rect 381154 472350 381774 489922
rect 381154 472294 381250 472350
rect 381306 472294 381374 472350
rect 381430 472294 381498 472350
rect 381554 472294 381622 472350
rect 381678 472294 381774 472350
rect 381154 472226 381774 472294
rect 381154 472170 381250 472226
rect 381306 472170 381374 472226
rect 381430 472170 381498 472226
rect 381554 472170 381622 472226
rect 381678 472170 381774 472226
rect 381154 472102 381774 472170
rect 381154 472046 381250 472102
rect 381306 472046 381374 472102
rect 381430 472046 381498 472102
rect 381554 472046 381622 472102
rect 381678 472046 381774 472102
rect 381154 471978 381774 472046
rect 381154 471922 381250 471978
rect 381306 471922 381374 471978
rect 381430 471922 381498 471978
rect 381554 471922 381622 471978
rect 381678 471922 381774 471978
rect 381154 454350 381774 471922
rect 381154 454294 381250 454350
rect 381306 454294 381374 454350
rect 381430 454294 381498 454350
rect 381554 454294 381622 454350
rect 381678 454294 381774 454350
rect 381154 454226 381774 454294
rect 381154 454170 381250 454226
rect 381306 454170 381374 454226
rect 381430 454170 381498 454226
rect 381554 454170 381622 454226
rect 381678 454170 381774 454226
rect 381154 454102 381774 454170
rect 381154 454046 381250 454102
rect 381306 454046 381374 454102
rect 381430 454046 381498 454102
rect 381554 454046 381622 454102
rect 381678 454046 381774 454102
rect 381154 453978 381774 454046
rect 381154 453922 381250 453978
rect 381306 453922 381374 453978
rect 381430 453922 381498 453978
rect 381554 453922 381622 453978
rect 381678 453922 381774 453978
rect 381154 436350 381774 453922
rect 381154 436294 381250 436350
rect 381306 436294 381374 436350
rect 381430 436294 381498 436350
rect 381554 436294 381622 436350
rect 381678 436294 381774 436350
rect 381154 436226 381774 436294
rect 381154 436170 381250 436226
rect 381306 436170 381374 436226
rect 381430 436170 381498 436226
rect 381554 436170 381622 436226
rect 381678 436170 381774 436226
rect 381154 436102 381774 436170
rect 381154 436046 381250 436102
rect 381306 436046 381374 436102
rect 381430 436046 381498 436102
rect 381554 436046 381622 436102
rect 381678 436046 381774 436102
rect 381154 435978 381774 436046
rect 381154 435922 381250 435978
rect 381306 435922 381374 435978
rect 381430 435922 381498 435978
rect 381554 435922 381622 435978
rect 381678 435922 381774 435978
rect 381154 418350 381774 435922
rect 381154 418294 381250 418350
rect 381306 418294 381374 418350
rect 381430 418294 381498 418350
rect 381554 418294 381622 418350
rect 381678 418294 381774 418350
rect 381154 418226 381774 418294
rect 381154 418170 381250 418226
rect 381306 418170 381374 418226
rect 381430 418170 381498 418226
rect 381554 418170 381622 418226
rect 381678 418170 381774 418226
rect 381154 418102 381774 418170
rect 381154 418046 381250 418102
rect 381306 418046 381374 418102
rect 381430 418046 381498 418102
rect 381554 418046 381622 418102
rect 381678 418046 381774 418102
rect 381154 417978 381774 418046
rect 381154 417922 381250 417978
rect 381306 417922 381374 417978
rect 381430 417922 381498 417978
rect 381554 417922 381622 417978
rect 381678 417922 381774 417978
rect 381154 400350 381774 417922
rect 381154 400294 381250 400350
rect 381306 400294 381374 400350
rect 381430 400294 381498 400350
rect 381554 400294 381622 400350
rect 381678 400294 381774 400350
rect 381154 400226 381774 400294
rect 381154 400170 381250 400226
rect 381306 400170 381374 400226
rect 381430 400170 381498 400226
rect 381554 400170 381622 400226
rect 381678 400170 381774 400226
rect 381154 400102 381774 400170
rect 381154 400046 381250 400102
rect 381306 400046 381374 400102
rect 381430 400046 381498 400102
rect 381554 400046 381622 400102
rect 381678 400046 381774 400102
rect 381154 399978 381774 400046
rect 381154 399922 381250 399978
rect 381306 399922 381374 399978
rect 381430 399922 381498 399978
rect 381554 399922 381622 399978
rect 381678 399922 381774 399978
rect 381154 382350 381774 399922
rect 381154 382294 381250 382350
rect 381306 382294 381374 382350
rect 381430 382294 381498 382350
rect 381554 382294 381622 382350
rect 381678 382294 381774 382350
rect 381154 382226 381774 382294
rect 381154 382170 381250 382226
rect 381306 382170 381374 382226
rect 381430 382170 381498 382226
rect 381554 382170 381622 382226
rect 381678 382170 381774 382226
rect 381154 382102 381774 382170
rect 381154 382046 381250 382102
rect 381306 382046 381374 382102
rect 381430 382046 381498 382102
rect 381554 382046 381622 382102
rect 381678 382046 381774 382102
rect 381154 381978 381774 382046
rect 381154 381922 381250 381978
rect 381306 381922 381374 381978
rect 381430 381922 381498 381978
rect 381554 381922 381622 381978
rect 381678 381922 381774 381978
rect 381154 364350 381774 381922
rect 381154 364294 381250 364350
rect 381306 364294 381374 364350
rect 381430 364294 381498 364350
rect 381554 364294 381622 364350
rect 381678 364294 381774 364350
rect 381154 364226 381774 364294
rect 381154 364170 381250 364226
rect 381306 364170 381374 364226
rect 381430 364170 381498 364226
rect 381554 364170 381622 364226
rect 381678 364170 381774 364226
rect 381154 364102 381774 364170
rect 381154 364046 381250 364102
rect 381306 364046 381374 364102
rect 381430 364046 381498 364102
rect 381554 364046 381622 364102
rect 381678 364046 381774 364102
rect 381154 363978 381774 364046
rect 381154 363922 381250 363978
rect 381306 363922 381374 363978
rect 381430 363922 381498 363978
rect 381554 363922 381622 363978
rect 381678 363922 381774 363978
rect 381154 346350 381774 363922
rect 381154 346294 381250 346350
rect 381306 346294 381374 346350
rect 381430 346294 381498 346350
rect 381554 346294 381622 346350
rect 381678 346294 381774 346350
rect 381154 346226 381774 346294
rect 381154 346170 381250 346226
rect 381306 346170 381374 346226
rect 381430 346170 381498 346226
rect 381554 346170 381622 346226
rect 381678 346170 381774 346226
rect 381154 346102 381774 346170
rect 381154 346046 381250 346102
rect 381306 346046 381374 346102
rect 381430 346046 381498 346102
rect 381554 346046 381622 346102
rect 381678 346046 381774 346102
rect 381154 345978 381774 346046
rect 381154 345922 381250 345978
rect 381306 345922 381374 345978
rect 381430 345922 381498 345978
rect 381554 345922 381622 345978
rect 381678 345922 381774 345978
rect 381154 328350 381774 345922
rect 381154 328294 381250 328350
rect 381306 328294 381374 328350
rect 381430 328294 381498 328350
rect 381554 328294 381622 328350
rect 381678 328294 381774 328350
rect 381154 328226 381774 328294
rect 381154 328170 381250 328226
rect 381306 328170 381374 328226
rect 381430 328170 381498 328226
rect 381554 328170 381622 328226
rect 381678 328170 381774 328226
rect 381154 328102 381774 328170
rect 381154 328046 381250 328102
rect 381306 328046 381374 328102
rect 381430 328046 381498 328102
rect 381554 328046 381622 328102
rect 381678 328046 381774 328102
rect 381154 327978 381774 328046
rect 381154 327922 381250 327978
rect 381306 327922 381374 327978
rect 381430 327922 381498 327978
rect 381554 327922 381622 327978
rect 381678 327922 381774 327978
rect 381154 310350 381774 327922
rect 381154 310294 381250 310350
rect 381306 310294 381374 310350
rect 381430 310294 381498 310350
rect 381554 310294 381622 310350
rect 381678 310294 381774 310350
rect 381154 310226 381774 310294
rect 381154 310170 381250 310226
rect 381306 310170 381374 310226
rect 381430 310170 381498 310226
rect 381554 310170 381622 310226
rect 381678 310170 381774 310226
rect 381154 310102 381774 310170
rect 381154 310046 381250 310102
rect 381306 310046 381374 310102
rect 381430 310046 381498 310102
rect 381554 310046 381622 310102
rect 381678 310046 381774 310102
rect 381154 309978 381774 310046
rect 381154 309922 381250 309978
rect 381306 309922 381374 309978
rect 381430 309922 381498 309978
rect 381554 309922 381622 309978
rect 381678 309922 381774 309978
rect 381154 292350 381774 309922
rect 381154 292294 381250 292350
rect 381306 292294 381374 292350
rect 381430 292294 381498 292350
rect 381554 292294 381622 292350
rect 381678 292294 381774 292350
rect 381154 292226 381774 292294
rect 381154 292170 381250 292226
rect 381306 292170 381374 292226
rect 381430 292170 381498 292226
rect 381554 292170 381622 292226
rect 381678 292170 381774 292226
rect 381154 292102 381774 292170
rect 381154 292046 381250 292102
rect 381306 292046 381374 292102
rect 381430 292046 381498 292102
rect 381554 292046 381622 292102
rect 381678 292046 381774 292102
rect 381154 291978 381774 292046
rect 381154 291922 381250 291978
rect 381306 291922 381374 291978
rect 381430 291922 381498 291978
rect 381554 291922 381622 291978
rect 381678 291922 381774 291978
rect 381154 274350 381774 291922
rect 381154 274294 381250 274350
rect 381306 274294 381374 274350
rect 381430 274294 381498 274350
rect 381554 274294 381622 274350
rect 381678 274294 381774 274350
rect 381154 274226 381774 274294
rect 381154 274170 381250 274226
rect 381306 274170 381374 274226
rect 381430 274170 381498 274226
rect 381554 274170 381622 274226
rect 381678 274170 381774 274226
rect 381154 274102 381774 274170
rect 381154 274046 381250 274102
rect 381306 274046 381374 274102
rect 381430 274046 381498 274102
rect 381554 274046 381622 274102
rect 381678 274046 381774 274102
rect 381154 273978 381774 274046
rect 381154 273922 381250 273978
rect 381306 273922 381374 273978
rect 381430 273922 381498 273978
rect 381554 273922 381622 273978
rect 381678 273922 381774 273978
rect 381154 256350 381774 273922
rect 381154 256294 381250 256350
rect 381306 256294 381374 256350
rect 381430 256294 381498 256350
rect 381554 256294 381622 256350
rect 381678 256294 381774 256350
rect 381154 256226 381774 256294
rect 381154 256170 381250 256226
rect 381306 256170 381374 256226
rect 381430 256170 381498 256226
rect 381554 256170 381622 256226
rect 381678 256170 381774 256226
rect 381154 256102 381774 256170
rect 381154 256046 381250 256102
rect 381306 256046 381374 256102
rect 381430 256046 381498 256102
rect 381554 256046 381622 256102
rect 381678 256046 381774 256102
rect 381154 255978 381774 256046
rect 381154 255922 381250 255978
rect 381306 255922 381374 255978
rect 381430 255922 381498 255978
rect 381554 255922 381622 255978
rect 381678 255922 381774 255978
rect 381154 238350 381774 255922
rect 381154 238294 381250 238350
rect 381306 238294 381374 238350
rect 381430 238294 381498 238350
rect 381554 238294 381622 238350
rect 381678 238294 381774 238350
rect 381154 238226 381774 238294
rect 381154 238170 381250 238226
rect 381306 238170 381374 238226
rect 381430 238170 381498 238226
rect 381554 238170 381622 238226
rect 381678 238170 381774 238226
rect 381154 238102 381774 238170
rect 381154 238046 381250 238102
rect 381306 238046 381374 238102
rect 381430 238046 381498 238102
rect 381554 238046 381622 238102
rect 381678 238046 381774 238102
rect 381154 237978 381774 238046
rect 381154 237922 381250 237978
rect 381306 237922 381374 237978
rect 381430 237922 381498 237978
rect 381554 237922 381622 237978
rect 381678 237922 381774 237978
rect 381154 220350 381774 237922
rect 381154 220294 381250 220350
rect 381306 220294 381374 220350
rect 381430 220294 381498 220350
rect 381554 220294 381622 220350
rect 381678 220294 381774 220350
rect 381154 220226 381774 220294
rect 381154 220170 381250 220226
rect 381306 220170 381374 220226
rect 381430 220170 381498 220226
rect 381554 220170 381622 220226
rect 381678 220170 381774 220226
rect 381154 220102 381774 220170
rect 381154 220046 381250 220102
rect 381306 220046 381374 220102
rect 381430 220046 381498 220102
rect 381554 220046 381622 220102
rect 381678 220046 381774 220102
rect 381154 219978 381774 220046
rect 381154 219922 381250 219978
rect 381306 219922 381374 219978
rect 381430 219922 381498 219978
rect 381554 219922 381622 219978
rect 381678 219922 381774 219978
rect 381154 217934 381774 219922
rect 399154 597212 399774 598268
rect 399154 597156 399250 597212
rect 399306 597156 399374 597212
rect 399430 597156 399498 597212
rect 399554 597156 399622 597212
rect 399678 597156 399774 597212
rect 399154 597088 399774 597156
rect 399154 597032 399250 597088
rect 399306 597032 399374 597088
rect 399430 597032 399498 597088
rect 399554 597032 399622 597088
rect 399678 597032 399774 597088
rect 399154 596964 399774 597032
rect 399154 596908 399250 596964
rect 399306 596908 399374 596964
rect 399430 596908 399498 596964
rect 399554 596908 399622 596964
rect 399678 596908 399774 596964
rect 399154 596840 399774 596908
rect 399154 596784 399250 596840
rect 399306 596784 399374 596840
rect 399430 596784 399498 596840
rect 399554 596784 399622 596840
rect 399678 596784 399774 596840
rect 399154 580350 399774 596784
rect 399154 580294 399250 580350
rect 399306 580294 399374 580350
rect 399430 580294 399498 580350
rect 399554 580294 399622 580350
rect 399678 580294 399774 580350
rect 399154 580226 399774 580294
rect 399154 580170 399250 580226
rect 399306 580170 399374 580226
rect 399430 580170 399498 580226
rect 399554 580170 399622 580226
rect 399678 580170 399774 580226
rect 399154 580102 399774 580170
rect 399154 580046 399250 580102
rect 399306 580046 399374 580102
rect 399430 580046 399498 580102
rect 399554 580046 399622 580102
rect 399678 580046 399774 580102
rect 399154 579978 399774 580046
rect 399154 579922 399250 579978
rect 399306 579922 399374 579978
rect 399430 579922 399498 579978
rect 399554 579922 399622 579978
rect 399678 579922 399774 579978
rect 399154 562350 399774 579922
rect 399154 562294 399250 562350
rect 399306 562294 399374 562350
rect 399430 562294 399498 562350
rect 399554 562294 399622 562350
rect 399678 562294 399774 562350
rect 399154 562226 399774 562294
rect 399154 562170 399250 562226
rect 399306 562170 399374 562226
rect 399430 562170 399498 562226
rect 399554 562170 399622 562226
rect 399678 562170 399774 562226
rect 399154 562102 399774 562170
rect 399154 562046 399250 562102
rect 399306 562046 399374 562102
rect 399430 562046 399498 562102
rect 399554 562046 399622 562102
rect 399678 562046 399774 562102
rect 399154 561978 399774 562046
rect 399154 561922 399250 561978
rect 399306 561922 399374 561978
rect 399430 561922 399498 561978
rect 399554 561922 399622 561978
rect 399678 561922 399774 561978
rect 399154 544350 399774 561922
rect 399154 544294 399250 544350
rect 399306 544294 399374 544350
rect 399430 544294 399498 544350
rect 399554 544294 399622 544350
rect 399678 544294 399774 544350
rect 399154 544226 399774 544294
rect 399154 544170 399250 544226
rect 399306 544170 399374 544226
rect 399430 544170 399498 544226
rect 399554 544170 399622 544226
rect 399678 544170 399774 544226
rect 399154 544102 399774 544170
rect 399154 544046 399250 544102
rect 399306 544046 399374 544102
rect 399430 544046 399498 544102
rect 399554 544046 399622 544102
rect 399678 544046 399774 544102
rect 399154 543978 399774 544046
rect 399154 543922 399250 543978
rect 399306 543922 399374 543978
rect 399430 543922 399498 543978
rect 399554 543922 399622 543978
rect 399678 543922 399774 543978
rect 399154 526350 399774 543922
rect 399154 526294 399250 526350
rect 399306 526294 399374 526350
rect 399430 526294 399498 526350
rect 399554 526294 399622 526350
rect 399678 526294 399774 526350
rect 399154 526226 399774 526294
rect 399154 526170 399250 526226
rect 399306 526170 399374 526226
rect 399430 526170 399498 526226
rect 399554 526170 399622 526226
rect 399678 526170 399774 526226
rect 399154 526102 399774 526170
rect 399154 526046 399250 526102
rect 399306 526046 399374 526102
rect 399430 526046 399498 526102
rect 399554 526046 399622 526102
rect 399678 526046 399774 526102
rect 399154 525978 399774 526046
rect 399154 525922 399250 525978
rect 399306 525922 399374 525978
rect 399430 525922 399498 525978
rect 399554 525922 399622 525978
rect 399678 525922 399774 525978
rect 399154 508350 399774 525922
rect 399154 508294 399250 508350
rect 399306 508294 399374 508350
rect 399430 508294 399498 508350
rect 399554 508294 399622 508350
rect 399678 508294 399774 508350
rect 399154 508226 399774 508294
rect 399154 508170 399250 508226
rect 399306 508170 399374 508226
rect 399430 508170 399498 508226
rect 399554 508170 399622 508226
rect 399678 508170 399774 508226
rect 399154 508102 399774 508170
rect 399154 508046 399250 508102
rect 399306 508046 399374 508102
rect 399430 508046 399498 508102
rect 399554 508046 399622 508102
rect 399678 508046 399774 508102
rect 399154 507978 399774 508046
rect 399154 507922 399250 507978
rect 399306 507922 399374 507978
rect 399430 507922 399498 507978
rect 399554 507922 399622 507978
rect 399678 507922 399774 507978
rect 399154 490350 399774 507922
rect 399154 490294 399250 490350
rect 399306 490294 399374 490350
rect 399430 490294 399498 490350
rect 399554 490294 399622 490350
rect 399678 490294 399774 490350
rect 399154 490226 399774 490294
rect 399154 490170 399250 490226
rect 399306 490170 399374 490226
rect 399430 490170 399498 490226
rect 399554 490170 399622 490226
rect 399678 490170 399774 490226
rect 399154 490102 399774 490170
rect 399154 490046 399250 490102
rect 399306 490046 399374 490102
rect 399430 490046 399498 490102
rect 399554 490046 399622 490102
rect 399678 490046 399774 490102
rect 399154 489978 399774 490046
rect 399154 489922 399250 489978
rect 399306 489922 399374 489978
rect 399430 489922 399498 489978
rect 399554 489922 399622 489978
rect 399678 489922 399774 489978
rect 399154 472350 399774 489922
rect 399154 472294 399250 472350
rect 399306 472294 399374 472350
rect 399430 472294 399498 472350
rect 399554 472294 399622 472350
rect 399678 472294 399774 472350
rect 399154 472226 399774 472294
rect 399154 472170 399250 472226
rect 399306 472170 399374 472226
rect 399430 472170 399498 472226
rect 399554 472170 399622 472226
rect 399678 472170 399774 472226
rect 399154 472102 399774 472170
rect 399154 472046 399250 472102
rect 399306 472046 399374 472102
rect 399430 472046 399498 472102
rect 399554 472046 399622 472102
rect 399678 472046 399774 472102
rect 399154 471978 399774 472046
rect 399154 471922 399250 471978
rect 399306 471922 399374 471978
rect 399430 471922 399498 471978
rect 399554 471922 399622 471978
rect 399678 471922 399774 471978
rect 399154 454350 399774 471922
rect 399154 454294 399250 454350
rect 399306 454294 399374 454350
rect 399430 454294 399498 454350
rect 399554 454294 399622 454350
rect 399678 454294 399774 454350
rect 399154 454226 399774 454294
rect 399154 454170 399250 454226
rect 399306 454170 399374 454226
rect 399430 454170 399498 454226
rect 399554 454170 399622 454226
rect 399678 454170 399774 454226
rect 399154 454102 399774 454170
rect 399154 454046 399250 454102
rect 399306 454046 399374 454102
rect 399430 454046 399498 454102
rect 399554 454046 399622 454102
rect 399678 454046 399774 454102
rect 399154 453978 399774 454046
rect 399154 453922 399250 453978
rect 399306 453922 399374 453978
rect 399430 453922 399498 453978
rect 399554 453922 399622 453978
rect 399678 453922 399774 453978
rect 399154 436350 399774 453922
rect 399154 436294 399250 436350
rect 399306 436294 399374 436350
rect 399430 436294 399498 436350
rect 399554 436294 399622 436350
rect 399678 436294 399774 436350
rect 399154 436226 399774 436294
rect 399154 436170 399250 436226
rect 399306 436170 399374 436226
rect 399430 436170 399498 436226
rect 399554 436170 399622 436226
rect 399678 436170 399774 436226
rect 399154 436102 399774 436170
rect 399154 436046 399250 436102
rect 399306 436046 399374 436102
rect 399430 436046 399498 436102
rect 399554 436046 399622 436102
rect 399678 436046 399774 436102
rect 399154 435978 399774 436046
rect 399154 435922 399250 435978
rect 399306 435922 399374 435978
rect 399430 435922 399498 435978
rect 399554 435922 399622 435978
rect 399678 435922 399774 435978
rect 399154 418350 399774 435922
rect 399154 418294 399250 418350
rect 399306 418294 399374 418350
rect 399430 418294 399498 418350
rect 399554 418294 399622 418350
rect 399678 418294 399774 418350
rect 399154 418226 399774 418294
rect 399154 418170 399250 418226
rect 399306 418170 399374 418226
rect 399430 418170 399498 418226
rect 399554 418170 399622 418226
rect 399678 418170 399774 418226
rect 399154 418102 399774 418170
rect 399154 418046 399250 418102
rect 399306 418046 399374 418102
rect 399430 418046 399498 418102
rect 399554 418046 399622 418102
rect 399678 418046 399774 418102
rect 399154 417978 399774 418046
rect 399154 417922 399250 417978
rect 399306 417922 399374 417978
rect 399430 417922 399498 417978
rect 399554 417922 399622 417978
rect 399678 417922 399774 417978
rect 399154 400350 399774 417922
rect 399154 400294 399250 400350
rect 399306 400294 399374 400350
rect 399430 400294 399498 400350
rect 399554 400294 399622 400350
rect 399678 400294 399774 400350
rect 399154 400226 399774 400294
rect 399154 400170 399250 400226
rect 399306 400170 399374 400226
rect 399430 400170 399498 400226
rect 399554 400170 399622 400226
rect 399678 400170 399774 400226
rect 399154 400102 399774 400170
rect 399154 400046 399250 400102
rect 399306 400046 399374 400102
rect 399430 400046 399498 400102
rect 399554 400046 399622 400102
rect 399678 400046 399774 400102
rect 399154 399978 399774 400046
rect 399154 399922 399250 399978
rect 399306 399922 399374 399978
rect 399430 399922 399498 399978
rect 399554 399922 399622 399978
rect 399678 399922 399774 399978
rect 399154 382350 399774 399922
rect 399154 382294 399250 382350
rect 399306 382294 399374 382350
rect 399430 382294 399498 382350
rect 399554 382294 399622 382350
rect 399678 382294 399774 382350
rect 399154 382226 399774 382294
rect 399154 382170 399250 382226
rect 399306 382170 399374 382226
rect 399430 382170 399498 382226
rect 399554 382170 399622 382226
rect 399678 382170 399774 382226
rect 399154 382102 399774 382170
rect 399154 382046 399250 382102
rect 399306 382046 399374 382102
rect 399430 382046 399498 382102
rect 399554 382046 399622 382102
rect 399678 382046 399774 382102
rect 399154 381978 399774 382046
rect 399154 381922 399250 381978
rect 399306 381922 399374 381978
rect 399430 381922 399498 381978
rect 399554 381922 399622 381978
rect 399678 381922 399774 381978
rect 399154 364350 399774 381922
rect 399154 364294 399250 364350
rect 399306 364294 399374 364350
rect 399430 364294 399498 364350
rect 399554 364294 399622 364350
rect 399678 364294 399774 364350
rect 399154 364226 399774 364294
rect 399154 364170 399250 364226
rect 399306 364170 399374 364226
rect 399430 364170 399498 364226
rect 399554 364170 399622 364226
rect 399678 364170 399774 364226
rect 399154 364102 399774 364170
rect 399154 364046 399250 364102
rect 399306 364046 399374 364102
rect 399430 364046 399498 364102
rect 399554 364046 399622 364102
rect 399678 364046 399774 364102
rect 399154 363978 399774 364046
rect 399154 363922 399250 363978
rect 399306 363922 399374 363978
rect 399430 363922 399498 363978
rect 399554 363922 399622 363978
rect 399678 363922 399774 363978
rect 399154 346350 399774 363922
rect 399154 346294 399250 346350
rect 399306 346294 399374 346350
rect 399430 346294 399498 346350
rect 399554 346294 399622 346350
rect 399678 346294 399774 346350
rect 399154 346226 399774 346294
rect 399154 346170 399250 346226
rect 399306 346170 399374 346226
rect 399430 346170 399498 346226
rect 399554 346170 399622 346226
rect 399678 346170 399774 346226
rect 399154 346102 399774 346170
rect 399154 346046 399250 346102
rect 399306 346046 399374 346102
rect 399430 346046 399498 346102
rect 399554 346046 399622 346102
rect 399678 346046 399774 346102
rect 399154 345978 399774 346046
rect 399154 345922 399250 345978
rect 399306 345922 399374 345978
rect 399430 345922 399498 345978
rect 399554 345922 399622 345978
rect 399678 345922 399774 345978
rect 399154 328350 399774 345922
rect 399154 328294 399250 328350
rect 399306 328294 399374 328350
rect 399430 328294 399498 328350
rect 399554 328294 399622 328350
rect 399678 328294 399774 328350
rect 399154 328226 399774 328294
rect 399154 328170 399250 328226
rect 399306 328170 399374 328226
rect 399430 328170 399498 328226
rect 399554 328170 399622 328226
rect 399678 328170 399774 328226
rect 399154 328102 399774 328170
rect 399154 328046 399250 328102
rect 399306 328046 399374 328102
rect 399430 328046 399498 328102
rect 399554 328046 399622 328102
rect 399678 328046 399774 328102
rect 399154 327978 399774 328046
rect 399154 327922 399250 327978
rect 399306 327922 399374 327978
rect 399430 327922 399498 327978
rect 399554 327922 399622 327978
rect 399678 327922 399774 327978
rect 399154 310350 399774 327922
rect 399154 310294 399250 310350
rect 399306 310294 399374 310350
rect 399430 310294 399498 310350
rect 399554 310294 399622 310350
rect 399678 310294 399774 310350
rect 399154 310226 399774 310294
rect 399154 310170 399250 310226
rect 399306 310170 399374 310226
rect 399430 310170 399498 310226
rect 399554 310170 399622 310226
rect 399678 310170 399774 310226
rect 399154 310102 399774 310170
rect 399154 310046 399250 310102
rect 399306 310046 399374 310102
rect 399430 310046 399498 310102
rect 399554 310046 399622 310102
rect 399678 310046 399774 310102
rect 399154 309978 399774 310046
rect 399154 309922 399250 309978
rect 399306 309922 399374 309978
rect 399430 309922 399498 309978
rect 399554 309922 399622 309978
rect 399678 309922 399774 309978
rect 399154 292350 399774 309922
rect 399154 292294 399250 292350
rect 399306 292294 399374 292350
rect 399430 292294 399498 292350
rect 399554 292294 399622 292350
rect 399678 292294 399774 292350
rect 399154 292226 399774 292294
rect 399154 292170 399250 292226
rect 399306 292170 399374 292226
rect 399430 292170 399498 292226
rect 399554 292170 399622 292226
rect 399678 292170 399774 292226
rect 399154 292102 399774 292170
rect 399154 292046 399250 292102
rect 399306 292046 399374 292102
rect 399430 292046 399498 292102
rect 399554 292046 399622 292102
rect 399678 292046 399774 292102
rect 399154 291978 399774 292046
rect 399154 291922 399250 291978
rect 399306 291922 399374 291978
rect 399430 291922 399498 291978
rect 399554 291922 399622 291978
rect 399678 291922 399774 291978
rect 399154 274350 399774 291922
rect 399154 274294 399250 274350
rect 399306 274294 399374 274350
rect 399430 274294 399498 274350
rect 399554 274294 399622 274350
rect 399678 274294 399774 274350
rect 399154 274226 399774 274294
rect 399154 274170 399250 274226
rect 399306 274170 399374 274226
rect 399430 274170 399498 274226
rect 399554 274170 399622 274226
rect 399678 274170 399774 274226
rect 399154 274102 399774 274170
rect 399154 274046 399250 274102
rect 399306 274046 399374 274102
rect 399430 274046 399498 274102
rect 399554 274046 399622 274102
rect 399678 274046 399774 274102
rect 399154 273978 399774 274046
rect 399154 273922 399250 273978
rect 399306 273922 399374 273978
rect 399430 273922 399498 273978
rect 399554 273922 399622 273978
rect 399678 273922 399774 273978
rect 399154 256350 399774 273922
rect 399154 256294 399250 256350
rect 399306 256294 399374 256350
rect 399430 256294 399498 256350
rect 399554 256294 399622 256350
rect 399678 256294 399774 256350
rect 399154 256226 399774 256294
rect 399154 256170 399250 256226
rect 399306 256170 399374 256226
rect 399430 256170 399498 256226
rect 399554 256170 399622 256226
rect 399678 256170 399774 256226
rect 399154 256102 399774 256170
rect 399154 256046 399250 256102
rect 399306 256046 399374 256102
rect 399430 256046 399498 256102
rect 399554 256046 399622 256102
rect 399678 256046 399774 256102
rect 399154 255978 399774 256046
rect 399154 255922 399250 255978
rect 399306 255922 399374 255978
rect 399430 255922 399498 255978
rect 399554 255922 399622 255978
rect 399678 255922 399774 255978
rect 399154 238350 399774 255922
rect 399154 238294 399250 238350
rect 399306 238294 399374 238350
rect 399430 238294 399498 238350
rect 399554 238294 399622 238350
rect 399678 238294 399774 238350
rect 399154 238226 399774 238294
rect 399154 238170 399250 238226
rect 399306 238170 399374 238226
rect 399430 238170 399498 238226
rect 399554 238170 399622 238226
rect 399678 238170 399774 238226
rect 399154 238102 399774 238170
rect 399154 238046 399250 238102
rect 399306 238046 399374 238102
rect 399430 238046 399498 238102
rect 399554 238046 399622 238102
rect 399678 238046 399774 238102
rect 399154 237978 399774 238046
rect 399154 237922 399250 237978
rect 399306 237922 399374 237978
rect 399430 237922 399498 237978
rect 399554 237922 399622 237978
rect 399678 237922 399774 237978
rect 399154 220350 399774 237922
rect 399154 220294 399250 220350
rect 399306 220294 399374 220350
rect 399430 220294 399498 220350
rect 399554 220294 399622 220350
rect 399678 220294 399774 220350
rect 399154 220226 399774 220294
rect 399154 220170 399250 220226
rect 399306 220170 399374 220226
rect 399430 220170 399498 220226
rect 399554 220170 399622 220226
rect 399678 220170 399774 220226
rect 399154 220102 399774 220170
rect 399154 220046 399250 220102
rect 399306 220046 399374 220102
rect 399430 220046 399498 220102
rect 399554 220046 399622 220102
rect 399678 220046 399774 220102
rect 399154 219978 399774 220046
rect 399154 219922 399250 219978
rect 399306 219922 399374 219978
rect 399430 219922 399498 219978
rect 399554 219922 399622 219978
rect 399678 219922 399774 219978
rect 399154 217934 399774 219922
rect 402874 598172 403494 598268
rect 402874 598116 402970 598172
rect 403026 598116 403094 598172
rect 403150 598116 403218 598172
rect 403274 598116 403342 598172
rect 403398 598116 403494 598172
rect 402874 598048 403494 598116
rect 402874 597992 402970 598048
rect 403026 597992 403094 598048
rect 403150 597992 403218 598048
rect 403274 597992 403342 598048
rect 403398 597992 403494 598048
rect 402874 597924 403494 597992
rect 402874 597868 402970 597924
rect 403026 597868 403094 597924
rect 403150 597868 403218 597924
rect 403274 597868 403342 597924
rect 403398 597868 403494 597924
rect 402874 597800 403494 597868
rect 402874 597744 402970 597800
rect 403026 597744 403094 597800
rect 403150 597744 403218 597800
rect 403274 597744 403342 597800
rect 403398 597744 403494 597800
rect 402874 586350 403494 597744
rect 417154 597212 417774 598268
rect 417154 597156 417250 597212
rect 417306 597156 417374 597212
rect 417430 597156 417498 597212
rect 417554 597156 417622 597212
rect 417678 597156 417774 597212
rect 417154 597088 417774 597156
rect 417154 597032 417250 597088
rect 417306 597032 417374 597088
rect 417430 597032 417498 597088
rect 417554 597032 417622 597088
rect 417678 597032 417774 597088
rect 417154 596964 417774 597032
rect 417154 596908 417250 596964
rect 417306 596908 417374 596964
rect 417430 596908 417498 596964
rect 417554 596908 417622 596964
rect 417678 596908 417774 596964
rect 417154 596840 417774 596908
rect 417154 596784 417250 596840
rect 417306 596784 417374 596840
rect 417430 596784 417498 596840
rect 417554 596784 417622 596840
rect 417678 596784 417774 596840
rect 408380 589764 408436 589774
rect 408380 588868 408436 589708
rect 408380 588802 408436 588812
rect 402874 586294 402970 586350
rect 403026 586294 403094 586350
rect 403150 586294 403218 586350
rect 403274 586294 403342 586350
rect 403398 586294 403494 586350
rect 402874 586226 403494 586294
rect 402874 586170 402970 586226
rect 403026 586170 403094 586226
rect 403150 586170 403218 586226
rect 403274 586170 403342 586226
rect 403398 586170 403494 586226
rect 402874 586102 403494 586170
rect 402874 586046 402970 586102
rect 403026 586046 403094 586102
rect 403150 586046 403218 586102
rect 403274 586046 403342 586102
rect 403398 586046 403494 586102
rect 402874 585978 403494 586046
rect 402874 585922 402970 585978
rect 403026 585922 403094 585978
rect 403150 585922 403218 585978
rect 403274 585922 403342 585978
rect 403398 585922 403494 585978
rect 402874 568350 403494 585922
rect 402874 568294 402970 568350
rect 403026 568294 403094 568350
rect 403150 568294 403218 568350
rect 403274 568294 403342 568350
rect 403398 568294 403494 568350
rect 402874 568226 403494 568294
rect 402874 568170 402970 568226
rect 403026 568170 403094 568226
rect 403150 568170 403218 568226
rect 403274 568170 403342 568226
rect 403398 568170 403494 568226
rect 402874 568102 403494 568170
rect 402874 568046 402970 568102
rect 403026 568046 403094 568102
rect 403150 568046 403218 568102
rect 403274 568046 403342 568102
rect 403398 568046 403494 568102
rect 402874 567978 403494 568046
rect 402874 567922 402970 567978
rect 403026 567922 403094 567978
rect 403150 567922 403218 567978
rect 403274 567922 403342 567978
rect 403398 567922 403494 567978
rect 402874 550350 403494 567922
rect 402874 550294 402970 550350
rect 403026 550294 403094 550350
rect 403150 550294 403218 550350
rect 403274 550294 403342 550350
rect 403398 550294 403494 550350
rect 402874 550226 403494 550294
rect 402874 550170 402970 550226
rect 403026 550170 403094 550226
rect 403150 550170 403218 550226
rect 403274 550170 403342 550226
rect 403398 550170 403494 550226
rect 402874 550102 403494 550170
rect 402874 550046 402970 550102
rect 403026 550046 403094 550102
rect 403150 550046 403218 550102
rect 403274 550046 403342 550102
rect 403398 550046 403494 550102
rect 402874 549978 403494 550046
rect 402874 549922 402970 549978
rect 403026 549922 403094 549978
rect 403150 549922 403218 549978
rect 403274 549922 403342 549978
rect 403398 549922 403494 549978
rect 402874 532350 403494 549922
rect 402874 532294 402970 532350
rect 403026 532294 403094 532350
rect 403150 532294 403218 532350
rect 403274 532294 403342 532350
rect 403398 532294 403494 532350
rect 402874 532226 403494 532294
rect 402874 532170 402970 532226
rect 403026 532170 403094 532226
rect 403150 532170 403218 532226
rect 403274 532170 403342 532226
rect 403398 532170 403494 532226
rect 402874 532102 403494 532170
rect 402874 532046 402970 532102
rect 403026 532046 403094 532102
rect 403150 532046 403218 532102
rect 403274 532046 403342 532102
rect 403398 532046 403494 532102
rect 402874 531978 403494 532046
rect 402874 531922 402970 531978
rect 403026 531922 403094 531978
rect 403150 531922 403218 531978
rect 403274 531922 403342 531978
rect 403398 531922 403494 531978
rect 402874 514350 403494 531922
rect 402874 514294 402970 514350
rect 403026 514294 403094 514350
rect 403150 514294 403218 514350
rect 403274 514294 403342 514350
rect 403398 514294 403494 514350
rect 402874 514226 403494 514294
rect 402874 514170 402970 514226
rect 403026 514170 403094 514226
rect 403150 514170 403218 514226
rect 403274 514170 403342 514226
rect 403398 514170 403494 514226
rect 402874 514102 403494 514170
rect 402874 514046 402970 514102
rect 403026 514046 403094 514102
rect 403150 514046 403218 514102
rect 403274 514046 403342 514102
rect 403398 514046 403494 514102
rect 402874 513978 403494 514046
rect 402874 513922 402970 513978
rect 403026 513922 403094 513978
rect 403150 513922 403218 513978
rect 403274 513922 403342 513978
rect 403398 513922 403494 513978
rect 402874 496350 403494 513922
rect 402874 496294 402970 496350
rect 403026 496294 403094 496350
rect 403150 496294 403218 496350
rect 403274 496294 403342 496350
rect 403398 496294 403494 496350
rect 402874 496226 403494 496294
rect 402874 496170 402970 496226
rect 403026 496170 403094 496226
rect 403150 496170 403218 496226
rect 403274 496170 403342 496226
rect 403398 496170 403494 496226
rect 402874 496102 403494 496170
rect 402874 496046 402970 496102
rect 403026 496046 403094 496102
rect 403150 496046 403218 496102
rect 403274 496046 403342 496102
rect 403398 496046 403494 496102
rect 402874 495978 403494 496046
rect 402874 495922 402970 495978
rect 403026 495922 403094 495978
rect 403150 495922 403218 495978
rect 403274 495922 403342 495978
rect 403398 495922 403494 495978
rect 402874 478350 403494 495922
rect 402874 478294 402970 478350
rect 403026 478294 403094 478350
rect 403150 478294 403218 478350
rect 403274 478294 403342 478350
rect 403398 478294 403494 478350
rect 402874 478226 403494 478294
rect 402874 478170 402970 478226
rect 403026 478170 403094 478226
rect 403150 478170 403218 478226
rect 403274 478170 403342 478226
rect 403398 478170 403494 478226
rect 402874 478102 403494 478170
rect 402874 478046 402970 478102
rect 403026 478046 403094 478102
rect 403150 478046 403218 478102
rect 403274 478046 403342 478102
rect 403398 478046 403494 478102
rect 402874 477978 403494 478046
rect 402874 477922 402970 477978
rect 403026 477922 403094 477978
rect 403150 477922 403218 477978
rect 403274 477922 403342 477978
rect 403398 477922 403494 477978
rect 402874 460350 403494 477922
rect 402874 460294 402970 460350
rect 403026 460294 403094 460350
rect 403150 460294 403218 460350
rect 403274 460294 403342 460350
rect 403398 460294 403494 460350
rect 402874 460226 403494 460294
rect 402874 460170 402970 460226
rect 403026 460170 403094 460226
rect 403150 460170 403218 460226
rect 403274 460170 403342 460226
rect 403398 460170 403494 460226
rect 402874 460102 403494 460170
rect 402874 460046 402970 460102
rect 403026 460046 403094 460102
rect 403150 460046 403218 460102
rect 403274 460046 403342 460102
rect 403398 460046 403494 460102
rect 402874 459978 403494 460046
rect 402874 459922 402970 459978
rect 403026 459922 403094 459978
rect 403150 459922 403218 459978
rect 403274 459922 403342 459978
rect 403398 459922 403494 459978
rect 402874 442350 403494 459922
rect 402874 442294 402970 442350
rect 403026 442294 403094 442350
rect 403150 442294 403218 442350
rect 403274 442294 403342 442350
rect 403398 442294 403494 442350
rect 402874 442226 403494 442294
rect 402874 442170 402970 442226
rect 403026 442170 403094 442226
rect 403150 442170 403218 442226
rect 403274 442170 403342 442226
rect 403398 442170 403494 442226
rect 402874 442102 403494 442170
rect 402874 442046 402970 442102
rect 403026 442046 403094 442102
rect 403150 442046 403218 442102
rect 403274 442046 403342 442102
rect 403398 442046 403494 442102
rect 402874 441978 403494 442046
rect 402874 441922 402970 441978
rect 403026 441922 403094 441978
rect 403150 441922 403218 441978
rect 403274 441922 403342 441978
rect 403398 441922 403494 441978
rect 402874 424350 403494 441922
rect 402874 424294 402970 424350
rect 403026 424294 403094 424350
rect 403150 424294 403218 424350
rect 403274 424294 403342 424350
rect 403398 424294 403494 424350
rect 402874 424226 403494 424294
rect 402874 424170 402970 424226
rect 403026 424170 403094 424226
rect 403150 424170 403218 424226
rect 403274 424170 403342 424226
rect 403398 424170 403494 424226
rect 402874 424102 403494 424170
rect 402874 424046 402970 424102
rect 403026 424046 403094 424102
rect 403150 424046 403218 424102
rect 403274 424046 403342 424102
rect 403398 424046 403494 424102
rect 402874 423978 403494 424046
rect 402874 423922 402970 423978
rect 403026 423922 403094 423978
rect 403150 423922 403218 423978
rect 403274 423922 403342 423978
rect 403398 423922 403494 423978
rect 402874 406350 403494 423922
rect 402874 406294 402970 406350
rect 403026 406294 403094 406350
rect 403150 406294 403218 406350
rect 403274 406294 403342 406350
rect 403398 406294 403494 406350
rect 402874 406226 403494 406294
rect 402874 406170 402970 406226
rect 403026 406170 403094 406226
rect 403150 406170 403218 406226
rect 403274 406170 403342 406226
rect 403398 406170 403494 406226
rect 402874 406102 403494 406170
rect 402874 406046 402970 406102
rect 403026 406046 403094 406102
rect 403150 406046 403218 406102
rect 403274 406046 403342 406102
rect 403398 406046 403494 406102
rect 402874 405978 403494 406046
rect 402874 405922 402970 405978
rect 403026 405922 403094 405978
rect 403150 405922 403218 405978
rect 403274 405922 403342 405978
rect 403398 405922 403494 405978
rect 402874 388350 403494 405922
rect 402874 388294 402970 388350
rect 403026 388294 403094 388350
rect 403150 388294 403218 388350
rect 403274 388294 403342 388350
rect 403398 388294 403494 388350
rect 402874 388226 403494 388294
rect 402874 388170 402970 388226
rect 403026 388170 403094 388226
rect 403150 388170 403218 388226
rect 403274 388170 403342 388226
rect 403398 388170 403494 388226
rect 402874 388102 403494 388170
rect 402874 388046 402970 388102
rect 403026 388046 403094 388102
rect 403150 388046 403218 388102
rect 403274 388046 403342 388102
rect 403398 388046 403494 388102
rect 402874 387978 403494 388046
rect 402874 387922 402970 387978
rect 403026 387922 403094 387978
rect 403150 387922 403218 387978
rect 403274 387922 403342 387978
rect 403398 387922 403494 387978
rect 402874 370350 403494 387922
rect 402874 370294 402970 370350
rect 403026 370294 403094 370350
rect 403150 370294 403218 370350
rect 403274 370294 403342 370350
rect 403398 370294 403494 370350
rect 402874 370226 403494 370294
rect 402874 370170 402970 370226
rect 403026 370170 403094 370226
rect 403150 370170 403218 370226
rect 403274 370170 403342 370226
rect 403398 370170 403494 370226
rect 402874 370102 403494 370170
rect 402874 370046 402970 370102
rect 403026 370046 403094 370102
rect 403150 370046 403218 370102
rect 403274 370046 403342 370102
rect 403398 370046 403494 370102
rect 402874 369978 403494 370046
rect 402874 369922 402970 369978
rect 403026 369922 403094 369978
rect 403150 369922 403218 369978
rect 403274 369922 403342 369978
rect 403398 369922 403494 369978
rect 402874 352350 403494 369922
rect 402874 352294 402970 352350
rect 403026 352294 403094 352350
rect 403150 352294 403218 352350
rect 403274 352294 403342 352350
rect 403398 352294 403494 352350
rect 402874 352226 403494 352294
rect 402874 352170 402970 352226
rect 403026 352170 403094 352226
rect 403150 352170 403218 352226
rect 403274 352170 403342 352226
rect 403398 352170 403494 352226
rect 402874 352102 403494 352170
rect 402874 352046 402970 352102
rect 403026 352046 403094 352102
rect 403150 352046 403218 352102
rect 403274 352046 403342 352102
rect 403398 352046 403494 352102
rect 402874 351978 403494 352046
rect 402874 351922 402970 351978
rect 403026 351922 403094 351978
rect 403150 351922 403218 351978
rect 403274 351922 403342 351978
rect 403398 351922 403494 351978
rect 402874 334350 403494 351922
rect 402874 334294 402970 334350
rect 403026 334294 403094 334350
rect 403150 334294 403218 334350
rect 403274 334294 403342 334350
rect 403398 334294 403494 334350
rect 402874 334226 403494 334294
rect 402874 334170 402970 334226
rect 403026 334170 403094 334226
rect 403150 334170 403218 334226
rect 403274 334170 403342 334226
rect 403398 334170 403494 334226
rect 402874 334102 403494 334170
rect 402874 334046 402970 334102
rect 403026 334046 403094 334102
rect 403150 334046 403218 334102
rect 403274 334046 403342 334102
rect 403398 334046 403494 334102
rect 402874 333978 403494 334046
rect 402874 333922 402970 333978
rect 403026 333922 403094 333978
rect 403150 333922 403218 333978
rect 403274 333922 403342 333978
rect 403398 333922 403494 333978
rect 402874 316350 403494 333922
rect 402874 316294 402970 316350
rect 403026 316294 403094 316350
rect 403150 316294 403218 316350
rect 403274 316294 403342 316350
rect 403398 316294 403494 316350
rect 402874 316226 403494 316294
rect 402874 316170 402970 316226
rect 403026 316170 403094 316226
rect 403150 316170 403218 316226
rect 403274 316170 403342 316226
rect 403398 316170 403494 316226
rect 402874 316102 403494 316170
rect 402874 316046 402970 316102
rect 403026 316046 403094 316102
rect 403150 316046 403218 316102
rect 403274 316046 403342 316102
rect 403398 316046 403494 316102
rect 402874 315978 403494 316046
rect 402874 315922 402970 315978
rect 403026 315922 403094 315978
rect 403150 315922 403218 315978
rect 403274 315922 403342 315978
rect 403398 315922 403494 315978
rect 402874 298350 403494 315922
rect 402874 298294 402970 298350
rect 403026 298294 403094 298350
rect 403150 298294 403218 298350
rect 403274 298294 403342 298350
rect 403398 298294 403494 298350
rect 402874 298226 403494 298294
rect 402874 298170 402970 298226
rect 403026 298170 403094 298226
rect 403150 298170 403218 298226
rect 403274 298170 403342 298226
rect 403398 298170 403494 298226
rect 402874 298102 403494 298170
rect 402874 298046 402970 298102
rect 403026 298046 403094 298102
rect 403150 298046 403218 298102
rect 403274 298046 403342 298102
rect 403398 298046 403494 298102
rect 402874 297978 403494 298046
rect 402874 297922 402970 297978
rect 403026 297922 403094 297978
rect 403150 297922 403218 297978
rect 403274 297922 403342 297978
rect 403398 297922 403494 297978
rect 402874 280350 403494 297922
rect 402874 280294 402970 280350
rect 403026 280294 403094 280350
rect 403150 280294 403218 280350
rect 403274 280294 403342 280350
rect 403398 280294 403494 280350
rect 402874 280226 403494 280294
rect 402874 280170 402970 280226
rect 403026 280170 403094 280226
rect 403150 280170 403218 280226
rect 403274 280170 403342 280226
rect 403398 280170 403494 280226
rect 402874 280102 403494 280170
rect 402874 280046 402970 280102
rect 403026 280046 403094 280102
rect 403150 280046 403218 280102
rect 403274 280046 403342 280102
rect 403398 280046 403494 280102
rect 402874 279978 403494 280046
rect 402874 279922 402970 279978
rect 403026 279922 403094 279978
rect 403150 279922 403218 279978
rect 403274 279922 403342 279978
rect 403398 279922 403494 279978
rect 402874 262350 403494 279922
rect 402874 262294 402970 262350
rect 403026 262294 403094 262350
rect 403150 262294 403218 262350
rect 403274 262294 403342 262350
rect 403398 262294 403494 262350
rect 402874 262226 403494 262294
rect 402874 262170 402970 262226
rect 403026 262170 403094 262226
rect 403150 262170 403218 262226
rect 403274 262170 403342 262226
rect 403398 262170 403494 262226
rect 402874 262102 403494 262170
rect 402874 262046 402970 262102
rect 403026 262046 403094 262102
rect 403150 262046 403218 262102
rect 403274 262046 403342 262102
rect 403398 262046 403494 262102
rect 402874 261978 403494 262046
rect 402874 261922 402970 261978
rect 403026 261922 403094 261978
rect 403150 261922 403218 261978
rect 403274 261922 403342 261978
rect 403398 261922 403494 261978
rect 402874 244350 403494 261922
rect 402874 244294 402970 244350
rect 403026 244294 403094 244350
rect 403150 244294 403218 244350
rect 403274 244294 403342 244350
rect 403398 244294 403494 244350
rect 402874 244226 403494 244294
rect 402874 244170 402970 244226
rect 403026 244170 403094 244226
rect 403150 244170 403218 244226
rect 403274 244170 403342 244226
rect 403398 244170 403494 244226
rect 402874 244102 403494 244170
rect 402874 244046 402970 244102
rect 403026 244046 403094 244102
rect 403150 244046 403218 244102
rect 403274 244046 403342 244102
rect 403398 244046 403494 244102
rect 402874 243978 403494 244046
rect 402874 243922 402970 243978
rect 403026 243922 403094 243978
rect 403150 243922 403218 243978
rect 403274 243922 403342 243978
rect 403398 243922 403494 243978
rect 402874 226350 403494 243922
rect 402874 226294 402970 226350
rect 403026 226294 403094 226350
rect 403150 226294 403218 226350
rect 403274 226294 403342 226350
rect 403398 226294 403494 226350
rect 402874 226226 403494 226294
rect 402874 226170 402970 226226
rect 403026 226170 403094 226226
rect 403150 226170 403218 226226
rect 403274 226170 403342 226226
rect 403398 226170 403494 226226
rect 402874 226102 403494 226170
rect 402874 226046 402970 226102
rect 403026 226046 403094 226102
rect 403150 226046 403218 226102
rect 403274 226046 403342 226102
rect 403398 226046 403494 226102
rect 402874 225978 403494 226046
rect 402874 225922 402970 225978
rect 403026 225922 403094 225978
rect 403150 225922 403218 225978
rect 403274 225922 403342 225978
rect 403398 225922 403494 225978
rect 402874 217934 403494 225922
rect 417154 580350 417774 596784
rect 417154 580294 417250 580350
rect 417306 580294 417374 580350
rect 417430 580294 417498 580350
rect 417554 580294 417622 580350
rect 417678 580294 417774 580350
rect 417154 580226 417774 580294
rect 417154 580170 417250 580226
rect 417306 580170 417374 580226
rect 417430 580170 417498 580226
rect 417554 580170 417622 580226
rect 417678 580170 417774 580226
rect 417154 580102 417774 580170
rect 417154 580046 417250 580102
rect 417306 580046 417374 580102
rect 417430 580046 417498 580102
rect 417554 580046 417622 580102
rect 417678 580046 417774 580102
rect 417154 579978 417774 580046
rect 417154 579922 417250 579978
rect 417306 579922 417374 579978
rect 417430 579922 417498 579978
rect 417554 579922 417622 579978
rect 417678 579922 417774 579978
rect 417154 562350 417774 579922
rect 417154 562294 417250 562350
rect 417306 562294 417374 562350
rect 417430 562294 417498 562350
rect 417554 562294 417622 562350
rect 417678 562294 417774 562350
rect 417154 562226 417774 562294
rect 417154 562170 417250 562226
rect 417306 562170 417374 562226
rect 417430 562170 417498 562226
rect 417554 562170 417622 562226
rect 417678 562170 417774 562226
rect 417154 562102 417774 562170
rect 417154 562046 417250 562102
rect 417306 562046 417374 562102
rect 417430 562046 417498 562102
rect 417554 562046 417622 562102
rect 417678 562046 417774 562102
rect 417154 561978 417774 562046
rect 417154 561922 417250 561978
rect 417306 561922 417374 561978
rect 417430 561922 417498 561978
rect 417554 561922 417622 561978
rect 417678 561922 417774 561978
rect 417154 544350 417774 561922
rect 417154 544294 417250 544350
rect 417306 544294 417374 544350
rect 417430 544294 417498 544350
rect 417554 544294 417622 544350
rect 417678 544294 417774 544350
rect 417154 544226 417774 544294
rect 417154 544170 417250 544226
rect 417306 544170 417374 544226
rect 417430 544170 417498 544226
rect 417554 544170 417622 544226
rect 417678 544170 417774 544226
rect 417154 544102 417774 544170
rect 417154 544046 417250 544102
rect 417306 544046 417374 544102
rect 417430 544046 417498 544102
rect 417554 544046 417622 544102
rect 417678 544046 417774 544102
rect 417154 543978 417774 544046
rect 417154 543922 417250 543978
rect 417306 543922 417374 543978
rect 417430 543922 417498 543978
rect 417554 543922 417622 543978
rect 417678 543922 417774 543978
rect 417154 526350 417774 543922
rect 417154 526294 417250 526350
rect 417306 526294 417374 526350
rect 417430 526294 417498 526350
rect 417554 526294 417622 526350
rect 417678 526294 417774 526350
rect 417154 526226 417774 526294
rect 417154 526170 417250 526226
rect 417306 526170 417374 526226
rect 417430 526170 417498 526226
rect 417554 526170 417622 526226
rect 417678 526170 417774 526226
rect 417154 526102 417774 526170
rect 417154 526046 417250 526102
rect 417306 526046 417374 526102
rect 417430 526046 417498 526102
rect 417554 526046 417622 526102
rect 417678 526046 417774 526102
rect 417154 525978 417774 526046
rect 417154 525922 417250 525978
rect 417306 525922 417374 525978
rect 417430 525922 417498 525978
rect 417554 525922 417622 525978
rect 417678 525922 417774 525978
rect 417154 508350 417774 525922
rect 417154 508294 417250 508350
rect 417306 508294 417374 508350
rect 417430 508294 417498 508350
rect 417554 508294 417622 508350
rect 417678 508294 417774 508350
rect 417154 508226 417774 508294
rect 417154 508170 417250 508226
rect 417306 508170 417374 508226
rect 417430 508170 417498 508226
rect 417554 508170 417622 508226
rect 417678 508170 417774 508226
rect 417154 508102 417774 508170
rect 417154 508046 417250 508102
rect 417306 508046 417374 508102
rect 417430 508046 417498 508102
rect 417554 508046 417622 508102
rect 417678 508046 417774 508102
rect 417154 507978 417774 508046
rect 417154 507922 417250 507978
rect 417306 507922 417374 507978
rect 417430 507922 417498 507978
rect 417554 507922 417622 507978
rect 417678 507922 417774 507978
rect 417154 490350 417774 507922
rect 417154 490294 417250 490350
rect 417306 490294 417374 490350
rect 417430 490294 417498 490350
rect 417554 490294 417622 490350
rect 417678 490294 417774 490350
rect 417154 490226 417774 490294
rect 417154 490170 417250 490226
rect 417306 490170 417374 490226
rect 417430 490170 417498 490226
rect 417554 490170 417622 490226
rect 417678 490170 417774 490226
rect 417154 490102 417774 490170
rect 417154 490046 417250 490102
rect 417306 490046 417374 490102
rect 417430 490046 417498 490102
rect 417554 490046 417622 490102
rect 417678 490046 417774 490102
rect 417154 489978 417774 490046
rect 417154 489922 417250 489978
rect 417306 489922 417374 489978
rect 417430 489922 417498 489978
rect 417554 489922 417622 489978
rect 417678 489922 417774 489978
rect 417154 472350 417774 489922
rect 417154 472294 417250 472350
rect 417306 472294 417374 472350
rect 417430 472294 417498 472350
rect 417554 472294 417622 472350
rect 417678 472294 417774 472350
rect 417154 472226 417774 472294
rect 417154 472170 417250 472226
rect 417306 472170 417374 472226
rect 417430 472170 417498 472226
rect 417554 472170 417622 472226
rect 417678 472170 417774 472226
rect 417154 472102 417774 472170
rect 417154 472046 417250 472102
rect 417306 472046 417374 472102
rect 417430 472046 417498 472102
rect 417554 472046 417622 472102
rect 417678 472046 417774 472102
rect 417154 471978 417774 472046
rect 417154 471922 417250 471978
rect 417306 471922 417374 471978
rect 417430 471922 417498 471978
rect 417554 471922 417622 471978
rect 417678 471922 417774 471978
rect 417154 454350 417774 471922
rect 417154 454294 417250 454350
rect 417306 454294 417374 454350
rect 417430 454294 417498 454350
rect 417554 454294 417622 454350
rect 417678 454294 417774 454350
rect 417154 454226 417774 454294
rect 417154 454170 417250 454226
rect 417306 454170 417374 454226
rect 417430 454170 417498 454226
rect 417554 454170 417622 454226
rect 417678 454170 417774 454226
rect 417154 454102 417774 454170
rect 417154 454046 417250 454102
rect 417306 454046 417374 454102
rect 417430 454046 417498 454102
rect 417554 454046 417622 454102
rect 417678 454046 417774 454102
rect 417154 453978 417774 454046
rect 417154 453922 417250 453978
rect 417306 453922 417374 453978
rect 417430 453922 417498 453978
rect 417554 453922 417622 453978
rect 417678 453922 417774 453978
rect 417154 436350 417774 453922
rect 417154 436294 417250 436350
rect 417306 436294 417374 436350
rect 417430 436294 417498 436350
rect 417554 436294 417622 436350
rect 417678 436294 417774 436350
rect 417154 436226 417774 436294
rect 417154 436170 417250 436226
rect 417306 436170 417374 436226
rect 417430 436170 417498 436226
rect 417554 436170 417622 436226
rect 417678 436170 417774 436226
rect 417154 436102 417774 436170
rect 417154 436046 417250 436102
rect 417306 436046 417374 436102
rect 417430 436046 417498 436102
rect 417554 436046 417622 436102
rect 417678 436046 417774 436102
rect 417154 435978 417774 436046
rect 417154 435922 417250 435978
rect 417306 435922 417374 435978
rect 417430 435922 417498 435978
rect 417554 435922 417622 435978
rect 417678 435922 417774 435978
rect 417154 418350 417774 435922
rect 417154 418294 417250 418350
rect 417306 418294 417374 418350
rect 417430 418294 417498 418350
rect 417554 418294 417622 418350
rect 417678 418294 417774 418350
rect 417154 418226 417774 418294
rect 417154 418170 417250 418226
rect 417306 418170 417374 418226
rect 417430 418170 417498 418226
rect 417554 418170 417622 418226
rect 417678 418170 417774 418226
rect 417154 418102 417774 418170
rect 417154 418046 417250 418102
rect 417306 418046 417374 418102
rect 417430 418046 417498 418102
rect 417554 418046 417622 418102
rect 417678 418046 417774 418102
rect 417154 417978 417774 418046
rect 417154 417922 417250 417978
rect 417306 417922 417374 417978
rect 417430 417922 417498 417978
rect 417554 417922 417622 417978
rect 417678 417922 417774 417978
rect 417154 400350 417774 417922
rect 417154 400294 417250 400350
rect 417306 400294 417374 400350
rect 417430 400294 417498 400350
rect 417554 400294 417622 400350
rect 417678 400294 417774 400350
rect 417154 400226 417774 400294
rect 417154 400170 417250 400226
rect 417306 400170 417374 400226
rect 417430 400170 417498 400226
rect 417554 400170 417622 400226
rect 417678 400170 417774 400226
rect 417154 400102 417774 400170
rect 417154 400046 417250 400102
rect 417306 400046 417374 400102
rect 417430 400046 417498 400102
rect 417554 400046 417622 400102
rect 417678 400046 417774 400102
rect 417154 399978 417774 400046
rect 417154 399922 417250 399978
rect 417306 399922 417374 399978
rect 417430 399922 417498 399978
rect 417554 399922 417622 399978
rect 417678 399922 417774 399978
rect 417154 382350 417774 399922
rect 417154 382294 417250 382350
rect 417306 382294 417374 382350
rect 417430 382294 417498 382350
rect 417554 382294 417622 382350
rect 417678 382294 417774 382350
rect 417154 382226 417774 382294
rect 417154 382170 417250 382226
rect 417306 382170 417374 382226
rect 417430 382170 417498 382226
rect 417554 382170 417622 382226
rect 417678 382170 417774 382226
rect 417154 382102 417774 382170
rect 417154 382046 417250 382102
rect 417306 382046 417374 382102
rect 417430 382046 417498 382102
rect 417554 382046 417622 382102
rect 417678 382046 417774 382102
rect 417154 381978 417774 382046
rect 417154 381922 417250 381978
rect 417306 381922 417374 381978
rect 417430 381922 417498 381978
rect 417554 381922 417622 381978
rect 417678 381922 417774 381978
rect 417154 364350 417774 381922
rect 417154 364294 417250 364350
rect 417306 364294 417374 364350
rect 417430 364294 417498 364350
rect 417554 364294 417622 364350
rect 417678 364294 417774 364350
rect 417154 364226 417774 364294
rect 417154 364170 417250 364226
rect 417306 364170 417374 364226
rect 417430 364170 417498 364226
rect 417554 364170 417622 364226
rect 417678 364170 417774 364226
rect 417154 364102 417774 364170
rect 417154 364046 417250 364102
rect 417306 364046 417374 364102
rect 417430 364046 417498 364102
rect 417554 364046 417622 364102
rect 417678 364046 417774 364102
rect 417154 363978 417774 364046
rect 417154 363922 417250 363978
rect 417306 363922 417374 363978
rect 417430 363922 417498 363978
rect 417554 363922 417622 363978
rect 417678 363922 417774 363978
rect 417154 346350 417774 363922
rect 417154 346294 417250 346350
rect 417306 346294 417374 346350
rect 417430 346294 417498 346350
rect 417554 346294 417622 346350
rect 417678 346294 417774 346350
rect 417154 346226 417774 346294
rect 417154 346170 417250 346226
rect 417306 346170 417374 346226
rect 417430 346170 417498 346226
rect 417554 346170 417622 346226
rect 417678 346170 417774 346226
rect 417154 346102 417774 346170
rect 417154 346046 417250 346102
rect 417306 346046 417374 346102
rect 417430 346046 417498 346102
rect 417554 346046 417622 346102
rect 417678 346046 417774 346102
rect 417154 345978 417774 346046
rect 417154 345922 417250 345978
rect 417306 345922 417374 345978
rect 417430 345922 417498 345978
rect 417554 345922 417622 345978
rect 417678 345922 417774 345978
rect 417154 328350 417774 345922
rect 417154 328294 417250 328350
rect 417306 328294 417374 328350
rect 417430 328294 417498 328350
rect 417554 328294 417622 328350
rect 417678 328294 417774 328350
rect 417154 328226 417774 328294
rect 417154 328170 417250 328226
rect 417306 328170 417374 328226
rect 417430 328170 417498 328226
rect 417554 328170 417622 328226
rect 417678 328170 417774 328226
rect 417154 328102 417774 328170
rect 417154 328046 417250 328102
rect 417306 328046 417374 328102
rect 417430 328046 417498 328102
rect 417554 328046 417622 328102
rect 417678 328046 417774 328102
rect 417154 327978 417774 328046
rect 417154 327922 417250 327978
rect 417306 327922 417374 327978
rect 417430 327922 417498 327978
rect 417554 327922 417622 327978
rect 417678 327922 417774 327978
rect 417154 310350 417774 327922
rect 417154 310294 417250 310350
rect 417306 310294 417374 310350
rect 417430 310294 417498 310350
rect 417554 310294 417622 310350
rect 417678 310294 417774 310350
rect 417154 310226 417774 310294
rect 417154 310170 417250 310226
rect 417306 310170 417374 310226
rect 417430 310170 417498 310226
rect 417554 310170 417622 310226
rect 417678 310170 417774 310226
rect 417154 310102 417774 310170
rect 417154 310046 417250 310102
rect 417306 310046 417374 310102
rect 417430 310046 417498 310102
rect 417554 310046 417622 310102
rect 417678 310046 417774 310102
rect 417154 309978 417774 310046
rect 417154 309922 417250 309978
rect 417306 309922 417374 309978
rect 417430 309922 417498 309978
rect 417554 309922 417622 309978
rect 417678 309922 417774 309978
rect 417154 292350 417774 309922
rect 417154 292294 417250 292350
rect 417306 292294 417374 292350
rect 417430 292294 417498 292350
rect 417554 292294 417622 292350
rect 417678 292294 417774 292350
rect 417154 292226 417774 292294
rect 417154 292170 417250 292226
rect 417306 292170 417374 292226
rect 417430 292170 417498 292226
rect 417554 292170 417622 292226
rect 417678 292170 417774 292226
rect 417154 292102 417774 292170
rect 417154 292046 417250 292102
rect 417306 292046 417374 292102
rect 417430 292046 417498 292102
rect 417554 292046 417622 292102
rect 417678 292046 417774 292102
rect 417154 291978 417774 292046
rect 417154 291922 417250 291978
rect 417306 291922 417374 291978
rect 417430 291922 417498 291978
rect 417554 291922 417622 291978
rect 417678 291922 417774 291978
rect 417154 274350 417774 291922
rect 417154 274294 417250 274350
rect 417306 274294 417374 274350
rect 417430 274294 417498 274350
rect 417554 274294 417622 274350
rect 417678 274294 417774 274350
rect 417154 274226 417774 274294
rect 417154 274170 417250 274226
rect 417306 274170 417374 274226
rect 417430 274170 417498 274226
rect 417554 274170 417622 274226
rect 417678 274170 417774 274226
rect 417154 274102 417774 274170
rect 417154 274046 417250 274102
rect 417306 274046 417374 274102
rect 417430 274046 417498 274102
rect 417554 274046 417622 274102
rect 417678 274046 417774 274102
rect 417154 273978 417774 274046
rect 417154 273922 417250 273978
rect 417306 273922 417374 273978
rect 417430 273922 417498 273978
rect 417554 273922 417622 273978
rect 417678 273922 417774 273978
rect 417154 256350 417774 273922
rect 417154 256294 417250 256350
rect 417306 256294 417374 256350
rect 417430 256294 417498 256350
rect 417554 256294 417622 256350
rect 417678 256294 417774 256350
rect 417154 256226 417774 256294
rect 417154 256170 417250 256226
rect 417306 256170 417374 256226
rect 417430 256170 417498 256226
rect 417554 256170 417622 256226
rect 417678 256170 417774 256226
rect 417154 256102 417774 256170
rect 417154 256046 417250 256102
rect 417306 256046 417374 256102
rect 417430 256046 417498 256102
rect 417554 256046 417622 256102
rect 417678 256046 417774 256102
rect 417154 255978 417774 256046
rect 417154 255922 417250 255978
rect 417306 255922 417374 255978
rect 417430 255922 417498 255978
rect 417554 255922 417622 255978
rect 417678 255922 417774 255978
rect 417154 238350 417774 255922
rect 417154 238294 417250 238350
rect 417306 238294 417374 238350
rect 417430 238294 417498 238350
rect 417554 238294 417622 238350
rect 417678 238294 417774 238350
rect 417154 238226 417774 238294
rect 417154 238170 417250 238226
rect 417306 238170 417374 238226
rect 417430 238170 417498 238226
rect 417554 238170 417622 238226
rect 417678 238170 417774 238226
rect 417154 238102 417774 238170
rect 417154 238046 417250 238102
rect 417306 238046 417374 238102
rect 417430 238046 417498 238102
rect 417554 238046 417622 238102
rect 417678 238046 417774 238102
rect 417154 237978 417774 238046
rect 417154 237922 417250 237978
rect 417306 237922 417374 237978
rect 417430 237922 417498 237978
rect 417554 237922 417622 237978
rect 417678 237922 417774 237978
rect 417154 220350 417774 237922
rect 417154 220294 417250 220350
rect 417306 220294 417374 220350
rect 417430 220294 417498 220350
rect 417554 220294 417622 220350
rect 417678 220294 417774 220350
rect 417154 220226 417774 220294
rect 417154 220170 417250 220226
rect 417306 220170 417374 220226
rect 417430 220170 417498 220226
rect 417554 220170 417622 220226
rect 417678 220170 417774 220226
rect 417154 220102 417774 220170
rect 417154 220046 417250 220102
rect 417306 220046 417374 220102
rect 417430 220046 417498 220102
rect 417554 220046 417622 220102
rect 417678 220046 417774 220102
rect 417154 219978 417774 220046
rect 417154 219922 417250 219978
rect 417306 219922 417374 219978
rect 417430 219922 417498 219978
rect 417554 219922 417622 219978
rect 417678 219922 417774 219978
rect 417154 217934 417774 219922
rect 420874 598172 421494 598268
rect 420874 598116 420970 598172
rect 421026 598116 421094 598172
rect 421150 598116 421218 598172
rect 421274 598116 421342 598172
rect 421398 598116 421494 598172
rect 420874 598048 421494 598116
rect 420874 597992 420970 598048
rect 421026 597992 421094 598048
rect 421150 597992 421218 598048
rect 421274 597992 421342 598048
rect 421398 597992 421494 598048
rect 420874 597924 421494 597992
rect 420874 597868 420970 597924
rect 421026 597868 421094 597924
rect 421150 597868 421218 597924
rect 421274 597868 421342 597924
rect 421398 597868 421494 597924
rect 420874 597800 421494 597868
rect 420874 597744 420970 597800
rect 421026 597744 421094 597800
rect 421150 597744 421218 597800
rect 421274 597744 421342 597800
rect 421398 597744 421494 597800
rect 420874 586350 421494 597744
rect 420874 586294 420970 586350
rect 421026 586294 421094 586350
rect 421150 586294 421218 586350
rect 421274 586294 421342 586350
rect 421398 586294 421494 586350
rect 420874 586226 421494 586294
rect 420874 586170 420970 586226
rect 421026 586170 421094 586226
rect 421150 586170 421218 586226
rect 421274 586170 421342 586226
rect 421398 586170 421494 586226
rect 420874 586102 421494 586170
rect 420874 586046 420970 586102
rect 421026 586046 421094 586102
rect 421150 586046 421218 586102
rect 421274 586046 421342 586102
rect 421398 586046 421494 586102
rect 420874 585978 421494 586046
rect 420874 585922 420970 585978
rect 421026 585922 421094 585978
rect 421150 585922 421218 585978
rect 421274 585922 421342 585978
rect 421398 585922 421494 585978
rect 420874 568350 421494 585922
rect 420874 568294 420970 568350
rect 421026 568294 421094 568350
rect 421150 568294 421218 568350
rect 421274 568294 421342 568350
rect 421398 568294 421494 568350
rect 420874 568226 421494 568294
rect 420874 568170 420970 568226
rect 421026 568170 421094 568226
rect 421150 568170 421218 568226
rect 421274 568170 421342 568226
rect 421398 568170 421494 568226
rect 420874 568102 421494 568170
rect 420874 568046 420970 568102
rect 421026 568046 421094 568102
rect 421150 568046 421218 568102
rect 421274 568046 421342 568102
rect 421398 568046 421494 568102
rect 420874 567978 421494 568046
rect 420874 567922 420970 567978
rect 421026 567922 421094 567978
rect 421150 567922 421218 567978
rect 421274 567922 421342 567978
rect 421398 567922 421494 567978
rect 420874 550350 421494 567922
rect 420874 550294 420970 550350
rect 421026 550294 421094 550350
rect 421150 550294 421218 550350
rect 421274 550294 421342 550350
rect 421398 550294 421494 550350
rect 420874 550226 421494 550294
rect 420874 550170 420970 550226
rect 421026 550170 421094 550226
rect 421150 550170 421218 550226
rect 421274 550170 421342 550226
rect 421398 550170 421494 550226
rect 420874 550102 421494 550170
rect 420874 550046 420970 550102
rect 421026 550046 421094 550102
rect 421150 550046 421218 550102
rect 421274 550046 421342 550102
rect 421398 550046 421494 550102
rect 420874 549978 421494 550046
rect 420874 549922 420970 549978
rect 421026 549922 421094 549978
rect 421150 549922 421218 549978
rect 421274 549922 421342 549978
rect 421398 549922 421494 549978
rect 420874 532350 421494 549922
rect 420874 532294 420970 532350
rect 421026 532294 421094 532350
rect 421150 532294 421218 532350
rect 421274 532294 421342 532350
rect 421398 532294 421494 532350
rect 420874 532226 421494 532294
rect 420874 532170 420970 532226
rect 421026 532170 421094 532226
rect 421150 532170 421218 532226
rect 421274 532170 421342 532226
rect 421398 532170 421494 532226
rect 420874 532102 421494 532170
rect 420874 532046 420970 532102
rect 421026 532046 421094 532102
rect 421150 532046 421218 532102
rect 421274 532046 421342 532102
rect 421398 532046 421494 532102
rect 420874 531978 421494 532046
rect 420874 531922 420970 531978
rect 421026 531922 421094 531978
rect 421150 531922 421218 531978
rect 421274 531922 421342 531978
rect 421398 531922 421494 531978
rect 420874 514350 421494 531922
rect 420874 514294 420970 514350
rect 421026 514294 421094 514350
rect 421150 514294 421218 514350
rect 421274 514294 421342 514350
rect 421398 514294 421494 514350
rect 420874 514226 421494 514294
rect 420874 514170 420970 514226
rect 421026 514170 421094 514226
rect 421150 514170 421218 514226
rect 421274 514170 421342 514226
rect 421398 514170 421494 514226
rect 420874 514102 421494 514170
rect 420874 514046 420970 514102
rect 421026 514046 421094 514102
rect 421150 514046 421218 514102
rect 421274 514046 421342 514102
rect 421398 514046 421494 514102
rect 420874 513978 421494 514046
rect 420874 513922 420970 513978
rect 421026 513922 421094 513978
rect 421150 513922 421218 513978
rect 421274 513922 421342 513978
rect 421398 513922 421494 513978
rect 420874 496350 421494 513922
rect 420874 496294 420970 496350
rect 421026 496294 421094 496350
rect 421150 496294 421218 496350
rect 421274 496294 421342 496350
rect 421398 496294 421494 496350
rect 420874 496226 421494 496294
rect 420874 496170 420970 496226
rect 421026 496170 421094 496226
rect 421150 496170 421218 496226
rect 421274 496170 421342 496226
rect 421398 496170 421494 496226
rect 420874 496102 421494 496170
rect 420874 496046 420970 496102
rect 421026 496046 421094 496102
rect 421150 496046 421218 496102
rect 421274 496046 421342 496102
rect 421398 496046 421494 496102
rect 420874 495978 421494 496046
rect 420874 495922 420970 495978
rect 421026 495922 421094 495978
rect 421150 495922 421218 495978
rect 421274 495922 421342 495978
rect 421398 495922 421494 495978
rect 420874 478350 421494 495922
rect 420874 478294 420970 478350
rect 421026 478294 421094 478350
rect 421150 478294 421218 478350
rect 421274 478294 421342 478350
rect 421398 478294 421494 478350
rect 420874 478226 421494 478294
rect 420874 478170 420970 478226
rect 421026 478170 421094 478226
rect 421150 478170 421218 478226
rect 421274 478170 421342 478226
rect 421398 478170 421494 478226
rect 420874 478102 421494 478170
rect 420874 478046 420970 478102
rect 421026 478046 421094 478102
rect 421150 478046 421218 478102
rect 421274 478046 421342 478102
rect 421398 478046 421494 478102
rect 420874 477978 421494 478046
rect 420874 477922 420970 477978
rect 421026 477922 421094 477978
rect 421150 477922 421218 477978
rect 421274 477922 421342 477978
rect 421398 477922 421494 477978
rect 420874 460350 421494 477922
rect 420874 460294 420970 460350
rect 421026 460294 421094 460350
rect 421150 460294 421218 460350
rect 421274 460294 421342 460350
rect 421398 460294 421494 460350
rect 420874 460226 421494 460294
rect 420874 460170 420970 460226
rect 421026 460170 421094 460226
rect 421150 460170 421218 460226
rect 421274 460170 421342 460226
rect 421398 460170 421494 460226
rect 420874 460102 421494 460170
rect 420874 460046 420970 460102
rect 421026 460046 421094 460102
rect 421150 460046 421218 460102
rect 421274 460046 421342 460102
rect 421398 460046 421494 460102
rect 420874 459978 421494 460046
rect 420874 459922 420970 459978
rect 421026 459922 421094 459978
rect 421150 459922 421218 459978
rect 421274 459922 421342 459978
rect 421398 459922 421494 459978
rect 420874 442350 421494 459922
rect 420874 442294 420970 442350
rect 421026 442294 421094 442350
rect 421150 442294 421218 442350
rect 421274 442294 421342 442350
rect 421398 442294 421494 442350
rect 420874 442226 421494 442294
rect 420874 442170 420970 442226
rect 421026 442170 421094 442226
rect 421150 442170 421218 442226
rect 421274 442170 421342 442226
rect 421398 442170 421494 442226
rect 420874 442102 421494 442170
rect 420874 442046 420970 442102
rect 421026 442046 421094 442102
rect 421150 442046 421218 442102
rect 421274 442046 421342 442102
rect 421398 442046 421494 442102
rect 420874 441978 421494 442046
rect 420874 441922 420970 441978
rect 421026 441922 421094 441978
rect 421150 441922 421218 441978
rect 421274 441922 421342 441978
rect 421398 441922 421494 441978
rect 420874 424350 421494 441922
rect 420874 424294 420970 424350
rect 421026 424294 421094 424350
rect 421150 424294 421218 424350
rect 421274 424294 421342 424350
rect 421398 424294 421494 424350
rect 420874 424226 421494 424294
rect 420874 424170 420970 424226
rect 421026 424170 421094 424226
rect 421150 424170 421218 424226
rect 421274 424170 421342 424226
rect 421398 424170 421494 424226
rect 420874 424102 421494 424170
rect 420874 424046 420970 424102
rect 421026 424046 421094 424102
rect 421150 424046 421218 424102
rect 421274 424046 421342 424102
rect 421398 424046 421494 424102
rect 420874 423978 421494 424046
rect 420874 423922 420970 423978
rect 421026 423922 421094 423978
rect 421150 423922 421218 423978
rect 421274 423922 421342 423978
rect 421398 423922 421494 423978
rect 420874 406350 421494 423922
rect 420874 406294 420970 406350
rect 421026 406294 421094 406350
rect 421150 406294 421218 406350
rect 421274 406294 421342 406350
rect 421398 406294 421494 406350
rect 420874 406226 421494 406294
rect 420874 406170 420970 406226
rect 421026 406170 421094 406226
rect 421150 406170 421218 406226
rect 421274 406170 421342 406226
rect 421398 406170 421494 406226
rect 420874 406102 421494 406170
rect 420874 406046 420970 406102
rect 421026 406046 421094 406102
rect 421150 406046 421218 406102
rect 421274 406046 421342 406102
rect 421398 406046 421494 406102
rect 420874 405978 421494 406046
rect 420874 405922 420970 405978
rect 421026 405922 421094 405978
rect 421150 405922 421218 405978
rect 421274 405922 421342 405978
rect 421398 405922 421494 405978
rect 420874 388350 421494 405922
rect 420874 388294 420970 388350
rect 421026 388294 421094 388350
rect 421150 388294 421218 388350
rect 421274 388294 421342 388350
rect 421398 388294 421494 388350
rect 420874 388226 421494 388294
rect 420874 388170 420970 388226
rect 421026 388170 421094 388226
rect 421150 388170 421218 388226
rect 421274 388170 421342 388226
rect 421398 388170 421494 388226
rect 420874 388102 421494 388170
rect 420874 388046 420970 388102
rect 421026 388046 421094 388102
rect 421150 388046 421218 388102
rect 421274 388046 421342 388102
rect 421398 388046 421494 388102
rect 420874 387978 421494 388046
rect 420874 387922 420970 387978
rect 421026 387922 421094 387978
rect 421150 387922 421218 387978
rect 421274 387922 421342 387978
rect 421398 387922 421494 387978
rect 420874 370350 421494 387922
rect 420874 370294 420970 370350
rect 421026 370294 421094 370350
rect 421150 370294 421218 370350
rect 421274 370294 421342 370350
rect 421398 370294 421494 370350
rect 420874 370226 421494 370294
rect 420874 370170 420970 370226
rect 421026 370170 421094 370226
rect 421150 370170 421218 370226
rect 421274 370170 421342 370226
rect 421398 370170 421494 370226
rect 420874 370102 421494 370170
rect 420874 370046 420970 370102
rect 421026 370046 421094 370102
rect 421150 370046 421218 370102
rect 421274 370046 421342 370102
rect 421398 370046 421494 370102
rect 420874 369978 421494 370046
rect 420874 369922 420970 369978
rect 421026 369922 421094 369978
rect 421150 369922 421218 369978
rect 421274 369922 421342 369978
rect 421398 369922 421494 369978
rect 420874 352350 421494 369922
rect 420874 352294 420970 352350
rect 421026 352294 421094 352350
rect 421150 352294 421218 352350
rect 421274 352294 421342 352350
rect 421398 352294 421494 352350
rect 420874 352226 421494 352294
rect 420874 352170 420970 352226
rect 421026 352170 421094 352226
rect 421150 352170 421218 352226
rect 421274 352170 421342 352226
rect 421398 352170 421494 352226
rect 420874 352102 421494 352170
rect 420874 352046 420970 352102
rect 421026 352046 421094 352102
rect 421150 352046 421218 352102
rect 421274 352046 421342 352102
rect 421398 352046 421494 352102
rect 420874 351978 421494 352046
rect 420874 351922 420970 351978
rect 421026 351922 421094 351978
rect 421150 351922 421218 351978
rect 421274 351922 421342 351978
rect 421398 351922 421494 351978
rect 420874 334350 421494 351922
rect 420874 334294 420970 334350
rect 421026 334294 421094 334350
rect 421150 334294 421218 334350
rect 421274 334294 421342 334350
rect 421398 334294 421494 334350
rect 420874 334226 421494 334294
rect 420874 334170 420970 334226
rect 421026 334170 421094 334226
rect 421150 334170 421218 334226
rect 421274 334170 421342 334226
rect 421398 334170 421494 334226
rect 420874 334102 421494 334170
rect 420874 334046 420970 334102
rect 421026 334046 421094 334102
rect 421150 334046 421218 334102
rect 421274 334046 421342 334102
rect 421398 334046 421494 334102
rect 420874 333978 421494 334046
rect 420874 333922 420970 333978
rect 421026 333922 421094 333978
rect 421150 333922 421218 333978
rect 421274 333922 421342 333978
rect 421398 333922 421494 333978
rect 420874 316350 421494 333922
rect 420874 316294 420970 316350
rect 421026 316294 421094 316350
rect 421150 316294 421218 316350
rect 421274 316294 421342 316350
rect 421398 316294 421494 316350
rect 420874 316226 421494 316294
rect 420874 316170 420970 316226
rect 421026 316170 421094 316226
rect 421150 316170 421218 316226
rect 421274 316170 421342 316226
rect 421398 316170 421494 316226
rect 420874 316102 421494 316170
rect 420874 316046 420970 316102
rect 421026 316046 421094 316102
rect 421150 316046 421218 316102
rect 421274 316046 421342 316102
rect 421398 316046 421494 316102
rect 420874 315978 421494 316046
rect 420874 315922 420970 315978
rect 421026 315922 421094 315978
rect 421150 315922 421218 315978
rect 421274 315922 421342 315978
rect 421398 315922 421494 315978
rect 420874 298350 421494 315922
rect 420874 298294 420970 298350
rect 421026 298294 421094 298350
rect 421150 298294 421218 298350
rect 421274 298294 421342 298350
rect 421398 298294 421494 298350
rect 420874 298226 421494 298294
rect 420874 298170 420970 298226
rect 421026 298170 421094 298226
rect 421150 298170 421218 298226
rect 421274 298170 421342 298226
rect 421398 298170 421494 298226
rect 420874 298102 421494 298170
rect 420874 298046 420970 298102
rect 421026 298046 421094 298102
rect 421150 298046 421218 298102
rect 421274 298046 421342 298102
rect 421398 298046 421494 298102
rect 420874 297978 421494 298046
rect 420874 297922 420970 297978
rect 421026 297922 421094 297978
rect 421150 297922 421218 297978
rect 421274 297922 421342 297978
rect 421398 297922 421494 297978
rect 420874 280350 421494 297922
rect 420874 280294 420970 280350
rect 421026 280294 421094 280350
rect 421150 280294 421218 280350
rect 421274 280294 421342 280350
rect 421398 280294 421494 280350
rect 420874 280226 421494 280294
rect 420874 280170 420970 280226
rect 421026 280170 421094 280226
rect 421150 280170 421218 280226
rect 421274 280170 421342 280226
rect 421398 280170 421494 280226
rect 420874 280102 421494 280170
rect 420874 280046 420970 280102
rect 421026 280046 421094 280102
rect 421150 280046 421218 280102
rect 421274 280046 421342 280102
rect 421398 280046 421494 280102
rect 420874 279978 421494 280046
rect 420874 279922 420970 279978
rect 421026 279922 421094 279978
rect 421150 279922 421218 279978
rect 421274 279922 421342 279978
rect 421398 279922 421494 279978
rect 420874 262350 421494 279922
rect 420874 262294 420970 262350
rect 421026 262294 421094 262350
rect 421150 262294 421218 262350
rect 421274 262294 421342 262350
rect 421398 262294 421494 262350
rect 420874 262226 421494 262294
rect 420874 262170 420970 262226
rect 421026 262170 421094 262226
rect 421150 262170 421218 262226
rect 421274 262170 421342 262226
rect 421398 262170 421494 262226
rect 420874 262102 421494 262170
rect 420874 262046 420970 262102
rect 421026 262046 421094 262102
rect 421150 262046 421218 262102
rect 421274 262046 421342 262102
rect 421398 262046 421494 262102
rect 420874 261978 421494 262046
rect 420874 261922 420970 261978
rect 421026 261922 421094 261978
rect 421150 261922 421218 261978
rect 421274 261922 421342 261978
rect 421398 261922 421494 261978
rect 420874 244350 421494 261922
rect 420874 244294 420970 244350
rect 421026 244294 421094 244350
rect 421150 244294 421218 244350
rect 421274 244294 421342 244350
rect 421398 244294 421494 244350
rect 420874 244226 421494 244294
rect 420874 244170 420970 244226
rect 421026 244170 421094 244226
rect 421150 244170 421218 244226
rect 421274 244170 421342 244226
rect 421398 244170 421494 244226
rect 420874 244102 421494 244170
rect 420874 244046 420970 244102
rect 421026 244046 421094 244102
rect 421150 244046 421218 244102
rect 421274 244046 421342 244102
rect 421398 244046 421494 244102
rect 420874 243978 421494 244046
rect 420874 243922 420970 243978
rect 421026 243922 421094 243978
rect 421150 243922 421218 243978
rect 421274 243922 421342 243978
rect 421398 243922 421494 243978
rect 420874 226350 421494 243922
rect 438874 598172 439494 598268
rect 438874 598116 438970 598172
rect 439026 598116 439094 598172
rect 439150 598116 439218 598172
rect 439274 598116 439342 598172
rect 439398 598116 439494 598172
rect 438874 598048 439494 598116
rect 438874 597992 438970 598048
rect 439026 597992 439094 598048
rect 439150 597992 439218 598048
rect 439274 597992 439342 598048
rect 439398 597992 439494 598048
rect 438874 597924 439494 597992
rect 438874 597868 438970 597924
rect 439026 597868 439094 597924
rect 439150 597868 439218 597924
rect 439274 597868 439342 597924
rect 439398 597868 439494 597924
rect 438874 597800 439494 597868
rect 438874 597744 438970 597800
rect 439026 597744 439094 597800
rect 439150 597744 439218 597800
rect 439274 597744 439342 597800
rect 439398 597744 439494 597800
rect 438874 586350 439494 597744
rect 438874 586294 438970 586350
rect 439026 586294 439094 586350
rect 439150 586294 439218 586350
rect 439274 586294 439342 586350
rect 439398 586294 439494 586350
rect 438874 586226 439494 586294
rect 438874 586170 438970 586226
rect 439026 586170 439094 586226
rect 439150 586170 439218 586226
rect 439274 586170 439342 586226
rect 439398 586170 439494 586226
rect 438874 586102 439494 586170
rect 438874 586046 438970 586102
rect 439026 586046 439094 586102
rect 439150 586046 439218 586102
rect 439274 586046 439342 586102
rect 439398 586046 439494 586102
rect 438874 585978 439494 586046
rect 438874 585922 438970 585978
rect 439026 585922 439094 585978
rect 439150 585922 439218 585978
rect 439274 585922 439342 585978
rect 439398 585922 439494 585978
rect 438874 568350 439494 585922
rect 438874 568294 438970 568350
rect 439026 568294 439094 568350
rect 439150 568294 439218 568350
rect 439274 568294 439342 568350
rect 439398 568294 439494 568350
rect 438874 568226 439494 568294
rect 438874 568170 438970 568226
rect 439026 568170 439094 568226
rect 439150 568170 439218 568226
rect 439274 568170 439342 568226
rect 439398 568170 439494 568226
rect 438874 568102 439494 568170
rect 438874 568046 438970 568102
rect 439026 568046 439094 568102
rect 439150 568046 439218 568102
rect 439274 568046 439342 568102
rect 439398 568046 439494 568102
rect 438874 567978 439494 568046
rect 438874 567922 438970 567978
rect 439026 567922 439094 567978
rect 439150 567922 439218 567978
rect 439274 567922 439342 567978
rect 439398 567922 439494 567978
rect 438874 550350 439494 567922
rect 438874 550294 438970 550350
rect 439026 550294 439094 550350
rect 439150 550294 439218 550350
rect 439274 550294 439342 550350
rect 439398 550294 439494 550350
rect 438874 550226 439494 550294
rect 438874 550170 438970 550226
rect 439026 550170 439094 550226
rect 439150 550170 439218 550226
rect 439274 550170 439342 550226
rect 439398 550170 439494 550226
rect 438874 550102 439494 550170
rect 438874 550046 438970 550102
rect 439026 550046 439094 550102
rect 439150 550046 439218 550102
rect 439274 550046 439342 550102
rect 439398 550046 439494 550102
rect 438874 549978 439494 550046
rect 438874 549922 438970 549978
rect 439026 549922 439094 549978
rect 439150 549922 439218 549978
rect 439274 549922 439342 549978
rect 439398 549922 439494 549978
rect 438874 532350 439494 549922
rect 438874 532294 438970 532350
rect 439026 532294 439094 532350
rect 439150 532294 439218 532350
rect 439274 532294 439342 532350
rect 439398 532294 439494 532350
rect 438874 532226 439494 532294
rect 438874 532170 438970 532226
rect 439026 532170 439094 532226
rect 439150 532170 439218 532226
rect 439274 532170 439342 532226
rect 439398 532170 439494 532226
rect 438874 532102 439494 532170
rect 438874 532046 438970 532102
rect 439026 532046 439094 532102
rect 439150 532046 439218 532102
rect 439274 532046 439342 532102
rect 439398 532046 439494 532102
rect 438874 531978 439494 532046
rect 438874 531922 438970 531978
rect 439026 531922 439094 531978
rect 439150 531922 439218 531978
rect 439274 531922 439342 531978
rect 439398 531922 439494 531978
rect 438874 514350 439494 531922
rect 438874 514294 438970 514350
rect 439026 514294 439094 514350
rect 439150 514294 439218 514350
rect 439274 514294 439342 514350
rect 439398 514294 439494 514350
rect 438874 514226 439494 514294
rect 438874 514170 438970 514226
rect 439026 514170 439094 514226
rect 439150 514170 439218 514226
rect 439274 514170 439342 514226
rect 439398 514170 439494 514226
rect 438874 514102 439494 514170
rect 438874 514046 438970 514102
rect 439026 514046 439094 514102
rect 439150 514046 439218 514102
rect 439274 514046 439342 514102
rect 439398 514046 439494 514102
rect 438874 513978 439494 514046
rect 438874 513922 438970 513978
rect 439026 513922 439094 513978
rect 439150 513922 439218 513978
rect 439274 513922 439342 513978
rect 439398 513922 439494 513978
rect 438874 496350 439494 513922
rect 438874 496294 438970 496350
rect 439026 496294 439094 496350
rect 439150 496294 439218 496350
rect 439274 496294 439342 496350
rect 439398 496294 439494 496350
rect 438874 496226 439494 496294
rect 438874 496170 438970 496226
rect 439026 496170 439094 496226
rect 439150 496170 439218 496226
rect 439274 496170 439342 496226
rect 439398 496170 439494 496226
rect 438874 496102 439494 496170
rect 438874 496046 438970 496102
rect 439026 496046 439094 496102
rect 439150 496046 439218 496102
rect 439274 496046 439342 496102
rect 439398 496046 439494 496102
rect 438874 495978 439494 496046
rect 438874 495922 438970 495978
rect 439026 495922 439094 495978
rect 439150 495922 439218 495978
rect 439274 495922 439342 495978
rect 439398 495922 439494 495978
rect 438874 478350 439494 495922
rect 438874 478294 438970 478350
rect 439026 478294 439094 478350
rect 439150 478294 439218 478350
rect 439274 478294 439342 478350
rect 439398 478294 439494 478350
rect 438874 478226 439494 478294
rect 438874 478170 438970 478226
rect 439026 478170 439094 478226
rect 439150 478170 439218 478226
rect 439274 478170 439342 478226
rect 439398 478170 439494 478226
rect 438874 478102 439494 478170
rect 438874 478046 438970 478102
rect 439026 478046 439094 478102
rect 439150 478046 439218 478102
rect 439274 478046 439342 478102
rect 439398 478046 439494 478102
rect 438874 477978 439494 478046
rect 438874 477922 438970 477978
rect 439026 477922 439094 477978
rect 439150 477922 439218 477978
rect 439274 477922 439342 477978
rect 439398 477922 439494 477978
rect 438874 460350 439494 477922
rect 438874 460294 438970 460350
rect 439026 460294 439094 460350
rect 439150 460294 439218 460350
rect 439274 460294 439342 460350
rect 439398 460294 439494 460350
rect 438874 460226 439494 460294
rect 438874 460170 438970 460226
rect 439026 460170 439094 460226
rect 439150 460170 439218 460226
rect 439274 460170 439342 460226
rect 439398 460170 439494 460226
rect 438874 460102 439494 460170
rect 438874 460046 438970 460102
rect 439026 460046 439094 460102
rect 439150 460046 439218 460102
rect 439274 460046 439342 460102
rect 439398 460046 439494 460102
rect 438874 459978 439494 460046
rect 438874 459922 438970 459978
rect 439026 459922 439094 459978
rect 439150 459922 439218 459978
rect 439274 459922 439342 459978
rect 439398 459922 439494 459978
rect 438874 442350 439494 459922
rect 438874 442294 438970 442350
rect 439026 442294 439094 442350
rect 439150 442294 439218 442350
rect 439274 442294 439342 442350
rect 439398 442294 439494 442350
rect 438874 442226 439494 442294
rect 438874 442170 438970 442226
rect 439026 442170 439094 442226
rect 439150 442170 439218 442226
rect 439274 442170 439342 442226
rect 439398 442170 439494 442226
rect 438874 442102 439494 442170
rect 438874 442046 438970 442102
rect 439026 442046 439094 442102
rect 439150 442046 439218 442102
rect 439274 442046 439342 442102
rect 439398 442046 439494 442102
rect 438874 441978 439494 442046
rect 438874 441922 438970 441978
rect 439026 441922 439094 441978
rect 439150 441922 439218 441978
rect 439274 441922 439342 441978
rect 439398 441922 439494 441978
rect 438874 424350 439494 441922
rect 438874 424294 438970 424350
rect 439026 424294 439094 424350
rect 439150 424294 439218 424350
rect 439274 424294 439342 424350
rect 439398 424294 439494 424350
rect 438874 424226 439494 424294
rect 438874 424170 438970 424226
rect 439026 424170 439094 424226
rect 439150 424170 439218 424226
rect 439274 424170 439342 424226
rect 439398 424170 439494 424226
rect 438874 424102 439494 424170
rect 438874 424046 438970 424102
rect 439026 424046 439094 424102
rect 439150 424046 439218 424102
rect 439274 424046 439342 424102
rect 439398 424046 439494 424102
rect 438874 423978 439494 424046
rect 438874 423922 438970 423978
rect 439026 423922 439094 423978
rect 439150 423922 439218 423978
rect 439274 423922 439342 423978
rect 439398 423922 439494 423978
rect 438874 406350 439494 423922
rect 438874 406294 438970 406350
rect 439026 406294 439094 406350
rect 439150 406294 439218 406350
rect 439274 406294 439342 406350
rect 439398 406294 439494 406350
rect 438874 406226 439494 406294
rect 438874 406170 438970 406226
rect 439026 406170 439094 406226
rect 439150 406170 439218 406226
rect 439274 406170 439342 406226
rect 439398 406170 439494 406226
rect 438874 406102 439494 406170
rect 438874 406046 438970 406102
rect 439026 406046 439094 406102
rect 439150 406046 439218 406102
rect 439274 406046 439342 406102
rect 439398 406046 439494 406102
rect 438874 405978 439494 406046
rect 438874 405922 438970 405978
rect 439026 405922 439094 405978
rect 439150 405922 439218 405978
rect 439274 405922 439342 405978
rect 439398 405922 439494 405978
rect 438874 388350 439494 405922
rect 438874 388294 438970 388350
rect 439026 388294 439094 388350
rect 439150 388294 439218 388350
rect 439274 388294 439342 388350
rect 439398 388294 439494 388350
rect 438874 388226 439494 388294
rect 438874 388170 438970 388226
rect 439026 388170 439094 388226
rect 439150 388170 439218 388226
rect 439274 388170 439342 388226
rect 439398 388170 439494 388226
rect 438874 388102 439494 388170
rect 438874 388046 438970 388102
rect 439026 388046 439094 388102
rect 439150 388046 439218 388102
rect 439274 388046 439342 388102
rect 439398 388046 439494 388102
rect 438874 387978 439494 388046
rect 438874 387922 438970 387978
rect 439026 387922 439094 387978
rect 439150 387922 439218 387978
rect 439274 387922 439342 387978
rect 439398 387922 439494 387978
rect 438874 370350 439494 387922
rect 438874 370294 438970 370350
rect 439026 370294 439094 370350
rect 439150 370294 439218 370350
rect 439274 370294 439342 370350
rect 439398 370294 439494 370350
rect 438874 370226 439494 370294
rect 438874 370170 438970 370226
rect 439026 370170 439094 370226
rect 439150 370170 439218 370226
rect 439274 370170 439342 370226
rect 439398 370170 439494 370226
rect 438874 370102 439494 370170
rect 438874 370046 438970 370102
rect 439026 370046 439094 370102
rect 439150 370046 439218 370102
rect 439274 370046 439342 370102
rect 439398 370046 439494 370102
rect 438874 369978 439494 370046
rect 438874 369922 438970 369978
rect 439026 369922 439094 369978
rect 439150 369922 439218 369978
rect 439274 369922 439342 369978
rect 439398 369922 439494 369978
rect 438874 352350 439494 369922
rect 438874 352294 438970 352350
rect 439026 352294 439094 352350
rect 439150 352294 439218 352350
rect 439274 352294 439342 352350
rect 439398 352294 439494 352350
rect 438874 352226 439494 352294
rect 438874 352170 438970 352226
rect 439026 352170 439094 352226
rect 439150 352170 439218 352226
rect 439274 352170 439342 352226
rect 439398 352170 439494 352226
rect 438874 352102 439494 352170
rect 438874 352046 438970 352102
rect 439026 352046 439094 352102
rect 439150 352046 439218 352102
rect 439274 352046 439342 352102
rect 439398 352046 439494 352102
rect 438874 351978 439494 352046
rect 438874 351922 438970 351978
rect 439026 351922 439094 351978
rect 439150 351922 439218 351978
rect 439274 351922 439342 351978
rect 439398 351922 439494 351978
rect 438874 334350 439494 351922
rect 438874 334294 438970 334350
rect 439026 334294 439094 334350
rect 439150 334294 439218 334350
rect 439274 334294 439342 334350
rect 439398 334294 439494 334350
rect 438874 334226 439494 334294
rect 438874 334170 438970 334226
rect 439026 334170 439094 334226
rect 439150 334170 439218 334226
rect 439274 334170 439342 334226
rect 439398 334170 439494 334226
rect 438874 334102 439494 334170
rect 438874 334046 438970 334102
rect 439026 334046 439094 334102
rect 439150 334046 439218 334102
rect 439274 334046 439342 334102
rect 439398 334046 439494 334102
rect 438874 333978 439494 334046
rect 438874 333922 438970 333978
rect 439026 333922 439094 333978
rect 439150 333922 439218 333978
rect 439274 333922 439342 333978
rect 439398 333922 439494 333978
rect 438874 316350 439494 333922
rect 438874 316294 438970 316350
rect 439026 316294 439094 316350
rect 439150 316294 439218 316350
rect 439274 316294 439342 316350
rect 439398 316294 439494 316350
rect 438874 316226 439494 316294
rect 438874 316170 438970 316226
rect 439026 316170 439094 316226
rect 439150 316170 439218 316226
rect 439274 316170 439342 316226
rect 439398 316170 439494 316226
rect 438874 316102 439494 316170
rect 438874 316046 438970 316102
rect 439026 316046 439094 316102
rect 439150 316046 439218 316102
rect 439274 316046 439342 316102
rect 439398 316046 439494 316102
rect 438874 315978 439494 316046
rect 438874 315922 438970 315978
rect 439026 315922 439094 315978
rect 439150 315922 439218 315978
rect 439274 315922 439342 315978
rect 439398 315922 439494 315978
rect 438874 298350 439494 315922
rect 438874 298294 438970 298350
rect 439026 298294 439094 298350
rect 439150 298294 439218 298350
rect 439274 298294 439342 298350
rect 439398 298294 439494 298350
rect 438874 298226 439494 298294
rect 438874 298170 438970 298226
rect 439026 298170 439094 298226
rect 439150 298170 439218 298226
rect 439274 298170 439342 298226
rect 439398 298170 439494 298226
rect 438874 298102 439494 298170
rect 438874 298046 438970 298102
rect 439026 298046 439094 298102
rect 439150 298046 439218 298102
rect 439274 298046 439342 298102
rect 439398 298046 439494 298102
rect 438874 297978 439494 298046
rect 438874 297922 438970 297978
rect 439026 297922 439094 297978
rect 439150 297922 439218 297978
rect 439274 297922 439342 297978
rect 439398 297922 439494 297978
rect 438874 280350 439494 297922
rect 438874 280294 438970 280350
rect 439026 280294 439094 280350
rect 439150 280294 439218 280350
rect 439274 280294 439342 280350
rect 439398 280294 439494 280350
rect 438874 280226 439494 280294
rect 438874 280170 438970 280226
rect 439026 280170 439094 280226
rect 439150 280170 439218 280226
rect 439274 280170 439342 280226
rect 439398 280170 439494 280226
rect 438874 280102 439494 280170
rect 438874 280046 438970 280102
rect 439026 280046 439094 280102
rect 439150 280046 439218 280102
rect 439274 280046 439342 280102
rect 439398 280046 439494 280102
rect 438874 279978 439494 280046
rect 438874 279922 438970 279978
rect 439026 279922 439094 279978
rect 439150 279922 439218 279978
rect 439274 279922 439342 279978
rect 439398 279922 439494 279978
rect 438874 262350 439494 279922
rect 438874 262294 438970 262350
rect 439026 262294 439094 262350
rect 439150 262294 439218 262350
rect 439274 262294 439342 262350
rect 439398 262294 439494 262350
rect 438874 262226 439494 262294
rect 438874 262170 438970 262226
rect 439026 262170 439094 262226
rect 439150 262170 439218 262226
rect 439274 262170 439342 262226
rect 439398 262170 439494 262226
rect 438874 262102 439494 262170
rect 438874 262046 438970 262102
rect 439026 262046 439094 262102
rect 439150 262046 439218 262102
rect 439274 262046 439342 262102
rect 439398 262046 439494 262102
rect 438874 261978 439494 262046
rect 438874 261922 438970 261978
rect 439026 261922 439094 261978
rect 439150 261922 439218 261978
rect 439274 261922 439342 261978
rect 439398 261922 439494 261978
rect 438874 244350 439494 261922
rect 438874 244294 438970 244350
rect 439026 244294 439094 244350
rect 439150 244294 439218 244350
rect 439274 244294 439342 244350
rect 439398 244294 439494 244350
rect 438874 244226 439494 244294
rect 438874 244170 438970 244226
rect 439026 244170 439094 244226
rect 439150 244170 439218 244226
rect 439274 244170 439342 244226
rect 439398 244170 439494 244226
rect 438874 244102 439494 244170
rect 438874 244046 438970 244102
rect 439026 244046 439094 244102
rect 439150 244046 439218 244102
rect 439274 244046 439342 244102
rect 439398 244046 439494 244102
rect 438874 243978 439494 244046
rect 438874 243922 438970 243978
rect 439026 243922 439094 243978
rect 439150 243922 439218 243978
rect 439274 243922 439342 243978
rect 439398 243922 439494 243978
rect 420874 226294 420970 226350
rect 421026 226294 421094 226350
rect 421150 226294 421218 226350
rect 421274 226294 421342 226350
rect 421398 226294 421494 226350
rect 420874 226226 421494 226294
rect 420874 226170 420970 226226
rect 421026 226170 421094 226226
rect 421150 226170 421218 226226
rect 421274 226170 421342 226226
rect 421398 226170 421494 226226
rect 420874 226102 421494 226170
rect 420874 226046 420970 226102
rect 421026 226046 421094 226102
rect 421150 226046 421218 226102
rect 421274 226046 421342 226102
rect 421398 226046 421494 226102
rect 420874 225978 421494 226046
rect 420874 225922 420970 225978
rect 421026 225922 421094 225978
rect 421150 225922 421218 225978
rect 421274 225922 421342 225978
rect 421398 225922 421494 225978
rect 420874 217934 421494 225922
rect 435154 238350 435774 242964
rect 435154 238294 435250 238350
rect 435306 238294 435374 238350
rect 435430 238294 435498 238350
rect 435554 238294 435622 238350
rect 435678 238294 435774 238350
rect 435154 238226 435774 238294
rect 435154 238170 435250 238226
rect 435306 238170 435374 238226
rect 435430 238170 435498 238226
rect 435554 238170 435622 238226
rect 435678 238170 435774 238226
rect 435154 238102 435774 238170
rect 435154 238046 435250 238102
rect 435306 238046 435374 238102
rect 435430 238046 435498 238102
rect 435554 238046 435622 238102
rect 435678 238046 435774 238102
rect 435154 237978 435774 238046
rect 435154 237922 435250 237978
rect 435306 237922 435374 237978
rect 435430 237922 435498 237978
rect 435554 237922 435622 237978
rect 435678 237922 435774 237978
rect 435154 220350 435774 237922
rect 435154 220294 435250 220350
rect 435306 220294 435374 220350
rect 435430 220294 435498 220350
rect 435554 220294 435622 220350
rect 435678 220294 435774 220350
rect 435154 220226 435774 220294
rect 435154 220170 435250 220226
rect 435306 220170 435374 220226
rect 435430 220170 435498 220226
rect 435554 220170 435622 220226
rect 435678 220170 435774 220226
rect 435154 220102 435774 220170
rect 435154 220046 435250 220102
rect 435306 220046 435374 220102
rect 435430 220046 435498 220102
rect 435554 220046 435622 220102
rect 435678 220046 435774 220102
rect 435154 219978 435774 220046
rect 435154 219922 435250 219978
rect 435306 219922 435374 219978
rect 435430 219922 435498 219978
rect 435554 219922 435622 219978
rect 435678 219922 435774 219978
rect 435154 218572 435774 219922
rect 438874 226350 439494 243922
rect 438874 226294 438970 226350
rect 439026 226294 439094 226350
rect 439150 226294 439218 226350
rect 439274 226294 439342 226350
rect 439398 226294 439494 226350
rect 438874 226226 439494 226294
rect 438874 226170 438970 226226
rect 439026 226170 439094 226226
rect 439150 226170 439218 226226
rect 439274 226170 439342 226226
rect 439398 226170 439494 226226
rect 438874 226102 439494 226170
rect 438874 226046 438970 226102
rect 439026 226046 439094 226102
rect 439150 226046 439218 226102
rect 439274 226046 439342 226102
rect 439398 226046 439494 226102
rect 438874 225978 439494 226046
rect 438874 225922 438970 225978
rect 439026 225922 439094 225978
rect 439150 225922 439218 225978
rect 439274 225922 439342 225978
rect 439398 225922 439494 225978
rect 438874 217934 439494 225922
rect 453154 597212 453774 598268
rect 453154 597156 453250 597212
rect 453306 597156 453374 597212
rect 453430 597156 453498 597212
rect 453554 597156 453622 597212
rect 453678 597156 453774 597212
rect 453154 597088 453774 597156
rect 453154 597032 453250 597088
rect 453306 597032 453374 597088
rect 453430 597032 453498 597088
rect 453554 597032 453622 597088
rect 453678 597032 453774 597088
rect 453154 596964 453774 597032
rect 453154 596908 453250 596964
rect 453306 596908 453374 596964
rect 453430 596908 453498 596964
rect 453554 596908 453622 596964
rect 453678 596908 453774 596964
rect 453154 596840 453774 596908
rect 453154 596784 453250 596840
rect 453306 596784 453374 596840
rect 453430 596784 453498 596840
rect 453554 596784 453622 596840
rect 453678 596784 453774 596840
rect 453154 580350 453774 596784
rect 453154 580294 453250 580350
rect 453306 580294 453374 580350
rect 453430 580294 453498 580350
rect 453554 580294 453622 580350
rect 453678 580294 453774 580350
rect 453154 580226 453774 580294
rect 453154 580170 453250 580226
rect 453306 580170 453374 580226
rect 453430 580170 453498 580226
rect 453554 580170 453622 580226
rect 453678 580170 453774 580226
rect 453154 580102 453774 580170
rect 453154 580046 453250 580102
rect 453306 580046 453374 580102
rect 453430 580046 453498 580102
rect 453554 580046 453622 580102
rect 453678 580046 453774 580102
rect 453154 579978 453774 580046
rect 453154 579922 453250 579978
rect 453306 579922 453374 579978
rect 453430 579922 453498 579978
rect 453554 579922 453622 579978
rect 453678 579922 453774 579978
rect 453154 562350 453774 579922
rect 453154 562294 453250 562350
rect 453306 562294 453374 562350
rect 453430 562294 453498 562350
rect 453554 562294 453622 562350
rect 453678 562294 453774 562350
rect 453154 562226 453774 562294
rect 453154 562170 453250 562226
rect 453306 562170 453374 562226
rect 453430 562170 453498 562226
rect 453554 562170 453622 562226
rect 453678 562170 453774 562226
rect 453154 562102 453774 562170
rect 453154 562046 453250 562102
rect 453306 562046 453374 562102
rect 453430 562046 453498 562102
rect 453554 562046 453622 562102
rect 453678 562046 453774 562102
rect 453154 561978 453774 562046
rect 453154 561922 453250 561978
rect 453306 561922 453374 561978
rect 453430 561922 453498 561978
rect 453554 561922 453622 561978
rect 453678 561922 453774 561978
rect 453154 544350 453774 561922
rect 453154 544294 453250 544350
rect 453306 544294 453374 544350
rect 453430 544294 453498 544350
rect 453554 544294 453622 544350
rect 453678 544294 453774 544350
rect 453154 544226 453774 544294
rect 453154 544170 453250 544226
rect 453306 544170 453374 544226
rect 453430 544170 453498 544226
rect 453554 544170 453622 544226
rect 453678 544170 453774 544226
rect 453154 544102 453774 544170
rect 453154 544046 453250 544102
rect 453306 544046 453374 544102
rect 453430 544046 453498 544102
rect 453554 544046 453622 544102
rect 453678 544046 453774 544102
rect 453154 543978 453774 544046
rect 453154 543922 453250 543978
rect 453306 543922 453374 543978
rect 453430 543922 453498 543978
rect 453554 543922 453622 543978
rect 453678 543922 453774 543978
rect 453154 526350 453774 543922
rect 453154 526294 453250 526350
rect 453306 526294 453374 526350
rect 453430 526294 453498 526350
rect 453554 526294 453622 526350
rect 453678 526294 453774 526350
rect 453154 526226 453774 526294
rect 453154 526170 453250 526226
rect 453306 526170 453374 526226
rect 453430 526170 453498 526226
rect 453554 526170 453622 526226
rect 453678 526170 453774 526226
rect 453154 526102 453774 526170
rect 453154 526046 453250 526102
rect 453306 526046 453374 526102
rect 453430 526046 453498 526102
rect 453554 526046 453622 526102
rect 453678 526046 453774 526102
rect 453154 525978 453774 526046
rect 453154 525922 453250 525978
rect 453306 525922 453374 525978
rect 453430 525922 453498 525978
rect 453554 525922 453622 525978
rect 453678 525922 453774 525978
rect 453154 508350 453774 525922
rect 453154 508294 453250 508350
rect 453306 508294 453374 508350
rect 453430 508294 453498 508350
rect 453554 508294 453622 508350
rect 453678 508294 453774 508350
rect 453154 508226 453774 508294
rect 453154 508170 453250 508226
rect 453306 508170 453374 508226
rect 453430 508170 453498 508226
rect 453554 508170 453622 508226
rect 453678 508170 453774 508226
rect 453154 508102 453774 508170
rect 453154 508046 453250 508102
rect 453306 508046 453374 508102
rect 453430 508046 453498 508102
rect 453554 508046 453622 508102
rect 453678 508046 453774 508102
rect 453154 507978 453774 508046
rect 453154 507922 453250 507978
rect 453306 507922 453374 507978
rect 453430 507922 453498 507978
rect 453554 507922 453622 507978
rect 453678 507922 453774 507978
rect 453154 490350 453774 507922
rect 453154 490294 453250 490350
rect 453306 490294 453374 490350
rect 453430 490294 453498 490350
rect 453554 490294 453622 490350
rect 453678 490294 453774 490350
rect 453154 490226 453774 490294
rect 453154 490170 453250 490226
rect 453306 490170 453374 490226
rect 453430 490170 453498 490226
rect 453554 490170 453622 490226
rect 453678 490170 453774 490226
rect 453154 490102 453774 490170
rect 453154 490046 453250 490102
rect 453306 490046 453374 490102
rect 453430 490046 453498 490102
rect 453554 490046 453622 490102
rect 453678 490046 453774 490102
rect 453154 489978 453774 490046
rect 453154 489922 453250 489978
rect 453306 489922 453374 489978
rect 453430 489922 453498 489978
rect 453554 489922 453622 489978
rect 453678 489922 453774 489978
rect 453154 472350 453774 489922
rect 453154 472294 453250 472350
rect 453306 472294 453374 472350
rect 453430 472294 453498 472350
rect 453554 472294 453622 472350
rect 453678 472294 453774 472350
rect 453154 472226 453774 472294
rect 453154 472170 453250 472226
rect 453306 472170 453374 472226
rect 453430 472170 453498 472226
rect 453554 472170 453622 472226
rect 453678 472170 453774 472226
rect 453154 472102 453774 472170
rect 453154 472046 453250 472102
rect 453306 472046 453374 472102
rect 453430 472046 453498 472102
rect 453554 472046 453622 472102
rect 453678 472046 453774 472102
rect 453154 471978 453774 472046
rect 453154 471922 453250 471978
rect 453306 471922 453374 471978
rect 453430 471922 453498 471978
rect 453554 471922 453622 471978
rect 453678 471922 453774 471978
rect 453154 454350 453774 471922
rect 453154 454294 453250 454350
rect 453306 454294 453374 454350
rect 453430 454294 453498 454350
rect 453554 454294 453622 454350
rect 453678 454294 453774 454350
rect 453154 454226 453774 454294
rect 453154 454170 453250 454226
rect 453306 454170 453374 454226
rect 453430 454170 453498 454226
rect 453554 454170 453622 454226
rect 453678 454170 453774 454226
rect 453154 454102 453774 454170
rect 453154 454046 453250 454102
rect 453306 454046 453374 454102
rect 453430 454046 453498 454102
rect 453554 454046 453622 454102
rect 453678 454046 453774 454102
rect 453154 453978 453774 454046
rect 453154 453922 453250 453978
rect 453306 453922 453374 453978
rect 453430 453922 453498 453978
rect 453554 453922 453622 453978
rect 453678 453922 453774 453978
rect 453154 436350 453774 453922
rect 453154 436294 453250 436350
rect 453306 436294 453374 436350
rect 453430 436294 453498 436350
rect 453554 436294 453622 436350
rect 453678 436294 453774 436350
rect 453154 436226 453774 436294
rect 453154 436170 453250 436226
rect 453306 436170 453374 436226
rect 453430 436170 453498 436226
rect 453554 436170 453622 436226
rect 453678 436170 453774 436226
rect 453154 436102 453774 436170
rect 453154 436046 453250 436102
rect 453306 436046 453374 436102
rect 453430 436046 453498 436102
rect 453554 436046 453622 436102
rect 453678 436046 453774 436102
rect 453154 435978 453774 436046
rect 453154 435922 453250 435978
rect 453306 435922 453374 435978
rect 453430 435922 453498 435978
rect 453554 435922 453622 435978
rect 453678 435922 453774 435978
rect 453154 418350 453774 435922
rect 453154 418294 453250 418350
rect 453306 418294 453374 418350
rect 453430 418294 453498 418350
rect 453554 418294 453622 418350
rect 453678 418294 453774 418350
rect 453154 418226 453774 418294
rect 453154 418170 453250 418226
rect 453306 418170 453374 418226
rect 453430 418170 453498 418226
rect 453554 418170 453622 418226
rect 453678 418170 453774 418226
rect 453154 418102 453774 418170
rect 453154 418046 453250 418102
rect 453306 418046 453374 418102
rect 453430 418046 453498 418102
rect 453554 418046 453622 418102
rect 453678 418046 453774 418102
rect 453154 417978 453774 418046
rect 453154 417922 453250 417978
rect 453306 417922 453374 417978
rect 453430 417922 453498 417978
rect 453554 417922 453622 417978
rect 453678 417922 453774 417978
rect 453154 400350 453774 417922
rect 453154 400294 453250 400350
rect 453306 400294 453374 400350
rect 453430 400294 453498 400350
rect 453554 400294 453622 400350
rect 453678 400294 453774 400350
rect 453154 400226 453774 400294
rect 453154 400170 453250 400226
rect 453306 400170 453374 400226
rect 453430 400170 453498 400226
rect 453554 400170 453622 400226
rect 453678 400170 453774 400226
rect 453154 400102 453774 400170
rect 453154 400046 453250 400102
rect 453306 400046 453374 400102
rect 453430 400046 453498 400102
rect 453554 400046 453622 400102
rect 453678 400046 453774 400102
rect 453154 399978 453774 400046
rect 453154 399922 453250 399978
rect 453306 399922 453374 399978
rect 453430 399922 453498 399978
rect 453554 399922 453622 399978
rect 453678 399922 453774 399978
rect 453154 382350 453774 399922
rect 453154 382294 453250 382350
rect 453306 382294 453374 382350
rect 453430 382294 453498 382350
rect 453554 382294 453622 382350
rect 453678 382294 453774 382350
rect 453154 382226 453774 382294
rect 453154 382170 453250 382226
rect 453306 382170 453374 382226
rect 453430 382170 453498 382226
rect 453554 382170 453622 382226
rect 453678 382170 453774 382226
rect 453154 382102 453774 382170
rect 453154 382046 453250 382102
rect 453306 382046 453374 382102
rect 453430 382046 453498 382102
rect 453554 382046 453622 382102
rect 453678 382046 453774 382102
rect 453154 381978 453774 382046
rect 453154 381922 453250 381978
rect 453306 381922 453374 381978
rect 453430 381922 453498 381978
rect 453554 381922 453622 381978
rect 453678 381922 453774 381978
rect 453154 364350 453774 381922
rect 453154 364294 453250 364350
rect 453306 364294 453374 364350
rect 453430 364294 453498 364350
rect 453554 364294 453622 364350
rect 453678 364294 453774 364350
rect 453154 364226 453774 364294
rect 453154 364170 453250 364226
rect 453306 364170 453374 364226
rect 453430 364170 453498 364226
rect 453554 364170 453622 364226
rect 453678 364170 453774 364226
rect 453154 364102 453774 364170
rect 453154 364046 453250 364102
rect 453306 364046 453374 364102
rect 453430 364046 453498 364102
rect 453554 364046 453622 364102
rect 453678 364046 453774 364102
rect 453154 363978 453774 364046
rect 453154 363922 453250 363978
rect 453306 363922 453374 363978
rect 453430 363922 453498 363978
rect 453554 363922 453622 363978
rect 453678 363922 453774 363978
rect 453154 346350 453774 363922
rect 453154 346294 453250 346350
rect 453306 346294 453374 346350
rect 453430 346294 453498 346350
rect 453554 346294 453622 346350
rect 453678 346294 453774 346350
rect 453154 346226 453774 346294
rect 453154 346170 453250 346226
rect 453306 346170 453374 346226
rect 453430 346170 453498 346226
rect 453554 346170 453622 346226
rect 453678 346170 453774 346226
rect 453154 346102 453774 346170
rect 453154 346046 453250 346102
rect 453306 346046 453374 346102
rect 453430 346046 453498 346102
rect 453554 346046 453622 346102
rect 453678 346046 453774 346102
rect 453154 345978 453774 346046
rect 453154 345922 453250 345978
rect 453306 345922 453374 345978
rect 453430 345922 453498 345978
rect 453554 345922 453622 345978
rect 453678 345922 453774 345978
rect 453154 328350 453774 345922
rect 453154 328294 453250 328350
rect 453306 328294 453374 328350
rect 453430 328294 453498 328350
rect 453554 328294 453622 328350
rect 453678 328294 453774 328350
rect 453154 328226 453774 328294
rect 453154 328170 453250 328226
rect 453306 328170 453374 328226
rect 453430 328170 453498 328226
rect 453554 328170 453622 328226
rect 453678 328170 453774 328226
rect 453154 328102 453774 328170
rect 453154 328046 453250 328102
rect 453306 328046 453374 328102
rect 453430 328046 453498 328102
rect 453554 328046 453622 328102
rect 453678 328046 453774 328102
rect 453154 327978 453774 328046
rect 453154 327922 453250 327978
rect 453306 327922 453374 327978
rect 453430 327922 453498 327978
rect 453554 327922 453622 327978
rect 453678 327922 453774 327978
rect 453154 310350 453774 327922
rect 453154 310294 453250 310350
rect 453306 310294 453374 310350
rect 453430 310294 453498 310350
rect 453554 310294 453622 310350
rect 453678 310294 453774 310350
rect 453154 310226 453774 310294
rect 453154 310170 453250 310226
rect 453306 310170 453374 310226
rect 453430 310170 453498 310226
rect 453554 310170 453622 310226
rect 453678 310170 453774 310226
rect 453154 310102 453774 310170
rect 453154 310046 453250 310102
rect 453306 310046 453374 310102
rect 453430 310046 453498 310102
rect 453554 310046 453622 310102
rect 453678 310046 453774 310102
rect 453154 309978 453774 310046
rect 453154 309922 453250 309978
rect 453306 309922 453374 309978
rect 453430 309922 453498 309978
rect 453554 309922 453622 309978
rect 453678 309922 453774 309978
rect 453154 292350 453774 309922
rect 453154 292294 453250 292350
rect 453306 292294 453374 292350
rect 453430 292294 453498 292350
rect 453554 292294 453622 292350
rect 453678 292294 453774 292350
rect 453154 292226 453774 292294
rect 453154 292170 453250 292226
rect 453306 292170 453374 292226
rect 453430 292170 453498 292226
rect 453554 292170 453622 292226
rect 453678 292170 453774 292226
rect 453154 292102 453774 292170
rect 453154 292046 453250 292102
rect 453306 292046 453374 292102
rect 453430 292046 453498 292102
rect 453554 292046 453622 292102
rect 453678 292046 453774 292102
rect 453154 291978 453774 292046
rect 453154 291922 453250 291978
rect 453306 291922 453374 291978
rect 453430 291922 453498 291978
rect 453554 291922 453622 291978
rect 453678 291922 453774 291978
rect 453154 274350 453774 291922
rect 453154 274294 453250 274350
rect 453306 274294 453374 274350
rect 453430 274294 453498 274350
rect 453554 274294 453622 274350
rect 453678 274294 453774 274350
rect 453154 274226 453774 274294
rect 453154 274170 453250 274226
rect 453306 274170 453374 274226
rect 453430 274170 453498 274226
rect 453554 274170 453622 274226
rect 453678 274170 453774 274226
rect 453154 274102 453774 274170
rect 453154 274046 453250 274102
rect 453306 274046 453374 274102
rect 453430 274046 453498 274102
rect 453554 274046 453622 274102
rect 453678 274046 453774 274102
rect 453154 273978 453774 274046
rect 453154 273922 453250 273978
rect 453306 273922 453374 273978
rect 453430 273922 453498 273978
rect 453554 273922 453622 273978
rect 453678 273922 453774 273978
rect 453154 256350 453774 273922
rect 453154 256294 453250 256350
rect 453306 256294 453374 256350
rect 453430 256294 453498 256350
rect 453554 256294 453622 256350
rect 453678 256294 453774 256350
rect 453154 256226 453774 256294
rect 453154 256170 453250 256226
rect 453306 256170 453374 256226
rect 453430 256170 453498 256226
rect 453554 256170 453622 256226
rect 453678 256170 453774 256226
rect 453154 256102 453774 256170
rect 453154 256046 453250 256102
rect 453306 256046 453374 256102
rect 453430 256046 453498 256102
rect 453554 256046 453622 256102
rect 453678 256046 453774 256102
rect 453154 255978 453774 256046
rect 453154 255922 453250 255978
rect 453306 255922 453374 255978
rect 453430 255922 453498 255978
rect 453554 255922 453622 255978
rect 453678 255922 453774 255978
rect 453154 238350 453774 255922
rect 453154 238294 453250 238350
rect 453306 238294 453374 238350
rect 453430 238294 453498 238350
rect 453554 238294 453622 238350
rect 453678 238294 453774 238350
rect 453154 238226 453774 238294
rect 453154 238170 453250 238226
rect 453306 238170 453374 238226
rect 453430 238170 453498 238226
rect 453554 238170 453622 238226
rect 453678 238170 453774 238226
rect 453154 238102 453774 238170
rect 453154 238046 453250 238102
rect 453306 238046 453374 238102
rect 453430 238046 453498 238102
rect 453554 238046 453622 238102
rect 453678 238046 453774 238102
rect 453154 237978 453774 238046
rect 453154 237922 453250 237978
rect 453306 237922 453374 237978
rect 453430 237922 453498 237978
rect 453554 237922 453622 237978
rect 453678 237922 453774 237978
rect 453154 220350 453774 237922
rect 453154 220294 453250 220350
rect 453306 220294 453374 220350
rect 453430 220294 453498 220350
rect 453554 220294 453622 220350
rect 453678 220294 453774 220350
rect 453154 220226 453774 220294
rect 453154 220170 453250 220226
rect 453306 220170 453374 220226
rect 453430 220170 453498 220226
rect 453554 220170 453622 220226
rect 453678 220170 453774 220226
rect 453154 220102 453774 220170
rect 453154 220046 453250 220102
rect 453306 220046 453374 220102
rect 453430 220046 453498 220102
rect 453554 220046 453622 220102
rect 453678 220046 453774 220102
rect 453154 219978 453774 220046
rect 453154 219922 453250 219978
rect 453306 219922 453374 219978
rect 453430 219922 453498 219978
rect 453554 219922 453622 219978
rect 453678 219922 453774 219978
rect 453154 217934 453774 219922
rect 456874 598172 457494 598268
rect 456874 598116 456970 598172
rect 457026 598116 457094 598172
rect 457150 598116 457218 598172
rect 457274 598116 457342 598172
rect 457398 598116 457494 598172
rect 456874 598048 457494 598116
rect 456874 597992 456970 598048
rect 457026 597992 457094 598048
rect 457150 597992 457218 598048
rect 457274 597992 457342 598048
rect 457398 597992 457494 598048
rect 456874 597924 457494 597992
rect 456874 597868 456970 597924
rect 457026 597868 457094 597924
rect 457150 597868 457218 597924
rect 457274 597868 457342 597924
rect 457398 597868 457494 597924
rect 456874 597800 457494 597868
rect 456874 597744 456970 597800
rect 457026 597744 457094 597800
rect 457150 597744 457218 597800
rect 457274 597744 457342 597800
rect 457398 597744 457494 597800
rect 456874 586350 457494 597744
rect 456874 586294 456970 586350
rect 457026 586294 457094 586350
rect 457150 586294 457218 586350
rect 457274 586294 457342 586350
rect 457398 586294 457494 586350
rect 456874 586226 457494 586294
rect 456874 586170 456970 586226
rect 457026 586170 457094 586226
rect 457150 586170 457218 586226
rect 457274 586170 457342 586226
rect 457398 586170 457494 586226
rect 456874 586102 457494 586170
rect 456874 586046 456970 586102
rect 457026 586046 457094 586102
rect 457150 586046 457218 586102
rect 457274 586046 457342 586102
rect 457398 586046 457494 586102
rect 456874 585978 457494 586046
rect 456874 585922 456970 585978
rect 457026 585922 457094 585978
rect 457150 585922 457218 585978
rect 457274 585922 457342 585978
rect 457398 585922 457494 585978
rect 456874 568350 457494 585922
rect 456874 568294 456970 568350
rect 457026 568294 457094 568350
rect 457150 568294 457218 568350
rect 457274 568294 457342 568350
rect 457398 568294 457494 568350
rect 456874 568226 457494 568294
rect 456874 568170 456970 568226
rect 457026 568170 457094 568226
rect 457150 568170 457218 568226
rect 457274 568170 457342 568226
rect 457398 568170 457494 568226
rect 456874 568102 457494 568170
rect 456874 568046 456970 568102
rect 457026 568046 457094 568102
rect 457150 568046 457218 568102
rect 457274 568046 457342 568102
rect 457398 568046 457494 568102
rect 456874 567978 457494 568046
rect 456874 567922 456970 567978
rect 457026 567922 457094 567978
rect 457150 567922 457218 567978
rect 457274 567922 457342 567978
rect 457398 567922 457494 567978
rect 456874 550350 457494 567922
rect 456874 550294 456970 550350
rect 457026 550294 457094 550350
rect 457150 550294 457218 550350
rect 457274 550294 457342 550350
rect 457398 550294 457494 550350
rect 456874 550226 457494 550294
rect 456874 550170 456970 550226
rect 457026 550170 457094 550226
rect 457150 550170 457218 550226
rect 457274 550170 457342 550226
rect 457398 550170 457494 550226
rect 456874 550102 457494 550170
rect 456874 550046 456970 550102
rect 457026 550046 457094 550102
rect 457150 550046 457218 550102
rect 457274 550046 457342 550102
rect 457398 550046 457494 550102
rect 456874 549978 457494 550046
rect 456874 549922 456970 549978
rect 457026 549922 457094 549978
rect 457150 549922 457218 549978
rect 457274 549922 457342 549978
rect 457398 549922 457494 549978
rect 456874 532350 457494 549922
rect 456874 532294 456970 532350
rect 457026 532294 457094 532350
rect 457150 532294 457218 532350
rect 457274 532294 457342 532350
rect 457398 532294 457494 532350
rect 456874 532226 457494 532294
rect 456874 532170 456970 532226
rect 457026 532170 457094 532226
rect 457150 532170 457218 532226
rect 457274 532170 457342 532226
rect 457398 532170 457494 532226
rect 456874 532102 457494 532170
rect 456874 532046 456970 532102
rect 457026 532046 457094 532102
rect 457150 532046 457218 532102
rect 457274 532046 457342 532102
rect 457398 532046 457494 532102
rect 456874 531978 457494 532046
rect 456874 531922 456970 531978
rect 457026 531922 457094 531978
rect 457150 531922 457218 531978
rect 457274 531922 457342 531978
rect 457398 531922 457494 531978
rect 456874 514350 457494 531922
rect 456874 514294 456970 514350
rect 457026 514294 457094 514350
rect 457150 514294 457218 514350
rect 457274 514294 457342 514350
rect 457398 514294 457494 514350
rect 456874 514226 457494 514294
rect 456874 514170 456970 514226
rect 457026 514170 457094 514226
rect 457150 514170 457218 514226
rect 457274 514170 457342 514226
rect 457398 514170 457494 514226
rect 456874 514102 457494 514170
rect 456874 514046 456970 514102
rect 457026 514046 457094 514102
rect 457150 514046 457218 514102
rect 457274 514046 457342 514102
rect 457398 514046 457494 514102
rect 456874 513978 457494 514046
rect 456874 513922 456970 513978
rect 457026 513922 457094 513978
rect 457150 513922 457218 513978
rect 457274 513922 457342 513978
rect 457398 513922 457494 513978
rect 456874 496350 457494 513922
rect 456874 496294 456970 496350
rect 457026 496294 457094 496350
rect 457150 496294 457218 496350
rect 457274 496294 457342 496350
rect 457398 496294 457494 496350
rect 456874 496226 457494 496294
rect 456874 496170 456970 496226
rect 457026 496170 457094 496226
rect 457150 496170 457218 496226
rect 457274 496170 457342 496226
rect 457398 496170 457494 496226
rect 456874 496102 457494 496170
rect 456874 496046 456970 496102
rect 457026 496046 457094 496102
rect 457150 496046 457218 496102
rect 457274 496046 457342 496102
rect 457398 496046 457494 496102
rect 456874 495978 457494 496046
rect 456874 495922 456970 495978
rect 457026 495922 457094 495978
rect 457150 495922 457218 495978
rect 457274 495922 457342 495978
rect 457398 495922 457494 495978
rect 456874 478350 457494 495922
rect 456874 478294 456970 478350
rect 457026 478294 457094 478350
rect 457150 478294 457218 478350
rect 457274 478294 457342 478350
rect 457398 478294 457494 478350
rect 456874 478226 457494 478294
rect 456874 478170 456970 478226
rect 457026 478170 457094 478226
rect 457150 478170 457218 478226
rect 457274 478170 457342 478226
rect 457398 478170 457494 478226
rect 456874 478102 457494 478170
rect 456874 478046 456970 478102
rect 457026 478046 457094 478102
rect 457150 478046 457218 478102
rect 457274 478046 457342 478102
rect 457398 478046 457494 478102
rect 456874 477978 457494 478046
rect 456874 477922 456970 477978
rect 457026 477922 457094 477978
rect 457150 477922 457218 477978
rect 457274 477922 457342 477978
rect 457398 477922 457494 477978
rect 456874 460350 457494 477922
rect 456874 460294 456970 460350
rect 457026 460294 457094 460350
rect 457150 460294 457218 460350
rect 457274 460294 457342 460350
rect 457398 460294 457494 460350
rect 456874 460226 457494 460294
rect 456874 460170 456970 460226
rect 457026 460170 457094 460226
rect 457150 460170 457218 460226
rect 457274 460170 457342 460226
rect 457398 460170 457494 460226
rect 456874 460102 457494 460170
rect 456874 460046 456970 460102
rect 457026 460046 457094 460102
rect 457150 460046 457218 460102
rect 457274 460046 457342 460102
rect 457398 460046 457494 460102
rect 456874 459978 457494 460046
rect 456874 459922 456970 459978
rect 457026 459922 457094 459978
rect 457150 459922 457218 459978
rect 457274 459922 457342 459978
rect 457398 459922 457494 459978
rect 456874 442350 457494 459922
rect 456874 442294 456970 442350
rect 457026 442294 457094 442350
rect 457150 442294 457218 442350
rect 457274 442294 457342 442350
rect 457398 442294 457494 442350
rect 456874 442226 457494 442294
rect 456874 442170 456970 442226
rect 457026 442170 457094 442226
rect 457150 442170 457218 442226
rect 457274 442170 457342 442226
rect 457398 442170 457494 442226
rect 456874 442102 457494 442170
rect 456874 442046 456970 442102
rect 457026 442046 457094 442102
rect 457150 442046 457218 442102
rect 457274 442046 457342 442102
rect 457398 442046 457494 442102
rect 456874 441978 457494 442046
rect 456874 441922 456970 441978
rect 457026 441922 457094 441978
rect 457150 441922 457218 441978
rect 457274 441922 457342 441978
rect 457398 441922 457494 441978
rect 456874 424350 457494 441922
rect 456874 424294 456970 424350
rect 457026 424294 457094 424350
rect 457150 424294 457218 424350
rect 457274 424294 457342 424350
rect 457398 424294 457494 424350
rect 456874 424226 457494 424294
rect 456874 424170 456970 424226
rect 457026 424170 457094 424226
rect 457150 424170 457218 424226
rect 457274 424170 457342 424226
rect 457398 424170 457494 424226
rect 456874 424102 457494 424170
rect 456874 424046 456970 424102
rect 457026 424046 457094 424102
rect 457150 424046 457218 424102
rect 457274 424046 457342 424102
rect 457398 424046 457494 424102
rect 456874 423978 457494 424046
rect 456874 423922 456970 423978
rect 457026 423922 457094 423978
rect 457150 423922 457218 423978
rect 457274 423922 457342 423978
rect 457398 423922 457494 423978
rect 456874 406350 457494 423922
rect 456874 406294 456970 406350
rect 457026 406294 457094 406350
rect 457150 406294 457218 406350
rect 457274 406294 457342 406350
rect 457398 406294 457494 406350
rect 456874 406226 457494 406294
rect 456874 406170 456970 406226
rect 457026 406170 457094 406226
rect 457150 406170 457218 406226
rect 457274 406170 457342 406226
rect 457398 406170 457494 406226
rect 456874 406102 457494 406170
rect 456874 406046 456970 406102
rect 457026 406046 457094 406102
rect 457150 406046 457218 406102
rect 457274 406046 457342 406102
rect 457398 406046 457494 406102
rect 456874 405978 457494 406046
rect 456874 405922 456970 405978
rect 457026 405922 457094 405978
rect 457150 405922 457218 405978
rect 457274 405922 457342 405978
rect 457398 405922 457494 405978
rect 456874 388350 457494 405922
rect 456874 388294 456970 388350
rect 457026 388294 457094 388350
rect 457150 388294 457218 388350
rect 457274 388294 457342 388350
rect 457398 388294 457494 388350
rect 456874 388226 457494 388294
rect 456874 388170 456970 388226
rect 457026 388170 457094 388226
rect 457150 388170 457218 388226
rect 457274 388170 457342 388226
rect 457398 388170 457494 388226
rect 456874 388102 457494 388170
rect 456874 388046 456970 388102
rect 457026 388046 457094 388102
rect 457150 388046 457218 388102
rect 457274 388046 457342 388102
rect 457398 388046 457494 388102
rect 456874 387978 457494 388046
rect 456874 387922 456970 387978
rect 457026 387922 457094 387978
rect 457150 387922 457218 387978
rect 457274 387922 457342 387978
rect 457398 387922 457494 387978
rect 456874 370350 457494 387922
rect 456874 370294 456970 370350
rect 457026 370294 457094 370350
rect 457150 370294 457218 370350
rect 457274 370294 457342 370350
rect 457398 370294 457494 370350
rect 456874 370226 457494 370294
rect 456874 370170 456970 370226
rect 457026 370170 457094 370226
rect 457150 370170 457218 370226
rect 457274 370170 457342 370226
rect 457398 370170 457494 370226
rect 456874 370102 457494 370170
rect 456874 370046 456970 370102
rect 457026 370046 457094 370102
rect 457150 370046 457218 370102
rect 457274 370046 457342 370102
rect 457398 370046 457494 370102
rect 456874 369978 457494 370046
rect 456874 369922 456970 369978
rect 457026 369922 457094 369978
rect 457150 369922 457218 369978
rect 457274 369922 457342 369978
rect 457398 369922 457494 369978
rect 456874 352350 457494 369922
rect 456874 352294 456970 352350
rect 457026 352294 457094 352350
rect 457150 352294 457218 352350
rect 457274 352294 457342 352350
rect 457398 352294 457494 352350
rect 456874 352226 457494 352294
rect 456874 352170 456970 352226
rect 457026 352170 457094 352226
rect 457150 352170 457218 352226
rect 457274 352170 457342 352226
rect 457398 352170 457494 352226
rect 456874 352102 457494 352170
rect 456874 352046 456970 352102
rect 457026 352046 457094 352102
rect 457150 352046 457218 352102
rect 457274 352046 457342 352102
rect 457398 352046 457494 352102
rect 456874 351978 457494 352046
rect 456874 351922 456970 351978
rect 457026 351922 457094 351978
rect 457150 351922 457218 351978
rect 457274 351922 457342 351978
rect 457398 351922 457494 351978
rect 456874 334350 457494 351922
rect 456874 334294 456970 334350
rect 457026 334294 457094 334350
rect 457150 334294 457218 334350
rect 457274 334294 457342 334350
rect 457398 334294 457494 334350
rect 456874 334226 457494 334294
rect 456874 334170 456970 334226
rect 457026 334170 457094 334226
rect 457150 334170 457218 334226
rect 457274 334170 457342 334226
rect 457398 334170 457494 334226
rect 456874 334102 457494 334170
rect 456874 334046 456970 334102
rect 457026 334046 457094 334102
rect 457150 334046 457218 334102
rect 457274 334046 457342 334102
rect 457398 334046 457494 334102
rect 456874 333978 457494 334046
rect 456874 333922 456970 333978
rect 457026 333922 457094 333978
rect 457150 333922 457218 333978
rect 457274 333922 457342 333978
rect 457398 333922 457494 333978
rect 456874 316350 457494 333922
rect 456874 316294 456970 316350
rect 457026 316294 457094 316350
rect 457150 316294 457218 316350
rect 457274 316294 457342 316350
rect 457398 316294 457494 316350
rect 456874 316226 457494 316294
rect 456874 316170 456970 316226
rect 457026 316170 457094 316226
rect 457150 316170 457218 316226
rect 457274 316170 457342 316226
rect 457398 316170 457494 316226
rect 456874 316102 457494 316170
rect 456874 316046 456970 316102
rect 457026 316046 457094 316102
rect 457150 316046 457218 316102
rect 457274 316046 457342 316102
rect 457398 316046 457494 316102
rect 456874 315978 457494 316046
rect 456874 315922 456970 315978
rect 457026 315922 457094 315978
rect 457150 315922 457218 315978
rect 457274 315922 457342 315978
rect 457398 315922 457494 315978
rect 456874 298350 457494 315922
rect 456874 298294 456970 298350
rect 457026 298294 457094 298350
rect 457150 298294 457218 298350
rect 457274 298294 457342 298350
rect 457398 298294 457494 298350
rect 456874 298226 457494 298294
rect 456874 298170 456970 298226
rect 457026 298170 457094 298226
rect 457150 298170 457218 298226
rect 457274 298170 457342 298226
rect 457398 298170 457494 298226
rect 456874 298102 457494 298170
rect 456874 298046 456970 298102
rect 457026 298046 457094 298102
rect 457150 298046 457218 298102
rect 457274 298046 457342 298102
rect 457398 298046 457494 298102
rect 456874 297978 457494 298046
rect 456874 297922 456970 297978
rect 457026 297922 457094 297978
rect 457150 297922 457218 297978
rect 457274 297922 457342 297978
rect 457398 297922 457494 297978
rect 456874 280350 457494 297922
rect 456874 280294 456970 280350
rect 457026 280294 457094 280350
rect 457150 280294 457218 280350
rect 457274 280294 457342 280350
rect 457398 280294 457494 280350
rect 456874 280226 457494 280294
rect 456874 280170 456970 280226
rect 457026 280170 457094 280226
rect 457150 280170 457218 280226
rect 457274 280170 457342 280226
rect 457398 280170 457494 280226
rect 456874 280102 457494 280170
rect 456874 280046 456970 280102
rect 457026 280046 457094 280102
rect 457150 280046 457218 280102
rect 457274 280046 457342 280102
rect 457398 280046 457494 280102
rect 456874 279978 457494 280046
rect 456874 279922 456970 279978
rect 457026 279922 457094 279978
rect 457150 279922 457218 279978
rect 457274 279922 457342 279978
rect 457398 279922 457494 279978
rect 456874 262350 457494 279922
rect 456874 262294 456970 262350
rect 457026 262294 457094 262350
rect 457150 262294 457218 262350
rect 457274 262294 457342 262350
rect 457398 262294 457494 262350
rect 456874 262226 457494 262294
rect 456874 262170 456970 262226
rect 457026 262170 457094 262226
rect 457150 262170 457218 262226
rect 457274 262170 457342 262226
rect 457398 262170 457494 262226
rect 456874 262102 457494 262170
rect 456874 262046 456970 262102
rect 457026 262046 457094 262102
rect 457150 262046 457218 262102
rect 457274 262046 457342 262102
rect 457398 262046 457494 262102
rect 456874 261978 457494 262046
rect 456874 261922 456970 261978
rect 457026 261922 457094 261978
rect 457150 261922 457218 261978
rect 457274 261922 457342 261978
rect 457398 261922 457494 261978
rect 456874 244350 457494 261922
rect 456874 244294 456970 244350
rect 457026 244294 457094 244350
rect 457150 244294 457218 244350
rect 457274 244294 457342 244350
rect 457398 244294 457494 244350
rect 456874 244226 457494 244294
rect 456874 244170 456970 244226
rect 457026 244170 457094 244226
rect 457150 244170 457218 244226
rect 457274 244170 457342 244226
rect 457398 244170 457494 244226
rect 456874 244102 457494 244170
rect 456874 244046 456970 244102
rect 457026 244046 457094 244102
rect 457150 244046 457218 244102
rect 457274 244046 457342 244102
rect 457398 244046 457494 244102
rect 456874 243978 457494 244046
rect 456874 243922 456970 243978
rect 457026 243922 457094 243978
rect 457150 243922 457218 243978
rect 457274 243922 457342 243978
rect 457398 243922 457494 243978
rect 456874 226350 457494 243922
rect 456874 226294 456970 226350
rect 457026 226294 457094 226350
rect 457150 226294 457218 226350
rect 457274 226294 457342 226350
rect 457398 226294 457494 226350
rect 456874 226226 457494 226294
rect 456874 226170 456970 226226
rect 457026 226170 457094 226226
rect 457150 226170 457218 226226
rect 457274 226170 457342 226226
rect 457398 226170 457494 226226
rect 456874 226102 457494 226170
rect 456874 226046 456970 226102
rect 457026 226046 457094 226102
rect 457150 226046 457218 226102
rect 457274 226046 457342 226102
rect 457398 226046 457494 226102
rect 456874 225978 457494 226046
rect 456874 225922 456970 225978
rect 457026 225922 457094 225978
rect 457150 225922 457218 225978
rect 457274 225922 457342 225978
rect 457398 225922 457494 225978
rect 456874 217934 457494 225922
rect 471154 597212 471774 598268
rect 471154 597156 471250 597212
rect 471306 597156 471374 597212
rect 471430 597156 471498 597212
rect 471554 597156 471622 597212
rect 471678 597156 471774 597212
rect 471154 597088 471774 597156
rect 471154 597032 471250 597088
rect 471306 597032 471374 597088
rect 471430 597032 471498 597088
rect 471554 597032 471622 597088
rect 471678 597032 471774 597088
rect 471154 596964 471774 597032
rect 471154 596908 471250 596964
rect 471306 596908 471374 596964
rect 471430 596908 471498 596964
rect 471554 596908 471622 596964
rect 471678 596908 471774 596964
rect 471154 596840 471774 596908
rect 471154 596784 471250 596840
rect 471306 596784 471374 596840
rect 471430 596784 471498 596840
rect 471554 596784 471622 596840
rect 471678 596784 471774 596840
rect 471154 580350 471774 596784
rect 489154 597212 489774 598268
rect 489154 597156 489250 597212
rect 489306 597156 489374 597212
rect 489430 597156 489498 597212
rect 489554 597156 489622 597212
rect 489678 597156 489774 597212
rect 489154 597088 489774 597156
rect 489154 597032 489250 597088
rect 489306 597032 489374 597088
rect 489430 597032 489498 597088
rect 489554 597032 489622 597088
rect 489678 597032 489774 597088
rect 489154 596964 489774 597032
rect 489154 596908 489250 596964
rect 489306 596908 489374 596964
rect 489430 596908 489498 596964
rect 489554 596908 489622 596964
rect 489678 596908 489774 596964
rect 489154 596840 489774 596908
rect 489154 596784 489250 596840
rect 489306 596784 489374 596840
rect 489430 596784 489498 596840
rect 489554 596784 489622 596840
rect 489678 596784 489774 596840
rect 474572 589764 474628 589774
rect 474572 589316 474628 589708
rect 474572 589250 474628 589260
rect 471154 580294 471250 580350
rect 471306 580294 471374 580350
rect 471430 580294 471498 580350
rect 471554 580294 471622 580350
rect 471678 580294 471774 580350
rect 471154 580226 471774 580294
rect 471154 580170 471250 580226
rect 471306 580170 471374 580226
rect 471430 580170 471498 580226
rect 471554 580170 471622 580226
rect 471678 580170 471774 580226
rect 471154 580102 471774 580170
rect 471154 580046 471250 580102
rect 471306 580046 471374 580102
rect 471430 580046 471498 580102
rect 471554 580046 471622 580102
rect 471678 580046 471774 580102
rect 471154 579978 471774 580046
rect 471154 579922 471250 579978
rect 471306 579922 471374 579978
rect 471430 579922 471498 579978
rect 471554 579922 471622 579978
rect 471678 579922 471774 579978
rect 471154 562350 471774 579922
rect 471154 562294 471250 562350
rect 471306 562294 471374 562350
rect 471430 562294 471498 562350
rect 471554 562294 471622 562350
rect 471678 562294 471774 562350
rect 471154 562226 471774 562294
rect 471154 562170 471250 562226
rect 471306 562170 471374 562226
rect 471430 562170 471498 562226
rect 471554 562170 471622 562226
rect 471678 562170 471774 562226
rect 471154 562102 471774 562170
rect 471154 562046 471250 562102
rect 471306 562046 471374 562102
rect 471430 562046 471498 562102
rect 471554 562046 471622 562102
rect 471678 562046 471774 562102
rect 471154 561978 471774 562046
rect 471154 561922 471250 561978
rect 471306 561922 471374 561978
rect 471430 561922 471498 561978
rect 471554 561922 471622 561978
rect 471678 561922 471774 561978
rect 471154 544350 471774 561922
rect 471154 544294 471250 544350
rect 471306 544294 471374 544350
rect 471430 544294 471498 544350
rect 471554 544294 471622 544350
rect 471678 544294 471774 544350
rect 471154 544226 471774 544294
rect 471154 544170 471250 544226
rect 471306 544170 471374 544226
rect 471430 544170 471498 544226
rect 471554 544170 471622 544226
rect 471678 544170 471774 544226
rect 471154 544102 471774 544170
rect 471154 544046 471250 544102
rect 471306 544046 471374 544102
rect 471430 544046 471498 544102
rect 471554 544046 471622 544102
rect 471678 544046 471774 544102
rect 471154 543978 471774 544046
rect 471154 543922 471250 543978
rect 471306 543922 471374 543978
rect 471430 543922 471498 543978
rect 471554 543922 471622 543978
rect 471678 543922 471774 543978
rect 471154 526350 471774 543922
rect 471154 526294 471250 526350
rect 471306 526294 471374 526350
rect 471430 526294 471498 526350
rect 471554 526294 471622 526350
rect 471678 526294 471774 526350
rect 471154 526226 471774 526294
rect 471154 526170 471250 526226
rect 471306 526170 471374 526226
rect 471430 526170 471498 526226
rect 471554 526170 471622 526226
rect 471678 526170 471774 526226
rect 471154 526102 471774 526170
rect 471154 526046 471250 526102
rect 471306 526046 471374 526102
rect 471430 526046 471498 526102
rect 471554 526046 471622 526102
rect 471678 526046 471774 526102
rect 471154 525978 471774 526046
rect 471154 525922 471250 525978
rect 471306 525922 471374 525978
rect 471430 525922 471498 525978
rect 471554 525922 471622 525978
rect 471678 525922 471774 525978
rect 471154 508350 471774 525922
rect 471154 508294 471250 508350
rect 471306 508294 471374 508350
rect 471430 508294 471498 508350
rect 471554 508294 471622 508350
rect 471678 508294 471774 508350
rect 471154 508226 471774 508294
rect 471154 508170 471250 508226
rect 471306 508170 471374 508226
rect 471430 508170 471498 508226
rect 471554 508170 471622 508226
rect 471678 508170 471774 508226
rect 471154 508102 471774 508170
rect 471154 508046 471250 508102
rect 471306 508046 471374 508102
rect 471430 508046 471498 508102
rect 471554 508046 471622 508102
rect 471678 508046 471774 508102
rect 471154 507978 471774 508046
rect 471154 507922 471250 507978
rect 471306 507922 471374 507978
rect 471430 507922 471498 507978
rect 471554 507922 471622 507978
rect 471678 507922 471774 507978
rect 471154 490350 471774 507922
rect 471154 490294 471250 490350
rect 471306 490294 471374 490350
rect 471430 490294 471498 490350
rect 471554 490294 471622 490350
rect 471678 490294 471774 490350
rect 471154 490226 471774 490294
rect 471154 490170 471250 490226
rect 471306 490170 471374 490226
rect 471430 490170 471498 490226
rect 471554 490170 471622 490226
rect 471678 490170 471774 490226
rect 471154 490102 471774 490170
rect 471154 490046 471250 490102
rect 471306 490046 471374 490102
rect 471430 490046 471498 490102
rect 471554 490046 471622 490102
rect 471678 490046 471774 490102
rect 471154 489978 471774 490046
rect 471154 489922 471250 489978
rect 471306 489922 471374 489978
rect 471430 489922 471498 489978
rect 471554 489922 471622 489978
rect 471678 489922 471774 489978
rect 471154 472350 471774 489922
rect 471154 472294 471250 472350
rect 471306 472294 471374 472350
rect 471430 472294 471498 472350
rect 471554 472294 471622 472350
rect 471678 472294 471774 472350
rect 471154 472226 471774 472294
rect 471154 472170 471250 472226
rect 471306 472170 471374 472226
rect 471430 472170 471498 472226
rect 471554 472170 471622 472226
rect 471678 472170 471774 472226
rect 471154 472102 471774 472170
rect 471154 472046 471250 472102
rect 471306 472046 471374 472102
rect 471430 472046 471498 472102
rect 471554 472046 471622 472102
rect 471678 472046 471774 472102
rect 471154 471978 471774 472046
rect 471154 471922 471250 471978
rect 471306 471922 471374 471978
rect 471430 471922 471498 471978
rect 471554 471922 471622 471978
rect 471678 471922 471774 471978
rect 471154 454350 471774 471922
rect 471154 454294 471250 454350
rect 471306 454294 471374 454350
rect 471430 454294 471498 454350
rect 471554 454294 471622 454350
rect 471678 454294 471774 454350
rect 471154 454226 471774 454294
rect 471154 454170 471250 454226
rect 471306 454170 471374 454226
rect 471430 454170 471498 454226
rect 471554 454170 471622 454226
rect 471678 454170 471774 454226
rect 471154 454102 471774 454170
rect 471154 454046 471250 454102
rect 471306 454046 471374 454102
rect 471430 454046 471498 454102
rect 471554 454046 471622 454102
rect 471678 454046 471774 454102
rect 471154 453978 471774 454046
rect 471154 453922 471250 453978
rect 471306 453922 471374 453978
rect 471430 453922 471498 453978
rect 471554 453922 471622 453978
rect 471678 453922 471774 453978
rect 471154 436350 471774 453922
rect 471154 436294 471250 436350
rect 471306 436294 471374 436350
rect 471430 436294 471498 436350
rect 471554 436294 471622 436350
rect 471678 436294 471774 436350
rect 471154 436226 471774 436294
rect 471154 436170 471250 436226
rect 471306 436170 471374 436226
rect 471430 436170 471498 436226
rect 471554 436170 471622 436226
rect 471678 436170 471774 436226
rect 471154 436102 471774 436170
rect 471154 436046 471250 436102
rect 471306 436046 471374 436102
rect 471430 436046 471498 436102
rect 471554 436046 471622 436102
rect 471678 436046 471774 436102
rect 471154 435978 471774 436046
rect 471154 435922 471250 435978
rect 471306 435922 471374 435978
rect 471430 435922 471498 435978
rect 471554 435922 471622 435978
rect 471678 435922 471774 435978
rect 471154 418350 471774 435922
rect 471154 418294 471250 418350
rect 471306 418294 471374 418350
rect 471430 418294 471498 418350
rect 471554 418294 471622 418350
rect 471678 418294 471774 418350
rect 471154 418226 471774 418294
rect 471154 418170 471250 418226
rect 471306 418170 471374 418226
rect 471430 418170 471498 418226
rect 471554 418170 471622 418226
rect 471678 418170 471774 418226
rect 471154 418102 471774 418170
rect 471154 418046 471250 418102
rect 471306 418046 471374 418102
rect 471430 418046 471498 418102
rect 471554 418046 471622 418102
rect 471678 418046 471774 418102
rect 471154 417978 471774 418046
rect 471154 417922 471250 417978
rect 471306 417922 471374 417978
rect 471430 417922 471498 417978
rect 471554 417922 471622 417978
rect 471678 417922 471774 417978
rect 471154 400350 471774 417922
rect 471154 400294 471250 400350
rect 471306 400294 471374 400350
rect 471430 400294 471498 400350
rect 471554 400294 471622 400350
rect 471678 400294 471774 400350
rect 471154 400226 471774 400294
rect 471154 400170 471250 400226
rect 471306 400170 471374 400226
rect 471430 400170 471498 400226
rect 471554 400170 471622 400226
rect 471678 400170 471774 400226
rect 471154 400102 471774 400170
rect 471154 400046 471250 400102
rect 471306 400046 471374 400102
rect 471430 400046 471498 400102
rect 471554 400046 471622 400102
rect 471678 400046 471774 400102
rect 471154 399978 471774 400046
rect 471154 399922 471250 399978
rect 471306 399922 471374 399978
rect 471430 399922 471498 399978
rect 471554 399922 471622 399978
rect 471678 399922 471774 399978
rect 471154 382350 471774 399922
rect 471154 382294 471250 382350
rect 471306 382294 471374 382350
rect 471430 382294 471498 382350
rect 471554 382294 471622 382350
rect 471678 382294 471774 382350
rect 471154 382226 471774 382294
rect 471154 382170 471250 382226
rect 471306 382170 471374 382226
rect 471430 382170 471498 382226
rect 471554 382170 471622 382226
rect 471678 382170 471774 382226
rect 471154 382102 471774 382170
rect 471154 382046 471250 382102
rect 471306 382046 471374 382102
rect 471430 382046 471498 382102
rect 471554 382046 471622 382102
rect 471678 382046 471774 382102
rect 471154 381978 471774 382046
rect 471154 381922 471250 381978
rect 471306 381922 471374 381978
rect 471430 381922 471498 381978
rect 471554 381922 471622 381978
rect 471678 381922 471774 381978
rect 471154 364350 471774 381922
rect 471154 364294 471250 364350
rect 471306 364294 471374 364350
rect 471430 364294 471498 364350
rect 471554 364294 471622 364350
rect 471678 364294 471774 364350
rect 471154 364226 471774 364294
rect 471154 364170 471250 364226
rect 471306 364170 471374 364226
rect 471430 364170 471498 364226
rect 471554 364170 471622 364226
rect 471678 364170 471774 364226
rect 471154 364102 471774 364170
rect 471154 364046 471250 364102
rect 471306 364046 471374 364102
rect 471430 364046 471498 364102
rect 471554 364046 471622 364102
rect 471678 364046 471774 364102
rect 471154 363978 471774 364046
rect 471154 363922 471250 363978
rect 471306 363922 471374 363978
rect 471430 363922 471498 363978
rect 471554 363922 471622 363978
rect 471678 363922 471774 363978
rect 471154 346350 471774 363922
rect 471154 346294 471250 346350
rect 471306 346294 471374 346350
rect 471430 346294 471498 346350
rect 471554 346294 471622 346350
rect 471678 346294 471774 346350
rect 471154 346226 471774 346294
rect 471154 346170 471250 346226
rect 471306 346170 471374 346226
rect 471430 346170 471498 346226
rect 471554 346170 471622 346226
rect 471678 346170 471774 346226
rect 471154 346102 471774 346170
rect 471154 346046 471250 346102
rect 471306 346046 471374 346102
rect 471430 346046 471498 346102
rect 471554 346046 471622 346102
rect 471678 346046 471774 346102
rect 471154 345978 471774 346046
rect 471154 345922 471250 345978
rect 471306 345922 471374 345978
rect 471430 345922 471498 345978
rect 471554 345922 471622 345978
rect 471678 345922 471774 345978
rect 471154 328350 471774 345922
rect 471154 328294 471250 328350
rect 471306 328294 471374 328350
rect 471430 328294 471498 328350
rect 471554 328294 471622 328350
rect 471678 328294 471774 328350
rect 471154 328226 471774 328294
rect 471154 328170 471250 328226
rect 471306 328170 471374 328226
rect 471430 328170 471498 328226
rect 471554 328170 471622 328226
rect 471678 328170 471774 328226
rect 471154 328102 471774 328170
rect 471154 328046 471250 328102
rect 471306 328046 471374 328102
rect 471430 328046 471498 328102
rect 471554 328046 471622 328102
rect 471678 328046 471774 328102
rect 471154 327978 471774 328046
rect 471154 327922 471250 327978
rect 471306 327922 471374 327978
rect 471430 327922 471498 327978
rect 471554 327922 471622 327978
rect 471678 327922 471774 327978
rect 471154 310350 471774 327922
rect 471154 310294 471250 310350
rect 471306 310294 471374 310350
rect 471430 310294 471498 310350
rect 471554 310294 471622 310350
rect 471678 310294 471774 310350
rect 471154 310226 471774 310294
rect 471154 310170 471250 310226
rect 471306 310170 471374 310226
rect 471430 310170 471498 310226
rect 471554 310170 471622 310226
rect 471678 310170 471774 310226
rect 471154 310102 471774 310170
rect 471154 310046 471250 310102
rect 471306 310046 471374 310102
rect 471430 310046 471498 310102
rect 471554 310046 471622 310102
rect 471678 310046 471774 310102
rect 471154 309978 471774 310046
rect 471154 309922 471250 309978
rect 471306 309922 471374 309978
rect 471430 309922 471498 309978
rect 471554 309922 471622 309978
rect 471678 309922 471774 309978
rect 471154 292350 471774 309922
rect 471154 292294 471250 292350
rect 471306 292294 471374 292350
rect 471430 292294 471498 292350
rect 471554 292294 471622 292350
rect 471678 292294 471774 292350
rect 471154 292226 471774 292294
rect 471154 292170 471250 292226
rect 471306 292170 471374 292226
rect 471430 292170 471498 292226
rect 471554 292170 471622 292226
rect 471678 292170 471774 292226
rect 471154 292102 471774 292170
rect 471154 292046 471250 292102
rect 471306 292046 471374 292102
rect 471430 292046 471498 292102
rect 471554 292046 471622 292102
rect 471678 292046 471774 292102
rect 471154 291978 471774 292046
rect 471154 291922 471250 291978
rect 471306 291922 471374 291978
rect 471430 291922 471498 291978
rect 471554 291922 471622 291978
rect 471678 291922 471774 291978
rect 471154 274350 471774 291922
rect 471154 274294 471250 274350
rect 471306 274294 471374 274350
rect 471430 274294 471498 274350
rect 471554 274294 471622 274350
rect 471678 274294 471774 274350
rect 471154 274226 471774 274294
rect 471154 274170 471250 274226
rect 471306 274170 471374 274226
rect 471430 274170 471498 274226
rect 471554 274170 471622 274226
rect 471678 274170 471774 274226
rect 471154 274102 471774 274170
rect 471154 274046 471250 274102
rect 471306 274046 471374 274102
rect 471430 274046 471498 274102
rect 471554 274046 471622 274102
rect 471678 274046 471774 274102
rect 471154 273978 471774 274046
rect 471154 273922 471250 273978
rect 471306 273922 471374 273978
rect 471430 273922 471498 273978
rect 471554 273922 471622 273978
rect 471678 273922 471774 273978
rect 471154 256350 471774 273922
rect 471154 256294 471250 256350
rect 471306 256294 471374 256350
rect 471430 256294 471498 256350
rect 471554 256294 471622 256350
rect 471678 256294 471774 256350
rect 471154 256226 471774 256294
rect 471154 256170 471250 256226
rect 471306 256170 471374 256226
rect 471430 256170 471498 256226
rect 471554 256170 471622 256226
rect 471678 256170 471774 256226
rect 471154 256102 471774 256170
rect 471154 256046 471250 256102
rect 471306 256046 471374 256102
rect 471430 256046 471498 256102
rect 471554 256046 471622 256102
rect 471678 256046 471774 256102
rect 471154 255978 471774 256046
rect 471154 255922 471250 255978
rect 471306 255922 471374 255978
rect 471430 255922 471498 255978
rect 471554 255922 471622 255978
rect 471678 255922 471774 255978
rect 471154 238350 471774 255922
rect 471154 238294 471250 238350
rect 471306 238294 471374 238350
rect 471430 238294 471498 238350
rect 471554 238294 471622 238350
rect 471678 238294 471774 238350
rect 471154 238226 471774 238294
rect 471154 238170 471250 238226
rect 471306 238170 471374 238226
rect 471430 238170 471498 238226
rect 471554 238170 471622 238226
rect 471678 238170 471774 238226
rect 471154 238102 471774 238170
rect 471154 238046 471250 238102
rect 471306 238046 471374 238102
rect 471430 238046 471498 238102
rect 471554 238046 471622 238102
rect 471678 238046 471774 238102
rect 471154 237978 471774 238046
rect 471154 237922 471250 237978
rect 471306 237922 471374 237978
rect 471430 237922 471498 237978
rect 471554 237922 471622 237978
rect 471678 237922 471774 237978
rect 471154 220350 471774 237922
rect 471154 220294 471250 220350
rect 471306 220294 471374 220350
rect 471430 220294 471498 220350
rect 471554 220294 471622 220350
rect 471678 220294 471774 220350
rect 471154 220226 471774 220294
rect 471154 220170 471250 220226
rect 471306 220170 471374 220226
rect 471430 220170 471498 220226
rect 471554 220170 471622 220226
rect 471678 220170 471774 220226
rect 471154 220102 471774 220170
rect 471154 220046 471250 220102
rect 471306 220046 471374 220102
rect 471430 220046 471498 220102
rect 471554 220046 471622 220102
rect 471678 220046 471774 220102
rect 471154 219978 471774 220046
rect 471154 219922 471250 219978
rect 471306 219922 471374 219978
rect 471430 219922 471498 219978
rect 471554 219922 471622 219978
rect 471678 219922 471774 219978
rect 471154 217934 471774 219922
rect 489154 580350 489774 596784
rect 489154 580294 489250 580350
rect 489306 580294 489374 580350
rect 489430 580294 489498 580350
rect 489554 580294 489622 580350
rect 489678 580294 489774 580350
rect 489154 580226 489774 580294
rect 489154 580170 489250 580226
rect 489306 580170 489374 580226
rect 489430 580170 489498 580226
rect 489554 580170 489622 580226
rect 489678 580170 489774 580226
rect 489154 580102 489774 580170
rect 489154 580046 489250 580102
rect 489306 580046 489374 580102
rect 489430 580046 489498 580102
rect 489554 580046 489622 580102
rect 489678 580046 489774 580102
rect 489154 579978 489774 580046
rect 489154 579922 489250 579978
rect 489306 579922 489374 579978
rect 489430 579922 489498 579978
rect 489554 579922 489622 579978
rect 489678 579922 489774 579978
rect 489154 562350 489774 579922
rect 489154 562294 489250 562350
rect 489306 562294 489374 562350
rect 489430 562294 489498 562350
rect 489554 562294 489622 562350
rect 489678 562294 489774 562350
rect 489154 562226 489774 562294
rect 489154 562170 489250 562226
rect 489306 562170 489374 562226
rect 489430 562170 489498 562226
rect 489554 562170 489622 562226
rect 489678 562170 489774 562226
rect 489154 562102 489774 562170
rect 489154 562046 489250 562102
rect 489306 562046 489374 562102
rect 489430 562046 489498 562102
rect 489554 562046 489622 562102
rect 489678 562046 489774 562102
rect 489154 561978 489774 562046
rect 489154 561922 489250 561978
rect 489306 561922 489374 561978
rect 489430 561922 489498 561978
rect 489554 561922 489622 561978
rect 489678 561922 489774 561978
rect 489154 544350 489774 561922
rect 489154 544294 489250 544350
rect 489306 544294 489374 544350
rect 489430 544294 489498 544350
rect 489554 544294 489622 544350
rect 489678 544294 489774 544350
rect 489154 544226 489774 544294
rect 489154 544170 489250 544226
rect 489306 544170 489374 544226
rect 489430 544170 489498 544226
rect 489554 544170 489622 544226
rect 489678 544170 489774 544226
rect 489154 544102 489774 544170
rect 489154 544046 489250 544102
rect 489306 544046 489374 544102
rect 489430 544046 489498 544102
rect 489554 544046 489622 544102
rect 489678 544046 489774 544102
rect 489154 543978 489774 544046
rect 489154 543922 489250 543978
rect 489306 543922 489374 543978
rect 489430 543922 489498 543978
rect 489554 543922 489622 543978
rect 489678 543922 489774 543978
rect 489154 526350 489774 543922
rect 489154 526294 489250 526350
rect 489306 526294 489374 526350
rect 489430 526294 489498 526350
rect 489554 526294 489622 526350
rect 489678 526294 489774 526350
rect 489154 526226 489774 526294
rect 489154 526170 489250 526226
rect 489306 526170 489374 526226
rect 489430 526170 489498 526226
rect 489554 526170 489622 526226
rect 489678 526170 489774 526226
rect 489154 526102 489774 526170
rect 489154 526046 489250 526102
rect 489306 526046 489374 526102
rect 489430 526046 489498 526102
rect 489554 526046 489622 526102
rect 489678 526046 489774 526102
rect 489154 525978 489774 526046
rect 489154 525922 489250 525978
rect 489306 525922 489374 525978
rect 489430 525922 489498 525978
rect 489554 525922 489622 525978
rect 489678 525922 489774 525978
rect 489154 508350 489774 525922
rect 489154 508294 489250 508350
rect 489306 508294 489374 508350
rect 489430 508294 489498 508350
rect 489554 508294 489622 508350
rect 489678 508294 489774 508350
rect 489154 508226 489774 508294
rect 489154 508170 489250 508226
rect 489306 508170 489374 508226
rect 489430 508170 489498 508226
rect 489554 508170 489622 508226
rect 489678 508170 489774 508226
rect 489154 508102 489774 508170
rect 489154 508046 489250 508102
rect 489306 508046 489374 508102
rect 489430 508046 489498 508102
rect 489554 508046 489622 508102
rect 489678 508046 489774 508102
rect 489154 507978 489774 508046
rect 489154 507922 489250 507978
rect 489306 507922 489374 507978
rect 489430 507922 489498 507978
rect 489554 507922 489622 507978
rect 489678 507922 489774 507978
rect 489154 490350 489774 507922
rect 489154 490294 489250 490350
rect 489306 490294 489374 490350
rect 489430 490294 489498 490350
rect 489554 490294 489622 490350
rect 489678 490294 489774 490350
rect 489154 490226 489774 490294
rect 489154 490170 489250 490226
rect 489306 490170 489374 490226
rect 489430 490170 489498 490226
rect 489554 490170 489622 490226
rect 489678 490170 489774 490226
rect 489154 490102 489774 490170
rect 489154 490046 489250 490102
rect 489306 490046 489374 490102
rect 489430 490046 489498 490102
rect 489554 490046 489622 490102
rect 489678 490046 489774 490102
rect 489154 489978 489774 490046
rect 489154 489922 489250 489978
rect 489306 489922 489374 489978
rect 489430 489922 489498 489978
rect 489554 489922 489622 489978
rect 489678 489922 489774 489978
rect 489154 472350 489774 489922
rect 489154 472294 489250 472350
rect 489306 472294 489374 472350
rect 489430 472294 489498 472350
rect 489554 472294 489622 472350
rect 489678 472294 489774 472350
rect 489154 472226 489774 472294
rect 489154 472170 489250 472226
rect 489306 472170 489374 472226
rect 489430 472170 489498 472226
rect 489554 472170 489622 472226
rect 489678 472170 489774 472226
rect 489154 472102 489774 472170
rect 489154 472046 489250 472102
rect 489306 472046 489374 472102
rect 489430 472046 489498 472102
rect 489554 472046 489622 472102
rect 489678 472046 489774 472102
rect 489154 471978 489774 472046
rect 489154 471922 489250 471978
rect 489306 471922 489374 471978
rect 489430 471922 489498 471978
rect 489554 471922 489622 471978
rect 489678 471922 489774 471978
rect 489154 454350 489774 471922
rect 489154 454294 489250 454350
rect 489306 454294 489374 454350
rect 489430 454294 489498 454350
rect 489554 454294 489622 454350
rect 489678 454294 489774 454350
rect 489154 454226 489774 454294
rect 489154 454170 489250 454226
rect 489306 454170 489374 454226
rect 489430 454170 489498 454226
rect 489554 454170 489622 454226
rect 489678 454170 489774 454226
rect 489154 454102 489774 454170
rect 489154 454046 489250 454102
rect 489306 454046 489374 454102
rect 489430 454046 489498 454102
rect 489554 454046 489622 454102
rect 489678 454046 489774 454102
rect 489154 453978 489774 454046
rect 489154 453922 489250 453978
rect 489306 453922 489374 453978
rect 489430 453922 489498 453978
rect 489554 453922 489622 453978
rect 489678 453922 489774 453978
rect 489154 436350 489774 453922
rect 489154 436294 489250 436350
rect 489306 436294 489374 436350
rect 489430 436294 489498 436350
rect 489554 436294 489622 436350
rect 489678 436294 489774 436350
rect 489154 436226 489774 436294
rect 489154 436170 489250 436226
rect 489306 436170 489374 436226
rect 489430 436170 489498 436226
rect 489554 436170 489622 436226
rect 489678 436170 489774 436226
rect 489154 436102 489774 436170
rect 489154 436046 489250 436102
rect 489306 436046 489374 436102
rect 489430 436046 489498 436102
rect 489554 436046 489622 436102
rect 489678 436046 489774 436102
rect 489154 435978 489774 436046
rect 489154 435922 489250 435978
rect 489306 435922 489374 435978
rect 489430 435922 489498 435978
rect 489554 435922 489622 435978
rect 489678 435922 489774 435978
rect 489154 418350 489774 435922
rect 489154 418294 489250 418350
rect 489306 418294 489374 418350
rect 489430 418294 489498 418350
rect 489554 418294 489622 418350
rect 489678 418294 489774 418350
rect 489154 418226 489774 418294
rect 489154 418170 489250 418226
rect 489306 418170 489374 418226
rect 489430 418170 489498 418226
rect 489554 418170 489622 418226
rect 489678 418170 489774 418226
rect 489154 418102 489774 418170
rect 489154 418046 489250 418102
rect 489306 418046 489374 418102
rect 489430 418046 489498 418102
rect 489554 418046 489622 418102
rect 489678 418046 489774 418102
rect 489154 417978 489774 418046
rect 489154 417922 489250 417978
rect 489306 417922 489374 417978
rect 489430 417922 489498 417978
rect 489554 417922 489622 417978
rect 489678 417922 489774 417978
rect 489154 400350 489774 417922
rect 489154 400294 489250 400350
rect 489306 400294 489374 400350
rect 489430 400294 489498 400350
rect 489554 400294 489622 400350
rect 489678 400294 489774 400350
rect 489154 400226 489774 400294
rect 489154 400170 489250 400226
rect 489306 400170 489374 400226
rect 489430 400170 489498 400226
rect 489554 400170 489622 400226
rect 489678 400170 489774 400226
rect 489154 400102 489774 400170
rect 489154 400046 489250 400102
rect 489306 400046 489374 400102
rect 489430 400046 489498 400102
rect 489554 400046 489622 400102
rect 489678 400046 489774 400102
rect 489154 399978 489774 400046
rect 489154 399922 489250 399978
rect 489306 399922 489374 399978
rect 489430 399922 489498 399978
rect 489554 399922 489622 399978
rect 489678 399922 489774 399978
rect 489154 382350 489774 399922
rect 489154 382294 489250 382350
rect 489306 382294 489374 382350
rect 489430 382294 489498 382350
rect 489554 382294 489622 382350
rect 489678 382294 489774 382350
rect 489154 382226 489774 382294
rect 489154 382170 489250 382226
rect 489306 382170 489374 382226
rect 489430 382170 489498 382226
rect 489554 382170 489622 382226
rect 489678 382170 489774 382226
rect 489154 382102 489774 382170
rect 489154 382046 489250 382102
rect 489306 382046 489374 382102
rect 489430 382046 489498 382102
rect 489554 382046 489622 382102
rect 489678 382046 489774 382102
rect 489154 381978 489774 382046
rect 489154 381922 489250 381978
rect 489306 381922 489374 381978
rect 489430 381922 489498 381978
rect 489554 381922 489622 381978
rect 489678 381922 489774 381978
rect 489154 364350 489774 381922
rect 489154 364294 489250 364350
rect 489306 364294 489374 364350
rect 489430 364294 489498 364350
rect 489554 364294 489622 364350
rect 489678 364294 489774 364350
rect 489154 364226 489774 364294
rect 489154 364170 489250 364226
rect 489306 364170 489374 364226
rect 489430 364170 489498 364226
rect 489554 364170 489622 364226
rect 489678 364170 489774 364226
rect 489154 364102 489774 364170
rect 489154 364046 489250 364102
rect 489306 364046 489374 364102
rect 489430 364046 489498 364102
rect 489554 364046 489622 364102
rect 489678 364046 489774 364102
rect 489154 363978 489774 364046
rect 489154 363922 489250 363978
rect 489306 363922 489374 363978
rect 489430 363922 489498 363978
rect 489554 363922 489622 363978
rect 489678 363922 489774 363978
rect 489154 346350 489774 363922
rect 489154 346294 489250 346350
rect 489306 346294 489374 346350
rect 489430 346294 489498 346350
rect 489554 346294 489622 346350
rect 489678 346294 489774 346350
rect 489154 346226 489774 346294
rect 489154 346170 489250 346226
rect 489306 346170 489374 346226
rect 489430 346170 489498 346226
rect 489554 346170 489622 346226
rect 489678 346170 489774 346226
rect 489154 346102 489774 346170
rect 489154 346046 489250 346102
rect 489306 346046 489374 346102
rect 489430 346046 489498 346102
rect 489554 346046 489622 346102
rect 489678 346046 489774 346102
rect 489154 345978 489774 346046
rect 489154 345922 489250 345978
rect 489306 345922 489374 345978
rect 489430 345922 489498 345978
rect 489554 345922 489622 345978
rect 489678 345922 489774 345978
rect 489154 328350 489774 345922
rect 489154 328294 489250 328350
rect 489306 328294 489374 328350
rect 489430 328294 489498 328350
rect 489554 328294 489622 328350
rect 489678 328294 489774 328350
rect 489154 328226 489774 328294
rect 489154 328170 489250 328226
rect 489306 328170 489374 328226
rect 489430 328170 489498 328226
rect 489554 328170 489622 328226
rect 489678 328170 489774 328226
rect 489154 328102 489774 328170
rect 489154 328046 489250 328102
rect 489306 328046 489374 328102
rect 489430 328046 489498 328102
rect 489554 328046 489622 328102
rect 489678 328046 489774 328102
rect 489154 327978 489774 328046
rect 489154 327922 489250 327978
rect 489306 327922 489374 327978
rect 489430 327922 489498 327978
rect 489554 327922 489622 327978
rect 489678 327922 489774 327978
rect 489154 310350 489774 327922
rect 489154 310294 489250 310350
rect 489306 310294 489374 310350
rect 489430 310294 489498 310350
rect 489554 310294 489622 310350
rect 489678 310294 489774 310350
rect 489154 310226 489774 310294
rect 489154 310170 489250 310226
rect 489306 310170 489374 310226
rect 489430 310170 489498 310226
rect 489554 310170 489622 310226
rect 489678 310170 489774 310226
rect 489154 310102 489774 310170
rect 489154 310046 489250 310102
rect 489306 310046 489374 310102
rect 489430 310046 489498 310102
rect 489554 310046 489622 310102
rect 489678 310046 489774 310102
rect 489154 309978 489774 310046
rect 489154 309922 489250 309978
rect 489306 309922 489374 309978
rect 489430 309922 489498 309978
rect 489554 309922 489622 309978
rect 489678 309922 489774 309978
rect 489154 292350 489774 309922
rect 489154 292294 489250 292350
rect 489306 292294 489374 292350
rect 489430 292294 489498 292350
rect 489554 292294 489622 292350
rect 489678 292294 489774 292350
rect 489154 292226 489774 292294
rect 489154 292170 489250 292226
rect 489306 292170 489374 292226
rect 489430 292170 489498 292226
rect 489554 292170 489622 292226
rect 489678 292170 489774 292226
rect 489154 292102 489774 292170
rect 489154 292046 489250 292102
rect 489306 292046 489374 292102
rect 489430 292046 489498 292102
rect 489554 292046 489622 292102
rect 489678 292046 489774 292102
rect 489154 291978 489774 292046
rect 489154 291922 489250 291978
rect 489306 291922 489374 291978
rect 489430 291922 489498 291978
rect 489554 291922 489622 291978
rect 489678 291922 489774 291978
rect 489154 274350 489774 291922
rect 489154 274294 489250 274350
rect 489306 274294 489374 274350
rect 489430 274294 489498 274350
rect 489554 274294 489622 274350
rect 489678 274294 489774 274350
rect 489154 274226 489774 274294
rect 489154 274170 489250 274226
rect 489306 274170 489374 274226
rect 489430 274170 489498 274226
rect 489554 274170 489622 274226
rect 489678 274170 489774 274226
rect 489154 274102 489774 274170
rect 489154 274046 489250 274102
rect 489306 274046 489374 274102
rect 489430 274046 489498 274102
rect 489554 274046 489622 274102
rect 489678 274046 489774 274102
rect 489154 273978 489774 274046
rect 489154 273922 489250 273978
rect 489306 273922 489374 273978
rect 489430 273922 489498 273978
rect 489554 273922 489622 273978
rect 489678 273922 489774 273978
rect 489154 256350 489774 273922
rect 489154 256294 489250 256350
rect 489306 256294 489374 256350
rect 489430 256294 489498 256350
rect 489554 256294 489622 256350
rect 489678 256294 489774 256350
rect 489154 256226 489774 256294
rect 489154 256170 489250 256226
rect 489306 256170 489374 256226
rect 489430 256170 489498 256226
rect 489554 256170 489622 256226
rect 489678 256170 489774 256226
rect 489154 256102 489774 256170
rect 489154 256046 489250 256102
rect 489306 256046 489374 256102
rect 489430 256046 489498 256102
rect 489554 256046 489622 256102
rect 489678 256046 489774 256102
rect 489154 255978 489774 256046
rect 489154 255922 489250 255978
rect 489306 255922 489374 255978
rect 489430 255922 489498 255978
rect 489554 255922 489622 255978
rect 489678 255922 489774 255978
rect 489154 238350 489774 255922
rect 489154 238294 489250 238350
rect 489306 238294 489374 238350
rect 489430 238294 489498 238350
rect 489554 238294 489622 238350
rect 489678 238294 489774 238350
rect 489154 238226 489774 238294
rect 489154 238170 489250 238226
rect 489306 238170 489374 238226
rect 489430 238170 489498 238226
rect 489554 238170 489622 238226
rect 489678 238170 489774 238226
rect 489154 238102 489774 238170
rect 489154 238046 489250 238102
rect 489306 238046 489374 238102
rect 489430 238046 489498 238102
rect 489554 238046 489622 238102
rect 489678 238046 489774 238102
rect 489154 237978 489774 238046
rect 489154 237922 489250 237978
rect 489306 237922 489374 237978
rect 489430 237922 489498 237978
rect 489554 237922 489622 237978
rect 489678 237922 489774 237978
rect 489154 220350 489774 237922
rect 489154 220294 489250 220350
rect 489306 220294 489374 220350
rect 489430 220294 489498 220350
rect 489554 220294 489622 220350
rect 489678 220294 489774 220350
rect 489154 220226 489774 220294
rect 489154 220170 489250 220226
rect 489306 220170 489374 220226
rect 489430 220170 489498 220226
rect 489554 220170 489622 220226
rect 489678 220170 489774 220226
rect 489154 220102 489774 220170
rect 489154 220046 489250 220102
rect 489306 220046 489374 220102
rect 489430 220046 489498 220102
rect 489554 220046 489622 220102
rect 489678 220046 489774 220102
rect 489154 219978 489774 220046
rect 489154 219922 489250 219978
rect 489306 219922 489374 219978
rect 489430 219922 489498 219978
rect 489554 219922 489622 219978
rect 489678 219922 489774 219978
rect 489154 217934 489774 219922
rect 492874 598172 493494 598268
rect 492874 598116 492970 598172
rect 493026 598116 493094 598172
rect 493150 598116 493218 598172
rect 493274 598116 493342 598172
rect 493398 598116 493494 598172
rect 492874 598048 493494 598116
rect 492874 597992 492970 598048
rect 493026 597992 493094 598048
rect 493150 597992 493218 598048
rect 493274 597992 493342 598048
rect 493398 597992 493494 598048
rect 492874 597924 493494 597992
rect 492874 597868 492970 597924
rect 493026 597868 493094 597924
rect 493150 597868 493218 597924
rect 493274 597868 493342 597924
rect 493398 597868 493494 597924
rect 492874 597800 493494 597868
rect 492874 597744 492970 597800
rect 493026 597744 493094 597800
rect 493150 597744 493218 597800
rect 493274 597744 493342 597800
rect 493398 597744 493494 597800
rect 492874 586350 493494 597744
rect 492874 586294 492970 586350
rect 493026 586294 493094 586350
rect 493150 586294 493218 586350
rect 493274 586294 493342 586350
rect 493398 586294 493494 586350
rect 492874 586226 493494 586294
rect 492874 586170 492970 586226
rect 493026 586170 493094 586226
rect 493150 586170 493218 586226
rect 493274 586170 493342 586226
rect 493398 586170 493494 586226
rect 492874 586102 493494 586170
rect 492874 586046 492970 586102
rect 493026 586046 493094 586102
rect 493150 586046 493218 586102
rect 493274 586046 493342 586102
rect 493398 586046 493494 586102
rect 492874 585978 493494 586046
rect 492874 585922 492970 585978
rect 493026 585922 493094 585978
rect 493150 585922 493218 585978
rect 493274 585922 493342 585978
rect 493398 585922 493494 585978
rect 492874 568350 493494 585922
rect 492874 568294 492970 568350
rect 493026 568294 493094 568350
rect 493150 568294 493218 568350
rect 493274 568294 493342 568350
rect 493398 568294 493494 568350
rect 492874 568226 493494 568294
rect 492874 568170 492970 568226
rect 493026 568170 493094 568226
rect 493150 568170 493218 568226
rect 493274 568170 493342 568226
rect 493398 568170 493494 568226
rect 492874 568102 493494 568170
rect 492874 568046 492970 568102
rect 493026 568046 493094 568102
rect 493150 568046 493218 568102
rect 493274 568046 493342 568102
rect 493398 568046 493494 568102
rect 492874 567978 493494 568046
rect 492874 567922 492970 567978
rect 493026 567922 493094 567978
rect 493150 567922 493218 567978
rect 493274 567922 493342 567978
rect 493398 567922 493494 567978
rect 492874 550350 493494 567922
rect 492874 550294 492970 550350
rect 493026 550294 493094 550350
rect 493150 550294 493218 550350
rect 493274 550294 493342 550350
rect 493398 550294 493494 550350
rect 492874 550226 493494 550294
rect 492874 550170 492970 550226
rect 493026 550170 493094 550226
rect 493150 550170 493218 550226
rect 493274 550170 493342 550226
rect 493398 550170 493494 550226
rect 492874 550102 493494 550170
rect 492874 550046 492970 550102
rect 493026 550046 493094 550102
rect 493150 550046 493218 550102
rect 493274 550046 493342 550102
rect 493398 550046 493494 550102
rect 492874 549978 493494 550046
rect 492874 549922 492970 549978
rect 493026 549922 493094 549978
rect 493150 549922 493218 549978
rect 493274 549922 493342 549978
rect 493398 549922 493494 549978
rect 492874 532350 493494 549922
rect 492874 532294 492970 532350
rect 493026 532294 493094 532350
rect 493150 532294 493218 532350
rect 493274 532294 493342 532350
rect 493398 532294 493494 532350
rect 492874 532226 493494 532294
rect 492874 532170 492970 532226
rect 493026 532170 493094 532226
rect 493150 532170 493218 532226
rect 493274 532170 493342 532226
rect 493398 532170 493494 532226
rect 492874 532102 493494 532170
rect 492874 532046 492970 532102
rect 493026 532046 493094 532102
rect 493150 532046 493218 532102
rect 493274 532046 493342 532102
rect 493398 532046 493494 532102
rect 492874 531978 493494 532046
rect 492874 531922 492970 531978
rect 493026 531922 493094 531978
rect 493150 531922 493218 531978
rect 493274 531922 493342 531978
rect 493398 531922 493494 531978
rect 492874 514350 493494 531922
rect 492874 514294 492970 514350
rect 493026 514294 493094 514350
rect 493150 514294 493218 514350
rect 493274 514294 493342 514350
rect 493398 514294 493494 514350
rect 492874 514226 493494 514294
rect 492874 514170 492970 514226
rect 493026 514170 493094 514226
rect 493150 514170 493218 514226
rect 493274 514170 493342 514226
rect 493398 514170 493494 514226
rect 492874 514102 493494 514170
rect 492874 514046 492970 514102
rect 493026 514046 493094 514102
rect 493150 514046 493218 514102
rect 493274 514046 493342 514102
rect 493398 514046 493494 514102
rect 492874 513978 493494 514046
rect 492874 513922 492970 513978
rect 493026 513922 493094 513978
rect 493150 513922 493218 513978
rect 493274 513922 493342 513978
rect 493398 513922 493494 513978
rect 492874 496350 493494 513922
rect 492874 496294 492970 496350
rect 493026 496294 493094 496350
rect 493150 496294 493218 496350
rect 493274 496294 493342 496350
rect 493398 496294 493494 496350
rect 492874 496226 493494 496294
rect 492874 496170 492970 496226
rect 493026 496170 493094 496226
rect 493150 496170 493218 496226
rect 493274 496170 493342 496226
rect 493398 496170 493494 496226
rect 492874 496102 493494 496170
rect 492874 496046 492970 496102
rect 493026 496046 493094 496102
rect 493150 496046 493218 496102
rect 493274 496046 493342 496102
rect 493398 496046 493494 496102
rect 492874 495978 493494 496046
rect 492874 495922 492970 495978
rect 493026 495922 493094 495978
rect 493150 495922 493218 495978
rect 493274 495922 493342 495978
rect 493398 495922 493494 495978
rect 492874 478350 493494 495922
rect 492874 478294 492970 478350
rect 493026 478294 493094 478350
rect 493150 478294 493218 478350
rect 493274 478294 493342 478350
rect 493398 478294 493494 478350
rect 492874 478226 493494 478294
rect 492874 478170 492970 478226
rect 493026 478170 493094 478226
rect 493150 478170 493218 478226
rect 493274 478170 493342 478226
rect 493398 478170 493494 478226
rect 492874 478102 493494 478170
rect 492874 478046 492970 478102
rect 493026 478046 493094 478102
rect 493150 478046 493218 478102
rect 493274 478046 493342 478102
rect 493398 478046 493494 478102
rect 492874 477978 493494 478046
rect 492874 477922 492970 477978
rect 493026 477922 493094 477978
rect 493150 477922 493218 477978
rect 493274 477922 493342 477978
rect 493398 477922 493494 477978
rect 492874 460350 493494 477922
rect 492874 460294 492970 460350
rect 493026 460294 493094 460350
rect 493150 460294 493218 460350
rect 493274 460294 493342 460350
rect 493398 460294 493494 460350
rect 492874 460226 493494 460294
rect 492874 460170 492970 460226
rect 493026 460170 493094 460226
rect 493150 460170 493218 460226
rect 493274 460170 493342 460226
rect 493398 460170 493494 460226
rect 492874 460102 493494 460170
rect 492874 460046 492970 460102
rect 493026 460046 493094 460102
rect 493150 460046 493218 460102
rect 493274 460046 493342 460102
rect 493398 460046 493494 460102
rect 492874 459978 493494 460046
rect 492874 459922 492970 459978
rect 493026 459922 493094 459978
rect 493150 459922 493218 459978
rect 493274 459922 493342 459978
rect 493398 459922 493494 459978
rect 492874 442350 493494 459922
rect 492874 442294 492970 442350
rect 493026 442294 493094 442350
rect 493150 442294 493218 442350
rect 493274 442294 493342 442350
rect 493398 442294 493494 442350
rect 492874 442226 493494 442294
rect 492874 442170 492970 442226
rect 493026 442170 493094 442226
rect 493150 442170 493218 442226
rect 493274 442170 493342 442226
rect 493398 442170 493494 442226
rect 492874 442102 493494 442170
rect 492874 442046 492970 442102
rect 493026 442046 493094 442102
rect 493150 442046 493218 442102
rect 493274 442046 493342 442102
rect 493398 442046 493494 442102
rect 492874 441978 493494 442046
rect 492874 441922 492970 441978
rect 493026 441922 493094 441978
rect 493150 441922 493218 441978
rect 493274 441922 493342 441978
rect 493398 441922 493494 441978
rect 492874 424350 493494 441922
rect 492874 424294 492970 424350
rect 493026 424294 493094 424350
rect 493150 424294 493218 424350
rect 493274 424294 493342 424350
rect 493398 424294 493494 424350
rect 492874 424226 493494 424294
rect 492874 424170 492970 424226
rect 493026 424170 493094 424226
rect 493150 424170 493218 424226
rect 493274 424170 493342 424226
rect 493398 424170 493494 424226
rect 492874 424102 493494 424170
rect 492874 424046 492970 424102
rect 493026 424046 493094 424102
rect 493150 424046 493218 424102
rect 493274 424046 493342 424102
rect 493398 424046 493494 424102
rect 492874 423978 493494 424046
rect 492874 423922 492970 423978
rect 493026 423922 493094 423978
rect 493150 423922 493218 423978
rect 493274 423922 493342 423978
rect 493398 423922 493494 423978
rect 492874 406350 493494 423922
rect 492874 406294 492970 406350
rect 493026 406294 493094 406350
rect 493150 406294 493218 406350
rect 493274 406294 493342 406350
rect 493398 406294 493494 406350
rect 492874 406226 493494 406294
rect 492874 406170 492970 406226
rect 493026 406170 493094 406226
rect 493150 406170 493218 406226
rect 493274 406170 493342 406226
rect 493398 406170 493494 406226
rect 492874 406102 493494 406170
rect 492874 406046 492970 406102
rect 493026 406046 493094 406102
rect 493150 406046 493218 406102
rect 493274 406046 493342 406102
rect 493398 406046 493494 406102
rect 492874 405978 493494 406046
rect 492874 405922 492970 405978
rect 493026 405922 493094 405978
rect 493150 405922 493218 405978
rect 493274 405922 493342 405978
rect 493398 405922 493494 405978
rect 492874 388350 493494 405922
rect 492874 388294 492970 388350
rect 493026 388294 493094 388350
rect 493150 388294 493218 388350
rect 493274 388294 493342 388350
rect 493398 388294 493494 388350
rect 492874 388226 493494 388294
rect 492874 388170 492970 388226
rect 493026 388170 493094 388226
rect 493150 388170 493218 388226
rect 493274 388170 493342 388226
rect 493398 388170 493494 388226
rect 492874 388102 493494 388170
rect 492874 388046 492970 388102
rect 493026 388046 493094 388102
rect 493150 388046 493218 388102
rect 493274 388046 493342 388102
rect 493398 388046 493494 388102
rect 492874 387978 493494 388046
rect 492874 387922 492970 387978
rect 493026 387922 493094 387978
rect 493150 387922 493218 387978
rect 493274 387922 493342 387978
rect 493398 387922 493494 387978
rect 492874 370350 493494 387922
rect 492874 370294 492970 370350
rect 493026 370294 493094 370350
rect 493150 370294 493218 370350
rect 493274 370294 493342 370350
rect 493398 370294 493494 370350
rect 492874 370226 493494 370294
rect 492874 370170 492970 370226
rect 493026 370170 493094 370226
rect 493150 370170 493218 370226
rect 493274 370170 493342 370226
rect 493398 370170 493494 370226
rect 492874 370102 493494 370170
rect 492874 370046 492970 370102
rect 493026 370046 493094 370102
rect 493150 370046 493218 370102
rect 493274 370046 493342 370102
rect 493398 370046 493494 370102
rect 492874 369978 493494 370046
rect 492874 369922 492970 369978
rect 493026 369922 493094 369978
rect 493150 369922 493218 369978
rect 493274 369922 493342 369978
rect 493398 369922 493494 369978
rect 492874 352350 493494 369922
rect 492874 352294 492970 352350
rect 493026 352294 493094 352350
rect 493150 352294 493218 352350
rect 493274 352294 493342 352350
rect 493398 352294 493494 352350
rect 492874 352226 493494 352294
rect 492874 352170 492970 352226
rect 493026 352170 493094 352226
rect 493150 352170 493218 352226
rect 493274 352170 493342 352226
rect 493398 352170 493494 352226
rect 492874 352102 493494 352170
rect 492874 352046 492970 352102
rect 493026 352046 493094 352102
rect 493150 352046 493218 352102
rect 493274 352046 493342 352102
rect 493398 352046 493494 352102
rect 492874 351978 493494 352046
rect 492874 351922 492970 351978
rect 493026 351922 493094 351978
rect 493150 351922 493218 351978
rect 493274 351922 493342 351978
rect 493398 351922 493494 351978
rect 492874 334350 493494 351922
rect 492874 334294 492970 334350
rect 493026 334294 493094 334350
rect 493150 334294 493218 334350
rect 493274 334294 493342 334350
rect 493398 334294 493494 334350
rect 492874 334226 493494 334294
rect 492874 334170 492970 334226
rect 493026 334170 493094 334226
rect 493150 334170 493218 334226
rect 493274 334170 493342 334226
rect 493398 334170 493494 334226
rect 492874 334102 493494 334170
rect 492874 334046 492970 334102
rect 493026 334046 493094 334102
rect 493150 334046 493218 334102
rect 493274 334046 493342 334102
rect 493398 334046 493494 334102
rect 492874 333978 493494 334046
rect 492874 333922 492970 333978
rect 493026 333922 493094 333978
rect 493150 333922 493218 333978
rect 493274 333922 493342 333978
rect 493398 333922 493494 333978
rect 492874 316350 493494 333922
rect 492874 316294 492970 316350
rect 493026 316294 493094 316350
rect 493150 316294 493218 316350
rect 493274 316294 493342 316350
rect 493398 316294 493494 316350
rect 492874 316226 493494 316294
rect 492874 316170 492970 316226
rect 493026 316170 493094 316226
rect 493150 316170 493218 316226
rect 493274 316170 493342 316226
rect 493398 316170 493494 316226
rect 492874 316102 493494 316170
rect 492874 316046 492970 316102
rect 493026 316046 493094 316102
rect 493150 316046 493218 316102
rect 493274 316046 493342 316102
rect 493398 316046 493494 316102
rect 492874 315978 493494 316046
rect 492874 315922 492970 315978
rect 493026 315922 493094 315978
rect 493150 315922 493218 315978
rect 493274 315922 493342 315978
rect 493398 315922 493494 315978
rect 492874 298350 493494 315922
rect 492874 298294 492970 298350
rect 493026 298294 493094 298350
rect 493150 298294 493218 298350
rect 493274 298294 493342 298350
rect 493398 298294 493494 298350
rect 492874 298226 493494 298294
rect 492874 298170 492970 298226
rect 493026 298170 493094 298226
rect 493150 298170 493218 298226
rect 493274 298170 493342 298226
rect 493398 298170 493494 298226
rect 492874 298102 493494 298170
rect 492874 298046 492970 298102
rect 493026 298046 493094 298102
rect 493150 298046 493218 298102
rect 493274 298046 493342 298102
rect 493398 298046 493494 298102
rect 492874 297978 493494 298046
rect 492874 297922 492970 297978
rect 493026 297922 493094 297978
rect 493150 297922 493218 297978
rect 493274 297922 493342 297978
rect 493398 297922 493494 297978
rect 492874 280350 493494 297922
rect 492874 280294 492970 280350
rect 493026 280294 493094 280350
rect 493150 280294 493218 280350
rect 493274 280294 493342 280350
rect 493398 280294 493494 280350
rect 492874 280226 493494 280294
rect 492874 280170 492970 280226
rect 493026 280170 493094 280226
rect 493150 280170 493218 280226
rect 493274 280170 493342 280226
rect 493398 280170 493494 280226
rect 492874 280102 493494 280170
rect 492874 280046 492970 280102
rect 493026 280046 493094 280102
rect 493150 280046 493218 280102
rect 493274 280046 493342 280102
rect 493398 280046 493494 280102
rect 492874 279978 493494 280046
rect 492874 279922 492970 279978
rect 493026 279922 493094 279978
rect 493150 279922 493218 279978
rect 493274 279922 493342 279978
rect 493398 279922 493494 279978
rect 492874 262350 493494 279922
rect 492874 262294 492970 262350
rect 493026 262294 493094 262350
rect 493150 262294 493218 262350
rect 493274 262294 493342 262350
rect 493398 262294 493494 262350
rect 492874 262226 493494 262294
rect 492874 262170 492970 262226
rect 493026 262170 493094 262226
rect 493150 262170 493218 262226
rect 493274 262170 493342 262226
rect 493398 262170 493494 262226
rect 492874 262102 493494 262170
rect 492874 262046 492970 262102
rect 493026 262046 493094 262102
rect 493150 262046 493218 262102
rect 493274 262046 493342 262102
rect 493398 262046 493494 262102
rect 492874 261978 493494 262046
rect 492874 261922 492970 261978
rect 493026 261922 493094 261978
rect 493150 261922 493218 261978
rect 493274 261922 493342 261978
rect 493398 261922 493494 261978
rect 492874 244350 493494 261922
rect 492874 244294 492970 244350
rect 493026 244294 493094 244350
rect 493150 244294 493218 244350
rect 493274 244294 493342 244350
rect 493398 244294 493494 244350
rect 492874 244226 493494 244294
rect 492874 244170 492970 244226
rect 493026 244170 493094 244226
rect 493150 244170 493218 244226
rect 493274 244170 493342 244226
rect 493398 244170 493494 244226
rect 492874 244102 493494 244170
rect 492874 244046 492970 244102
rect 493026 244046 493094 244102
rect 493150 244046 493218 244102
rect 493274 244046 493342 244102
rect 493398 244046 493494 244102
rect 492874 243978 493494 244046
rect 492874 243922 492970 243978
rect 493026 243922 493094 243978
rect 493150 243922 493218 243978
rect 493274 243922 493342 243978
rect 493398 243922 493494 243978
rect 492874 226350 493494 243922
rect 492874 226294 492970 226350
rect 493026 226294 493094 226350
rect 493150 226294 493218 226350
rect 493274 226294 493342 226350
rect 493398 226294 493494 226350
rect 492874 226226 493494 226294
rect 492874 226170 492970 226226
rect 493026 226170 493094 226226
rect 493150 226170 493218 226226
rect 493274 226170 493342 226226
rect 493398 226170 493494 226226
rect 492874 226102 493494 226170
rect 492874 226046 492970 226102
rect 493026 226046 493094 226102
rect 493150 226046 493218 226102
rect 493274 226046 493342 226102
rect 493398 226046 493494 226102
rect 492874 225978 493494 226046
rect 492874 225922 492970 225978
rect 493026 225922 493094 225978
rect 493150 225922 493218 225978
rect 493274 225922 493342 225978
rect 493398 225922 493494 225978
rect 492874 217934 493494 225922
rect 507154 597212 507774 598268
rect 507154 597156 507250 597212
rect 507306 597156 507374 597212
rect 507430 597156 507498 597212
rect 507554 597156 507622 597212
rect 507678 597156 507774 597212
rect 507154 597088 507774 597156
rect 507154 597032 507250 597088
rect 507306 597032 507374 597088
rect 507430 597032 507498 597088
rect 507554 597032 507622 597088
rect 507678 597032 507774 597088
rect 507154 596964 507774 597032
rect 507154 596908 507250 596964
rect 507306 596908 507374 596964
rect 507430 596908 507498 596964
rect 507554 596908 507622 596964
rect 507678 596908 507774 596964
rect 507154 596840 507774 596908
rect 507154 596784 507250 596840
rect 507306 596784 507374 596840
rect 507430 596784 507498 596840
rect 507554 596784 507622 596840
rect 507678 596784 507774 596840
rect 507154 580350 507774 596784
rect 507154 580294 507250 580350
rect 507306 580294 507374 580350
rect 507430 580294 507498 580350
rect 507554 580294 507622 580350
rect 507678 580294 507774 580350
rect 507154 580226 507774 580294
rect 507154 580170 507250 580226
rect 507306 580170 507374 580226
rect 507430 580170 507498 580226
rect 507554 580170 507622 580226
rect 507678 580170 507774 580226
rect 507154 580102 507774 580170
rect 507154 580046 507250 580102
rect 507306 580046 507374 580102
rect 507430 580046 507498 580102
rect 507554 580046 507622 580102
rect 507678 580046 507774 580102
rect 507154 579978 507774 580046
rect 507154 579922 507250 579978
rect 507306 579922 507374 579978
rect 507430 579922 507498 579978
rect 507554 579922 507622 579978
rect 507678 579922 507774 579978
rect 507154 562350 507774 579922
rect 507154 562294 507250 562350
rect 507306 562294 507374 562350
rect 507430 562294 507498 562350
rect 507554 562294 507622 562350
rect 507678 562294 507774 562350
rect 507154 562226 507774 562294
rect 507154 562170 507250 562226
rect 507306 562170 507374 562226
rect 507430 562170 507498 562226
rect 507554 562170 507622 562226
rect 507678 562170 507774 562226
rect 507154 562102 507774 562170
rect 507154 562046 507250 562102
rect 507306 562046 507374 562102
rect 507430 562046 507498 562102
rect 507554 562046 507622 562102
rect 507678 562046 507774 562102
rect 507154 561978 507774 562046
rect 507154 561922 507250 561978
rect 507306 561922 507374 561978
rect 507430 561922 507498 561978
rect 507554 561922 507622 561978
rect 507678 561922 507774 561978
rect 507154 544350 507774 561922
rect 507154 544294 507250 544350
rect 507306 544294 507374 544350
rect 507430 544294 507498 544350
rect 507554 544294 507622 544350
rect 507678 544294 507774 544350
rect 507154 544226 507774 544294
rect 507154 544170 507250 544226
rect 507306 544170 507374 544226
rect 507430 544170 507498 544226
rect 507554 544170 507622 544226
rect 507678 544170 507774 544226
rect 507154 544102 507774 544170
rect 507154 544046 507250 544102
rect 507306 544046 507374 544102
rect 507430 544046 507498 544102
rect 507554 544046 507622 544102
rect 507678 544046 507774 544102
rect 507154 543978 507774 544046
rect 507154 543922 507250 543978
rect 507306 543922 507374 543978
rect 507430 543922 507498 543978
rect 507554 543922 507622 543978
rect 507678 543922 507774 543978
rect 507154 526350 507774 543922
rect 507154 526294 507250 526350
rect 507306 526294 507374 526350
rect 507430 526294 507498 526350
rect 507554 526294 507622 526350
rect 507678 526294 507774 526350
rect 507154 526226 507774 526294
rect 507154 526170 507250 526226
rect 507306 526170 507374 526226
rect 507430 526170 507498 526226
rect 507554 526170 507622 526226
rect 507678 526170 507774 526226
rect 507154 526102 507774 526170
rect 507154 526046 507250 526102
rect 507306 526046 507374 526102
rect 507430 526046 507498 526102
rect 507554 526046 507622 526102
rect 507678 526046 507774 526102
rect 507154 525978 507774 526046
rect 507154 525922 507250 525978
rect 507306 525922 507374 525978
rect 507430 525922 507498 525978
rect 507554 525922 507622 525978
rect 507678 525922 507774 525978
rect 507154 508350 507774 525922
rect 507154 508294 507250 508350
rect 507306 508294 507374 508350
rect 507430 508294 507498 508350
rect 507554 508294 507622 508350
rect 507678 508294 507774 508350
rect 507154 508226 507774 508294
rect 507154 508170 507250 508226
rect 507306 508170 507374 508226
rect 507430 508170 507498 508226
rect 507554 508170 507622 508226
rect 507678 508170 507774 508226
rect 507154 508102 507774 508170
rect 507154 508046 507250 508102
rect 507306 508046 507374 508102
rect 507430 508046 507498 508102
rect 507554 508046 507622 508102
rect 507678 508046 507774 508102
rect 507154 507978 507774 508046
rect 507154 507922 507250 507978
rect 507306 507922 507374 507978
rect 507430 507922 507498 507978
rect 507554 507922 507622 507978
rect 507678 507922 507774 507978
rect 507154 490350 507774 507922
rect 507154 490294 507250 490350
rect 507306 490294 507374 490350
rect 507430 490294 507498 490350
rect 507554 490294 507622 490350
rect 507678 490294 507774 490350
rect 507154 490226 507774 490294
rect 507154 490170 507250 490226
rect 507306 490170 507374 490226
rect 507430 490170 507498 490226
rect 507554 490170 507622 490226
rect 507678 490170 507774 490226
rect 507154 490102 507774 490170
rect 507154 490046 507250 490102
rect 507306 490046 507374 490102
rect 507430 490046 507498 490102
rect 507554 490046 507622 490102
rect 507678 490046 507774 490102
rect 507154 489978 507774 490046
rect 507154 489922 507250 489978
rect 507306 489922 507374 489978
rect 507430 489922 507498 489978
rect 507554 489922 507622 489978
rect 507678 489922 507774 489978
rect 507154 472350 507774 489922
rect 507154 472294 507250 472350
rect 507306 472294 507374 472350
rect 507430 472294 507498 472350
rect 507554 472294 507622 472350
rect 507678 472294 507774 472350
rect 507154 472226 507774 472294
rect 507154 472170 507250 472226
rect 507306 472170 507374 472226
rect 507430 472170 507498 472226
rect 507554 472170 507622 472226
rect 507678 472170 507774 472226
rect 507154 472102 507774 472170
rect 507154 472046 507250 472102
rect 507306 472046 507374 472102
rect 507430 472046 507498 472102
rect 507554 472046 507622 472102
rect 507678 472046 507774 472102
rect 507154 471978 507774 472046
rect 507154 471922 507250 471978
rect 507306 471922 507374 471978
rect 507430 471922 507498 471978
rect 507554 471922 507622 471978
rect 507678 471922 507774 471978
rect 507154 454350 507774 471922
rect 507154 454294 507250 454350
rect 507306 454294 507374 454350
rect 507430 454294 507498 454350
rect 507554 454294 507622 454350
rect 507678 454294 507774 454350
rect 507154 454226 507774 454294
rect 507154 454170 507250 454226
rect 507306 454170 507374 454226
rect 507430 454170 507498 454226
rect 507554 454170 507622 454226
rect 507678 454170 507774 454226
rect 507154 454102 507774 454170
rect 507154 454046 507250 454102
rect 507306 454046 507374 454102
rect 507430 454046 507498 454102
rect 507554 454046 507622 454102
rect 507678 454046 507774 454102
rect 507154 453978 507774 454046
rect 507154 453922 507250 453978
rect 507306 453922 507374 453978
rect 507430 453922 507498 453978
rect 507554 453922 507622 453978
rect 507678 453922 507774 453978
rect 507154 436350 507774 453922
rect 507154 436294 507250 436350
rect 507306 436294 507374 436350
rect 507430 436294 507498 436350
rect 507554 436294 507622 436350
rect 507678 436294 507774 436350
rect 507154 436226 507774 436294
rect 507154 436170 507250 436226
rect 507306 436170 507374 436226
rect 507430 436170 507498 436226
rect 507554 436170 507622 436226
rect 507678 436170 507774 436226
rect 507154 436102 507774 436170
rect 507154 436046 507250 436102
rect 507306 436046 507374 436102
rect 507430 436046 507498 436102
rect 507554 436046 507622 436102
rect 507678 436046 507774 436102
rect 507154 435978 507774 436046
rect 507154 435922 507250 435978
rect 507306 435922 507374 435978
rect 507430 435922 507498 435978
rect 507554 435922 507622 435978
rect 507678 435922 507774 435978
rect 507154 418350 507774 435922
rect 507154 418294 507250 418350
rect 507306 418294 507374 418350
rect 507430 418294 507498 418350
rect 507554 418294 507622 418350
rect 507678 418294 507774 418350
rect 507154 418226 507774 418294
rect 507154 418170 507250 418226
rect 507306 418170 507374 418226
rect 507430 418170 507498 418226
rect 507554 418170 507622 418226
rect 507678 418170 507774 418226
rect 507154 418102 507774 418170
rect 507154 418046 507250 418102
rect 507306 418046 507374 418102
rect 507430 418046 507498 418102
rect 507554 418046 507622 418102
rect 507678 418046 507774 418102
rect 507154 417978 507774 418046
rect 507154 417922 507250 417978
rect 507306 417922 507374 417978
rect 507430 417922 507498 417978
rect 507554 417922 507622 417978
rect 507678 417922 507774 417978
rect 507154 400350 507774 417922
rect 507154 400294 507250 400350
rect 507306 400294 507374 400350
rect 507430 400294 507498 400350
rect 507554 400294 507622 400350
rect 507678 400294 507774 400350
rect 507154 400226 507774 400294
rect 507154 400170 507250 400226
rect 507306 400170 507374 400226
rect 507430 400170 507498 400226
rect 507554 400170 507622 400226
rect 507678 400170 507774 400226
rect 507154 400102 507774 400170
rect 507154 400046 507250 400102
rect 507306 400046 507374 400102
rect 507430 400046 507498 400102
rect 507554 400046 507622 400102
rect 507678 400046 507774 400102
rect 507154 399978 507774 400046
rect 507154 399922 507250 399978
rect 507306 399922 507374 399978
rect 507430 399922 507498 399978
rect 507554 399922 507622 399978
rect 507678 399922 507774 399978
rect 507154 382350 507774 399922
rect 507154 382294 507250 382350
rect 507306 382294 507374 382350
rect 507430 382294 507498 382350
rect 507554 382294 507622 382350
rect 507678 382294 507774 382350
rect 507154 382226 507774 382294
rect 507154 382170 507250 382226
rect 507306 382170 507374 382226
rect 507430 382170 507498 382226
rect 507554 382170 507622 382226
rect 507678 382170 507774 382226
rect 507154 382102 507774 382170
rect 507154 382046 507250 382102
rect 507306 382046 507374 382102
rect 507430 382046 507498 382102
rect 507554 382046 507622 382102
rect 507678 382046 507774 382102
rect 507154 381978 507774 382046
rect 507154 381922 507250 381978
rect 507306 381922 507374 381978
rect 507430 381922 507498 381978
rect 507554 381922 507622 381978
rect 507678 381922 507774 381978
rect 507154 364350 507774 381922
rect 507154 364294 507250 364350
rect 507306 364294 507374 364350
rect 507430 364294 507498 364350
rect 507554 364294 507622 364350
rect 507678 364294 507774 364350
rect 507154 364226 507774 364294
rect 507154 364170 507250 364226
rect 507306 364170 507374 364226
rect 507430 364170 507498 364226
rect 507554 364170 507622 364226
rect 507678 364170 507774 364226
rect 507154 364102 507774 364170
rect 507154 364046 507250 364102
rect 507306 364046 507374 364102
rect 507430 364046 507498 364102
rect 507554 364046 507622 364102
rect 507678 364046 507774 364102
rect 507154 363978 507774 364046
rect 507154 363922 507250 363978
rect 507306 363922 507374 363978
rect 507430 363922 507498 363978
rect 507554 363922 507622 363978
rect 507678 363922 507774 363978
rect 507154 346350 507774 363922
rect 507154 346294 507250 346350
rect 507306 346294 507374 346350
rect 507430 346294 507498 346350
rect 507554 346294 507622 346350
rect 507678 346294 507774 346350
rect 507154 346226 507774 346294
rect 507154 346170 507250 346226
rect 507306 346170 507374 346226
rect 507430 346170 507498 346226
rect 507554 346170 507622 346226
rect 507678 346170 507774 346226
rect 507154 346102 507774 346170
rect 507154 346046 507250 346102
rect 507306 346046 507374 346102
rect 507430 346046 507498 346102
rect 507554 346046 507622 346102
rect 507678 346046 507774 346102
rect 507154 345978 507774 346046
rect 507154 345922 507250 345978
rect 507306 345922 507374 345978
rect 507430 345922 507498 345978
rect 507554 345922 507622 345978
rect 507678 345922 507774 345978
rect 507154 328350 507774 345922
rect 507154 328294 507250 328350
rect 507306 328294 507374 328350
rect 507430 328294 507498 328350
rect 507554 328294 507622 328350
rect 507678 328294 507774 328350
rect 507154 328226 507774 328294
rect 507154 328170 507250 328226
rect 507306 328170 507374 328226
rect 507430 328170 507498 328226
rect 507554 328170 507622 328226
rect 507678 328170 507774 328226
rect 507154 328102 507774 328170
rect 507154 328046 507250 328102
rect 507306 328046 507374 328102
rect 507430 328046 507498 328102
rect 507554 328046 507622 328102
rect 507678 328046 507774 328102
rect 507154 327978 507774 328046
rect 507154 327922 507250 327978
rect 507306 327922 507374 327978
rect 507430 327922 507498 327978
rect 507554 327922 507622 327978
rect 507678 327922 507774 327978
rect 507154 310350 507774 327922
rect 507154 310294 507250 310350
rect 507306 310294 507374 310350
rect 507430 310294 507498 310350
rect 507554 310294 507622 310350
rect 507678 310294 507774 310350
rect 507154 310226 507774 310294
rect 507154 310170 507250 310226
rect 507306 310170 507374 310226
rect 507430 310170 507498 310226
rect 507554 310170 507622 310226
rect 507678 310170 507774 310226
rect 507154 310102 507774 310170
rect 507154 310046 507250 310102
rect 507306 310046 507374 310102
rect 507430 310046 507498 310102
rect 507554 310046 507622 310102
rect 507678 310046 507774 310102
rect 507154 309978 507774 310046
rect 507154 309922 507250 309978
rect 507306 309922 507374 309978
rect 507430 309922 507498 309978
rect 507554 309922 507622 309978
rect 507678 309922 507774 309978
rect 507154 292350 507774 309922
rect 507154 292294 507250 292350
rect 507306 292294 507374 292350
rect 507430 292294 507498 292350
rect 507554 292294 507622 292350
rect 507678 292294 507774 292350
rect 507154 292226 507774 292294
rect 507154 292170 507250 292226
rect 507306 292170 507374 292226
rect 507430 292170 507498 292226
rect 507554 292170 507622 292226
rect 507678 292170 507774 292226
rect 507154 292102 507774 292170
rect 507154 292046 507250 292102
rect 507306 292046 507374 292102
rect 507430 292046 507498 292102
rect 507554 292046 507622 292102
rect 507678 292046 507774 292102
rect 507154 291978 507774 292046
rect 507154 291922 507250 291978
rect 507306 291922 507374 291978
rect 507430 291922 507498 291978
rect 507554 291922 507622 291978
rect 507678 291922 507774 291978
rect 507154 274350 507774 291922
rect 507154 274294 507250 274350
rect 507306 274294 507374 274350
rect 507430 274294 507498 274350
rect 507554 274294 507622 274350
rect 507678 274294 507774 274350
rect 507154 274226 507774 274294
rect 507154 274170 507250 274226
rect 507306 274170 507374 274226
rect 507430 274170 507498 274226
rect 507554 274170 507622 274226
rect 507678 274170 507774 274226
rect 507154 274102 507774 274170
rect 507154 274046 507250 274102
rect 507306 274046 507374 274102
rect 507430 274046 507498 274102
rect 507554 274046 507622 274102
rect 507678 274046 507774 274102
rect 507154 273978 507774 274046
rect 507154 273922 507250 273978
rect 507306 273922 507374 273978
rect 507430 273922 507498 273978
rect 507554 273922 507622 273978
rect 507678 273922 507774 273978
rect 507154 256350 507774 273922
rect 507154 256294 507250 256350
rect 507306 256294 507374 256350
rect 507430 256294 507498 256350
rect 507554 256294 507622 256350
rect 507678 256294 507774 256350
rect 507154 256226 507774 256294
rect 507154 256170 507250 256226
rect 507306 256170 507374 256226
rect 507430 256170 507498 256226
rect 507554 256170 507622 256226
rect 507678 256170 507774 256226
rect 507154 256102 507774 256170
rect 507154 256046 507250 256102
rect 507306 256046 507374 256102
rect 507430 256046 507498 256102
rect 507554 256046 507622 256102
rect 507678 256046 507774 256102
rect 507154 255978 507774 256046
rect 507154 255922 507250 255978
rect 507306 255922 507374 255978
rect 507430 255922 507498 255978
rect 507554 255922 507622 255978
rect 507678 255922 507774 255978
rect 507154 238350 507774 255922
rect 507154 238294 507250 238350
rect 507306 238294 507374 238350
rect 507430 238294 507498 238350
rect 507554 238294 507622 238350
rect 507678 238294 507774 238350
rect 507154 238226 507774 238294
rect 507154 238170 507250 238226
rect 507306 238170 507374 238226
rect 507430 238170 507498 238226
rect 507554 238170 507622 238226
rect 507678 238170 507774 238226
rect 507154 238102 507774 238170
rect 507154 238046 507250 238102
rect 507306 238046 507374 238102
rect 507430 238046 507498 238102
rect 507554 238046 507622 238102
rect 507678 238046 507774 238102
rect 507154 237978 507774 238046
rect 507154 237922 507250 237978
rect 507306 237922 507374 237978
rect 507430 237922 507498 237978
rect 507554 237922 507622 237978
rect 507678 237922 507774 237978
rect 507154 220350 507774 237922
rect 507154 220294 507250 220350
rect 507306 220294 507374 220350
rect 507430 220294 507498 220350
rect 507554 220294 507622 220350
rect 507678 220294 507774 220350
rect 507154 220226 507774 220294
rect 507154 220170 507250 220226
rect 507306 220170 507374 220226
rect 507430 220170 507498 220226
rect 507554 220170 507622 220226
rect 507678 220170 507774 220226
rect 507154 220102 507774 220170
rect 507154 220046 507250 220102
rect 507306 220046 507374 220102
rect 507430 220046 507498 220102
rect 507554 220046 507622 220102
rect 507678 220046 507774 220102
rect 507154 219978 507774 220046
rect 507154 219922 507250 219978
rect 507306 219922 507374 219978
rect 507430 219922 507498 219978
rect 507554 219922 507622 219978
rect 507678 219922 507774 219978
rect 507154 217934 507774 219922
rect 510874 598172 511494 598268
rect 510874 598116 510970 598172
rect 511026 598116 511094 598172
rect 511150 598116 511218 598172
rect 511274 598116 511342 598172
rect 511398 598116 511494 598172
rect 510874 598048 511494 598116
rect 510874 597992 510970 598048
rect 511026 597992 511094 598048
rect 511150 597992 511218 598048
rect 511274 597992 511342 598048
rect 511398 597992 511494 598048
rect 510874 597924 511494 597992
rect 510874 597868 510970 597924
rect 511026 597868 511094 597924
rect 511150 597868 511218 597924
rect 511274 597868 511342 597924
rect 511398 597868 511494 597924
rect 510874 597800 511494 597868
rect 510874 597744 510970 597800
rect 511026 597744 511094 597800
rect 511150 597744 511218 597800
rect 511274 597744 511342 597800
rect 511398 597744 511494 597800
rect 510874 586350 511494 597744
rect 510874 586294 510970 586350
rect 511026 586294 511094 586350
rect 511150 586294 511218 586350
rect 511274 586294 511342 586350
rect 511398 586294 511494 586350
rect 510874 586226 511494 586294
rect 510874 586170 510970 586226
rect 511026 586170 511094 586226
rect 511150 586170 511218 586226
rect 511274 586170 511342 586226
rect 511398 586170 511494 586226
rect 510874 586102 511494 586170
rect 510874 586046 510970 586102
rect 511026 586046 511094 586102
rect 511150 586046 511218 586102
rect 511274 586046 511342 586102
rect 511398 586046 511494 586102
rect 510874 585978 511494 586046
rect 510874 585922 510970 585978
rect 511026 585922 511094 585978
rect 511150 585922 511218 585978
rect 511274 585922 511342 585978
rect 511398 585922 511494 585978
rect 510874 568350 511494 585922
rect 510874 568294 510970 568350
rect 511026 568294 511094 568350
rect 511150 568294 511218 568350
rect 511274 568294 511342 568350
rect 511398 568294 511494 568350
rect 510874 568226 511494 568294
rect 510874 568170 510970 568226
rect 511026 568170 511094 568226
rect 511150 568170 511218 568226
rect 511274 568170 511342 568226
rect 511398 568170 511494 568226
rect 510874 568102 511494 568170
rect 510874 568046 510970 568102
rect 511026 568046 511094 568102
rect 511150 568046 511218 568102
rect 511274 568046 511342 568102
rect 511398 568046 511494 568102
rect 510874 567978 511494 568046
rect 510874 567922 510970 567978
rect 511026 567922 511094 567978
rect 511150 567922 511218 567978
rect 511274 567922 511342 567978
rect 511398 567922 511494 567978
rect 510874 550350 511494 567922
rect 510874 550294 510970 550350
rect 511026 550294 511094 550350
rect 511150 550294 511218 550350
rect 511274 550294 511342 550350
rect 511398 550294 511494 550350
rect 510874 550226 511494 550294
rect 510874 550170 510970 550226
rect 511026 550170 511094 550226
rect 511150 550170 511218 550226
rect 511274 550170 511342 550226
rect 511398 550170 511494 550226
rect 510874 550102 511494 550170
rect 510874 550046 510970 550102
rect 511026 550046 511094 550102
rect 511150 550046 511218 550102
rect 511274 550046 511342 550102
rect 511398 550046 511494 550102
rect 510874 549978 511494 550046
rect 510874 549922 510970 549978
rect 511026 549922 511094 549978
rect 511150 549922 511218 549978
rect 511274 549922 511342 549978
rect 511398 549922 511494 549978
rect 510874 532350 511494 549922
rect 510874 532294 510970 532350
rect 511026 532294 511094 532350
rect 511150 532294 511218 532350
rect 511274 532294 511342 532350
rect 511398 532294 511494 532350
rect 510874 532226 511494 532294
rect 510874 532170 510970 532226
rect 511026 532170 511094 532226
rect 511150 532170 511218 532226
rect 511274 532170 511342 532226
rect 511398 532170 511494 532226
rect 510874 532102 511494 532170
rect 510874 532046 510970 532102
rect 511026 532046 511094 532102
rect 511150 532046 511218 532102
rect 511274 532046 511342 532102
rect 511398 532046 511494 532102
rect 510874 531978 511494 532046
rect 510874 531922 510970 531978
rect 511026 531922 511094 531978
rect 511150 531922 511218 531978
rect 511274 531922 511342 531978
rect 511398 531922 511494 531978
rect 510874 514350 511494 531922
rect 510874 514294 510970 514350
rect 511026 514294 511094 514350
rect 511150 514294 511218 514350
rect 511274 514294 511342 514350
rect 511398 514294 511494 514350
rect 510874 514226 511494 514294
rect 510874 514170 510970 514226
rect 511026 514170 511094 514226
rect 511150 514170 511218 514226
rect 511274 514170 511342 514226
rect 511398 514170 511494 514226
rect 510874 514102 511494 514170
rect 510874 514046 510970 514102
rect 511026 514046 511094 514102
rect 511150 514046 511218 514102
rect 511274 514046 511342 514102
rect 511398 514046 511494 514102
rect 510874 513978 511494 514046
rect 510874 513922 510970 513978
rect 511026 513922 511094 513978
rect 511150 513922 511218 513978
rect 511274 513922 511342 513978
rect 511398 513922 511494 513978
rect 510874 496350 511494 513922
rect 510874 496294 510970 496350
rect 511026 496294 511094 496350
rect 511150 496294 511218 496350
rect 511274 496294 511342 496350
rect 511398 496294 511494 496350
rect 510874 496226 511494 496294
rect 510874 496170 510970 496226
rect 511026 496170 511094 496226
rect 511150 496170 511218 496226
rect 511274 496170 511342 496226
rect 511398 496170 511494 496226
rect 510874 496102 511494 496170
rect 510874 496046 510970 496102
rect 511026 496046 511094 496102
rect 511150 496046 511218 496102
rect 511274 496046 511342 496102
rect 511398 496046 511494 496102
rect 510874 495978 511494 496046
rect 510874 495922 510970 495978
rect 511026 495922 511094 495978
rect 511150 495922 511218 495978
rect 511274 495922 511342 495978
rect 511398 495922 511494 495978
rect 510874 478350 511494 495922
rect 510874 478294 510970 478350
rect 511026 478294 511094 478350
rect 511150 478294 511218 478350
rect 511274 478294 511342 478350
rect 511398 478294 511494 478350
rect 510874 478226 511494 478294
rect 510874 478170 510970 478226
rect 511026 478170 511094 478226
rect 511150 478170 511218 478226
rect 511274 478170 511342 478226
rect 511398 478170 511494 478226
rect 510874 478102 511494 478170
rect 510874 478046 510970 478102
rect 511026 478046 511094 478102
rect 511150 478046 511218 478102
rect 511274 478046 511342 478102
rect 511398 478046 511494 478102
rect 510874 477978 511494 478046
rect 510874 477922 510970 477978
rect 511026 477922 511094 477978
rect 511150 477922 511218 477978
rect 511274 477922 511342 477978
rect 511398 477922 511494 477978
rect 510874 460350 511494 477922
rect 510874 460294 510970 460350
rect 511026 460294 511094 460350
rect 511150 460294 511218 460350
rect 511274 460294 511342 460350
rect 511398 460294 511494 460350
rect 510874 460226 511494 460294
rect 510874 460170 510970 460226
rect 511026 460170 511094 460226
rect 511150 460170 511218 460226
rect 511274 460170 511342 460226
rect 511398 460170 511494 460226
rect 510874 460102 511494 460170
rect 510874 460046 510970 460102
rect 511026 460046 511094 460102
rect 511150 460046 511218 460102
rect 511274 460046 511342 460102
rect 511398 460046 511494 460102
rect 510874 459978 511494 460046
rect 510874 459922 510970 459978
rect 511026 459922 511094 459978
rect 511150 459922 511218 459978
rect 511274 459922 511342 459978
rect 511398 459922 511494 459978
rect 510874 442350 511494 459922
rect 510874 442294 510970 442350
rect 511026 442294 511094 442350
rect 511150 442294 511218 442350
rect 511274 442294 511342 442350
rect 511398 442294 511494 442350
rect 510874 442226 511494 442294
rect 510874 442170 510970 442226
rect 511026 442170 511094 442226
rect 511150 442170 511218 442226
rect 511274 442170 511342 442226
rect 511398 442170 511494 442226
rect 510874 442102 511494 442170
rect 510874 442046 510970 442102
rect 511026 442046 511094 442102
rect 511150 442046 511218 442102
rect 511274 442046 511342 442102
rect 511398 442046 511494 442102
rect 510874 441978 511494 442046
rect 510874 441922 510970 441978
rect 511026 441922 511094 441978
rect 511150 441922 511218 441978
rect 511274 441922 511342 441978
rect 511398 441922 511494 441978
rect 510874 424350 511494 441922
rect 510874 424294 510970 424350
rect 511026 424294 511094 424350
rect 511150 424294 511218 424350
rect 511274 424294 511342 424350
rect 511398 424294 511494 424350
rect 510874 424226 511494 424294
rect 510874 424170 510970 424226
rect 511026 424170 511094 424226
rect 511150 424170 511218 424226
rect 511274 424170 511342 424226
rect 511398 424170 511494 424226
rect 510874 424102 511494 424170
rect 510874 424046 510970 424102
rect 511026 424046 511094 424102
rect 511150 424046 511218 424102
rect 511274 424046 511342 424102
rect 511398 424046 511494 424102
rect 510874 423978 511494 424046
rect 510874 423922 510970 423978
rect 511026 423922 511094 423978
rect 511150 423922 511218 423978
rect 511274 423922 511342 423978
rect 511398 423922 511494 423978
rect 510874 406350 511494 423922
rect 510874 406294 510970 406350
rect 511026 406294 511094 406350
rect 511150 406294 511218 406350
rect 511274 406294 511342 406350
rect 511398 406294 511494 406350
rect 510874 406226 511494 406294
rect 510874 406170 510970 406226
rect 511026 406170 511094 406226
rect 511150 406170 511218 406226
rect 511274 406170 511342 406226
rect 511398 406170 511494 406226
rect 510874 406102 511494 406170
rect 510874 406046 510970 406102
rect 511026 406046 511094 406102
rect 511150 406046 511218 406102
rect 511274 406046 511342 406102
rect 511398 406046 511494 406102
rect 510874 405978 511494 406046
rect 510874 405922 510970 405978
rect 511026 405922 511094 405978
rect 511150 405922 511218 405978
rect 511274 405922 511342 405978
rect 511398 405922 511494 405978
rect 510874 388350 511494 405922
rect 510874 388294 510970 388350
rect 511026 388294 511094 388350
rect 511150 388294 511218 388350
rect 511274 388294 511342 388350
rect 511398 388294 511494 388350
rect 510874 388226 511494 388294
rect 510874 388170 510970 388226
rect 511026 388170 511094 388226
rect 511150 388170 511218 388226
rect 511274 388170 511342 388226
rect 511398 388170 511494 388226
rect 510874 388102 511494 388170
rect 510874 388046 510970 388102
rect 511026 388046 511094 388102
rect 511150 388046 511218 388102
rect 511274 388046 511342 388102
rect 511398 388046 511494 388102
rect 510874 387978 511494 388046
rect 510874 387922 510970 387978
rect 511026 387922 511094 387978
rect 511150 387922 511218 387978
rect 511274 387922 511342 387978
rect 511398 387922 511494 387978
rect 510874 370350 511494 387922
rect 510874 370294 510970 370350
rect 511026 370294 511094 370350
rect 511150 370294 511218 370350
rect 511274 370294 511342 370350
rect 511398 370294 511494 370350
rect 510874 370226 511494 370294
rect 510874 370170 510970 370226
rect 511026 370170 511094 370226
rect 511150 370170 511218 370226
rect 511274 370170 511342 370226
rect 511398 370170 511494 370226
rect 510874 370102 511494 370170
rect 510874 370046 510970 370102
rect 511026 370046 511094 370102
rect 511150 370046 511218 370102
rect 511274 370046 511342 370102
rect 511398 370046 511494 370102
rect 510874 369978 511494 370046
rect 510874 369922 510970 369978
rect 511026 369922 511094 369978
rect 511150 369922 511218 369978
rect 511274 369922 511342 369978
rect 511398 369922 511494 369978
rect 510874 352350 511494 369922
rect 510874 352294 510970 352350
rect 511026 352294 511094 352350
rect 511150 352294 511218 352350
rect 511274 352294 511342 352350
rect 511398 352294 511494 352350
rect 510874 352226 511494 352294
rect 510874 352170 510970 352226
rect 511026 352170 511094 352226
rect 511150 352170 511218 352226
rect 511274 352170 511342 352226
rect 511398 352170 511494 352226
rect 510874 352102 511494 352170
rect 510874 352046 510970 352102
rect 511026 352046 511094 352102
rect 511150 352046 511218 352102
rect 511274 352046 511342 352102
rect 511398 352046 511494 352102
rect 510874 351978 511494 352046
rect 510874 351922 510970 351978
rect 511026 351922 511094 351978
rect 511150 351922 511218 351978
rect 511274 351922 511342 351978
rect 511398 351922 511494 351978
rect 510874 334350 511494 351922
rect 510874 334294 510970 334350
rect 511026 334294 511094 334350
rect 511150 334294 511218 334350
rect 511274 334294 511342 334350
rect 511398 334294 511494 334350
rect 510874 334226 511494 334294
rect 510874 334170 510970 334226
rect 511026 334170 511094 334226
rect 511150 334170 511218 334226
rect 511274 334170 511342 334226
rect 511398 334170 511494 334226
rect 510874 334102 511494 334170
rect 510874 334046 510970 334102
rect 511026 334046 511094 334102
rect 511150 334046 511218 334102
rect 511274 334046 511342 334102
rect 511398 334046 511494 334102
rect 510874 333978 511494 334046
rect 510874 333922 510970 333978
rect 511026 333922 511094 333978
rect 511150 333922 511218 333978
rect 511274 333922 511342 333978
rect 511398 333922 511494 333978
rect 510874 316350 511494 333922
rect 510874 316294 510970 316350
rect 511026 316294 511094 316350
rect 511150 316294 511218 316350
rect 511274 316294 511342 316350
rect 511398 316294 511494 316350
rect 510874 316226 511494 316294
rect 510874 316170 510970 316226
rect 511026 316170 511094 316226
rect 511150 316170 511218 316226
rect 511274 316170 511342 316226
rect 511398 316170 511494 316226
rect 510874 316102 511494 316170
rect 510874 316046 510970 316102
rect 511026 316046 511094 316102
rect 511150 316046 511218 316102
rect 511274 316046 511342 316102
rect 511398 316046 511494 316102
rect 510874 315978 511494 316046
rect 510874 315922 510970 315978
rect 511026 315922 511094 315978
rect 511150 315922 511218 315978
rect 511274 315922 511342 315978
rect 511398 315922 511494 315978
rect 510874 298350 511494 315922
rect 510874 298294 510970 298350
rect 511026 298294 511094 298350
rect 511150 298294 511218 298350
rect 511274 298294 511342 298350
rect 511398 298294 511494 298350
rect 510874 298226 511494 298294
rect 510874 298170 510970 298226
rect 511026 298170 511094 298226
rect 511150 298170 511218 298226
rect 511274 298170 511342 298226
rect 511398 298170 511494 298226
rect 510874 298102 511494 298170
rect 510874 298046 510970 298102
rect 511026 298046 511094 298102
rect 511150 298046 511218 298102
rect 511274 298046 511342 298102
rect 511398 298046 511494 298102
rect 510874 297978 511494 298046
rect 510874 297922 510970 297978
rect 511026 297922 511094 297978
rect 511150 297922 511218 297978
rect 511274 297922 511342 297978
rect 511398 297922 511494 297978
rect 510874 280350 511494 297922
rect 510874 280294 510970 280350
rect 511026 280294 511094 280350
rect 511150 280294 511218 280350
rect 511274 280294 511342 280350
rect 511398 280294 511494 280350
rect 510874 280226 511494 280294
rect 510874 280170 510970 280226
rect 511026 280170 511094 280226
rect 511150 280170 511218 280226
rect 511274 280170 511342 280226
rect 511398 280170 511494 280226
rect 510874 280102 511494 280170
rect 510874 280046 510970 280102
rect 511026 280046 511094 280102
rect 511150 280046 511218 280102
rect 511274 280046 511342 280102
rect 511398 280046 511494 280102
rect 510874 279978 511494 280046
rect 510874 279922 510970 279978
rect 511026 279922 511094 279978
rect 511150 279922 511218 279978
rect 511274 279922 511342 279978
rect 511398 279922 511494 279978
rect 510874 262350 511494 279922
rect 510874 262294 510970 262350
rect 511026 262294 511094 262350
rect 511150 262294 511218 262350
rect 511274 262294 511342 262350
rect 511398 262294 511494 262350
rect 510874 262226 511494 262294
rect 510874 262170 510970 262226
rect 511026 262170 511094 262226
rect 511150 262170 511218 262226
rect 511274 262170 511342 262226
rect 511398 262170 511494 262226
rect 510874 262102 511494 262170
rect 510874 262046 510970 262102
rect 511026 262046 511094 262102
rect 511150 262046 511218 262102
rect 511274 262046 511342 262102
rect 511398 262046 511494 262102
rect 510874 261978 511494 262046
rect 510874 261922 510970 261978
rect 511026 261922 511094 261978
rect 511150 261922 511218 261978
rect 511274 261922 511342 261978
rect 511398 261922 511494 261978
rect 510874 244350 511494 261922
rect 510874 244294 510970 244350
rect 511026 244294 511094 244350
rect 511150 244294 511218 244350
rect 511274 244294 511342 244350
rect 511398 244294 511494 244350
rect 510874 244226 511494 244294
rect 510874 244170 510970 244226
rect 511026 244170 511094 244226
rect 511150 244170 511218 244226
rect 511274 244170 511342 244226
rect 511398 244170 511494 244226
rect 510874 244102 511494 244170
rect 510874 244046 510970 244102
rect 511026 244046 511094 244102
rect 511150 244046 511218 244102
rect 511274 244046 511342 244102
rect 511398 244046 511494 244102
rect 510874 243978 511494 244046
rect 510874 243922 510970 243978
rect 511026 243922 511094 243978
rect 511150 243922 511218 243978
rect 511274 243922 511342 243978
rect 511398 243922 511494 243978
rect 510874 226350 511494 243922
rect 528874 598172 529494 598268
rect 528874 598116 528970 598172
rect 529026 598116 529094 598172
rect 529150 598116 529218 598172
rect 529274 598116 529342 598172
rect 529398 598116 529494 598172
rect 528874 598048 529494 598116
rect 528874 597992 528970 598048
rect 529026 597992 529094 598048
rect 529150 597992 529218 598048
rect 529274 597992 529342 598048
rect 529398 597992 529494 598048
rect 528874 597924 529494 597992
rect 528874 597868 528970 597924
rect 529026 597868 529094 597924
rect 529150 597868 529218 597924
rect 529274 597868 529342 597924
rect 529398 597868 529494 597924
rect 528874 597800 529494 597868
rect 528874 597744 528970 597800
rect 529026 597744 529094 597800
rect 529150 597744 529218 597800
rect 529274 597744 529342 597800
rect 529398 597744 529494 597800
rect 528874 586350 529494 597744
rect 543154 597212 543774 598268
rect 543154 597156 543250 597212
rect 543306 597156 543374 597212
rect 543430 597156 543498 597212
rect 543554 597156 543622 597212
rect 543678 597156 543774 597212
rect 543154 597088 543774 597156
rect 543154 597032 543250 597088
rect 543306 597032 543374 597088
rect 543430 597032 543498 597088
rect 543554 597032 543622 597088
rect 543678 597032 543774 597088
rect 543154 596964 543774 597032
rect 543154 596908 543250 596964
rect 543306 596908 543374 596964
rect 543430 596908 543498 596964
rect 543554 596908 543622 596964
rect 543678 596908 543774 596964
rect 543154 596840 543774 596908
rect 543154 596784 543250 596840
rect 543306 596784 543374 596840
rect 543430 596784 543498 596840
rect 543554 596784 543622 596840
rect 543678 596784 543774 596840
rect 540764 589764 540820 589774
rect 540764 589316 540820 589708
rect 540764 589250 540820 589260
rect 528874 586294 528970 586350
rect 529026 586294 529094 586350
rect 529150 586294 529218 586350
rect 529274 586294 529342 586350
rect 529398 586294 529494 586350
rect 528874 586226 529494 586294
rect 528874 586170 528970 586226
rect 529026 586170 529094 586226
rect 529150 586170 529218 586226
rect 529274 586170 529342 586226
rect 529398 586170 529494 586226
rect 528874 586102 529494 586170
rect 528874 586046 528970 586102
rect 529026 586046 529094 586102
rect 529150 586046 529218 586102
rect 529274 586046 529342 586102
rect 529398 586046 529494 586102
rect 528874 585978 529494 586046
rect 528874 585922 528970 585978
rect 529026 585922 529094 585978
rect 529150 585922 529218 585978
rect 529274 585922 529342 585978
rect 529398 585922 529494 585978
rect 528874 568350 529494 585922
rect 528874 568294 528970 568350
rect 529026 568294 529094 568350
rect 529150 568294 529218 568350
rect 529274 568294 529342 568350
rect 529398 568294 529494 568350
rect 528874 568226 529494 568294
rect 528874 568170 528970 568226
rect 529026 568170 529094 568226
rect 529150 568170 529218 568226
rect 529274 568170 529342 568226
rect 529398 568170 529494 568226
rect 528874 568102 529494 568170
rect 528874 568046 528970 568102
rect 529026 568046 529094 568102
rect 529150 568046 529218 568102
rect 529274 568046 529342 568102
rect 529398 568046 529494 568102
rect 528874 567978 529494 568046
rect 528874 567922 528970 567978
rect 529026 567922 529094 567978
rect 529150 567922 529218 567978
rect 529274 567922 529342 567978
rect 529398 567922 529494 567978
rect 528874 550350 529494 567922
rect 528874 550294 528970 550350
rect 529026 550294 529094 550350
rect 529150 550294 529218 550350
rect 529274 550294 529342 550350
rect 529398 550294 529494 550350
rect 528874 550226 529494 550294
rect 528874 550170 528970 550226
rect 529026 550170 529094 550226
rect 529150 550170 529218 550226
rect 529274 550170 529342 550226
rect 529398 550170 529494 550226
rect 528874 550102 529494 550170
rect 528874 550046 528970 550102
rect 529026 550046 529094 550102
rect 529150 550046 529218 550102
rect 529274 550046 529342 550102
rect 529398 550046 529494 550102
rect 528874 549978 529494 550046
rect 528874 549922 528970 549978
rect 529026 549922 529094 549978
rect 529150 549922 529218 549978
rect 529274 549922 529342 549978
rect 529398 549922 529494 549978
rect 528874 532350 529494 549922
rect 528874 532294 528970 532350
rect 529026 532294 529094 532350
rect 529150 532294 529218 532350
rect 529274 532294 529342 532350
rect 529398 532294 529494 532350
rect 528874 532226 529494 532294
rect 528874 532170 528970 532226
rect 529026 532170 529094 532226
rect 529150 532170 529218 532226
rect 529274 532170 529342 532226
rect 529398 532170 529494 532226
rect 528874 532102 529494 532170
rect 528874 532046 528970 532102
rect 529026 532046 529094 532102
rect 529150 532046 529218 532102
rect 529274 532046 529342 532102
rect 529398 532046 529494 532102
rect 528874 531978 529494 532046
rect 528874 531922 528970 531978
rect 529026 531922 529094 531978
rect 529150 531922 529218 531978
rect 529274 531922 529342 531978
rect 529398 531922 529494 531978
rect 528874 514350 529494 531922
rect 528874 514294 528970 514350
rect 529026 514294 529094 514350
rect 529150 514294 529218 514350
rect 529274 514294 529342 514350
rect 529398 514294 529494 514350
rect 528874 514226 529494 514294
rect 528874 514170 528970 514226
rect 529026 514170 529094 514226
rect 529150 514170 529218 514226
rect 529274 514170 529342 514226
rect 529398 514170 529494 514226
rect 528874 514102 529494 514170
rect 528874 514046 528970 514102
rect 529026 514046 529094 514102
rect 529150 514046 529218 514102
rect 529274 514046 529342 514102
rect 529398 514046 529494 514102
rect 528874 513978 529494 514046
rect 528874 513922 528970 513978
rect 529026 513922 529094 513978
rect 529150 513922 529218 513978
rect 529274 513922 529342 513978
rect 529398 513922 529494 513978
rect 528874 496350 529494 513922
rect 528874 496294 528970 496350
rect 529026 496294 529094 496350
rect 529150 496294 529218 496350
rect 529274 496294 529342 496350
rect 529398 496294 529494 496350
rect 528874 496226 529494 496294
rect 528874 496170 528970 496226
rect 529026 496170 529094 496226
rect 529150 496170 529218 496226
rect 529274 496170 529342 496226
rect 529398 496170 529494 496226
rect 528874 496102 529494 496170
rect 528874 496046 528970 496102
rect 529026 496046 529094 496102
rect 529150 496046 529218 496102
rect 529274 496046 529342 496102
rect 529398 496046 529494 496102
rect 528874 495978 529494 496046
rect 528874 495922 528970 495978
rect 529026 495922 529094 495978
rect 529150 495922 529218 495978
rect 529274 495922 529342 495978
rect 529398 495922 529494 495978
rect 528874 478350 529494 495922
rect 528874 478294 528970 478350
rect 529026 478294 529094 478350
rect 529150 478294 529218 478350
rect 529274 478294 529342 478350
rect 529398 478294 529494 478350
rect 528874 478226 529494 478294
rect 528874 478170 528970 478226
rect 529026 478170 529094 478226
rect 529150 478170 529218 478226
rect 529274 478170 529342 478226
rect 529398 478170 529494 478226
rect 528874 478102 529494 478170
rect 528874 478046 528970 478102
rect 529026 478046 529094 478102
rect 529150 478046 529218 478102
rect 529274 478046 529342 478102
rect 529398 478046 529494 478102
rect 528874 477978 529494 478046
rect 528874 477922 528970 477978
rect 529026 477922 529094 477978
rect 529150 477922 529218 477978
rect 529274 477922 529342 477978
rect 529398 477922 529494 477978
rect 528874 460350 529494 477922
rect 528874 460294 528970 460350
rect 529026 460294 529094 460350
rect 529150 460294 529218 460350
rect 529274 460294 529342 460350
rect 529398 460294 529494 460350
rect 528874 460226 529494 460294
rect 528874 460170 528970 460226
rect 529026 460170 529094 460226
rect 529150 460170 529218 460226
rect 529274 460170 529342 460226
rect 529398 460170 529494 460226
rect 528874 460102 529494 460170
rect 528874 460046 528970 460102
rect 529026 460046 529094 460102
rect 529150 460046 529218 460102
rect 529274 460046 529342 460102
rect 529398 460046 529494 460102
rect 528874 459978 529494 460046
rect 528874 459922 528970 459978
rect 529026 459922 529094 459978
rect 529150 459922 529218 459978
rect 529274 459922 529342 459978
rect 529398 459922 529494 459978
rect 528874 442350 529494 459922
rect 528874 442294 528970 442350
rect 529026 442294 529094 442350
rect 529150 442294 529218 442350
rect 529274 442294 529342 442350
rect 529398 442294 529494 442350
rect 528874 442226 529494 442294
rect 528874 442170 528970 442226
rect 529026 442170 529094 442226
rect 529150 442170 529218 442226
rect 529274 442170 529342 442226
rect 529398 442170 529494 442226
rect 528874 442102 529494 442170
rect 528874 442046 528970 442102
rect 529026 442046 529094 442102
rect 529150 442046 529218 442102
rect 529274 442046 529342 442102
rect 529398 442046 529494 442102
rect 528874 441978 529494 442046
rect 528874 441922 528970 441978
rect 529026 441922 529094 441978
rect 529150 441922 529218 441978
rect 529274 441922 529342 441978
rect 529398 441922 529494 441978
rect 528874 424350 529494 441922
rect 528874 424294 528970 424350
rect 529026 424294 529094 424350
rect 529150 424294 529218 424350
rect 529274 424294 529342 424350
rect 529398 424294 529494 424350
rect 528874 424226 529494 424294
rect 528874 424170 528970 424226
rect 529026 424170 529094 424226
rect 529150 424170 529218 424226
rect 529274 424170 529342 424226
rect 529398 424170 529494 424226
rect 528874 424102 529494 424170
rect 528874 424046 528970 424102
rect 529026 424046 529094 424102
rect 529150 424046 529218 424102
rect 529274 424046 529342 424102
rect 529398 424046 529494 424102
rect 528874 423978 529494 424046
rect 528874 423922 528970 423978
rect 529026 423922 529094 423978
rect 529150 423922 529218 423978
rect 529274 423922 529342 423978
rect 529398 423922 529494 423978
rect 528874 406350 529494 423922
rect 528874 406294 528970 406350
rect 529026 406294 529094 406350
rect 529150 406294 529218 406350
rect 529274 406294 529342 406350
rect 529398 406294 529494 406350
rect 528874 406226 529494 406294
rect 528874 406170 528970 406226
rect 529026 406170 529094 406226
rect 529150 406170 529218 406226
rect 529274 406170 529342 406226
rect 529398 406170 529494 406226
rect 528874 406102 529494 406170
rect 528874 406046 528970 406102
rect 529026 406046 529094 406102
rect 529150 406046 529218 406102
rect 529274 406046 529342 406102
rect 529398 406046 529494 406102
rect 528874 405978 529494 406046
rect 528874 405922 528970 405978
rect 529026 405922 529094 405978
rect 529150 405922 529218 405978
rect 529274 405922 529342 405978
rect 529398 405922 529494 405978
rect 528874 388350 529494 405922
rect 528874 388294 528970 388350
rect 529026 388294 529094 388350
rect 529150 388294 529218 388350
rect 529274 388294 529342 388350
rect 529398 388294 529494 388350
rect 528874 388226 529494 388294
rect 528874 388170 528970 388226
rect 529026 388170 529094 388226
rect 529150 388170 529218 388226
rect 529274 388170 529342 388226
rect 529398 388170 529494 388226
rect 528874 388102 529494 388170
rect 528874 388046 528970 388102
rect 529026 388046 529094 388102
rect 529150 388046 529218 388102
rect 529274 388046 529342 388102
rect 529398 388046 529494 388102
rect 528874 387978 529494 388046
rect 528874 387922 528970 387978
rect 529026 387922 529094 387978
rect 529150 387922 529218 387978
rect 529274 387922 529342 387978
rect 529398 387922 529494 387978
rect 528874 370350 529494 387922
rect 528874 370294 528970 370350
rect 529026 370294 529094 370350
rect 529150 370294 529218 370350
rect 529274 370294 529342 370350
rect 529398 370294 529494 370350
rect 528874 370226 529494 370294
rect 528874 370170 528970 370226
rect 529026 370170 529094 370226
rect 529150 370170 529218 370226
rect 529274 370170 529342 370226
rect 529398 370170 529494 370226
rect 528874 370102 529494 370170
rect 528874 370046 528970 370102
rect 529026 370046 529094 370102
rect 529150 370046 529218 370102
rect 529274 370046 529342 370102
rect 529398 370046 529494 370102
rect 528874 369978 529494 370046
rect 528874 369922 528970 369978
rect 529026 369922 529094 369978
rect 529150 369922 529218 369978
rect 529274 369922 529342 369978
rect 529398 369922 529494 369978
rect 528874 352350 529494 369922
rect 528874 352294 528970 352350
rect 529026 352294 529094 352350
rect 529150 352294 529218 352350
rect 529274 352294 529342 352350
rect 529398 352294 529494 352350
rect 528874 352226 529494 352294
rect 528874 352170 528970 352226
rect 529026 352170 529094 352226
rect 529150 352170 529218 352226
rect 529274 352170 529342 352226
rect 529398 352170 529494 352226
rect 528874 352102 529494 352170
rect 528874 352046 528970 352102
rect 529026 352046 529094 352102
rect 529150 352046 529218 352102
rect 529274 352046 529342 352102
rect 529398 352046 529494 352102
rect 528874 351978 529494 352046
rect 528874 351922 528970 351978
rect 529026 351922 529094 351978
rect 529150 351922 529218 351978
rect 529274 351922 529342 351978
rect 529398 351922 529494 351978
rect 528874 334350 529494 351922
rect 528874 334294 528970 334350
rect 529026 334294 529094 334350
rect 529150 334294 529218 334350
rect 529274 334294 529342 334350
rect 529398 334294 529494 334350
rect 528874 334226 529494 334294
rect 528874 334170 528970 334226
rect 529026 334170 529094 334226
rect 529150 334170 529218 334226
rect 529274 334170 529342 334226
rect 529398 334170 529494 334226
rect 528874 334102 529494 334170
rect 528874 334046 528970 334102
rect 529026 334046 529094 334102
rect 529150 334046 529218 334102
rect 529274 334046 529342 334102
rect 529398 334046 529494 334102
rect 528874 333978 529494 334046
rect 528874 333922 528970 333978
rect 529026 333922 529094 333978
rect 529150 333922 529218 333978
rect 529274 333922 529342 333978
rect 529398 333922 529494 333978
rect 528874 316350 529494 333922
rect 528874 316294 528970 316350
rect 529026 316294 529094 316350
rect 529150 316294 529218 316350
rect 529274 316294 529342 316350
rect 529398 316294 529494 316350
rect 528874 316226 529494 316294
rect 528874 316170 528970 316226
rect 529026 316170 529094 316226
rect 529150 316170 529218 316226
rect 529274 316170 529342 316226
rect 529398 316170 529494 316226
rect 528874 316102 529494 316170
rect 528874 316046 528970 316102
rect 529026 316046 529094 316102
rect 529150 316046 529218 316102
rect 529274 316046 529342 316102
rect 529398 316046 529494 316102
rect 528874 315978 529494 316046
rect 528874 315922 528970 315978
rect 529026 315922 529094 315978
rect 529150 315922 529218 315978
rect 529274 315922 529342 315978
rect 529398 315922 529494 315978
rect 528874 298350 529494 315922
rect 528874 298294 528970 298350
rect 529026 298294 529094 298350
rect 529150 298294 529218 298350
rect 529274 298294 529342 298350
rect 529398 298294 529494 298350
rect 528874 298226 529494 298294
rect 528874 298170 528970 298226
rect 529026 298170 529094 298226
rect 529150 298170 529218 298226
rect 529274 298170 529342 298226
rect 529398 298170 529494 298226
rect 528874 298102 529494 298170
rect 528874 298046 528970 298102
rect 529026 298046 529094 298102
rect 529150 298046 529218 298102
rect 529274 298046 529342 298102
rect 529398 298046 529494 298102
rect 528874 297978 529494 298046
rect 528874 297922 528970 297978
rect 529026 297922 529094 297978
rect 529150 297922 529218 297978
rect 529274 297922 529342 297978
rect 529398 297922 529494 297978
rect 528874 280350 529494 297922
rect 528874 280294 528970 280350
rect 529026 280294 529094 280350
rect 529150 280294 529218 280350
rect 529274 280294 529342 280350
rect 529398 280294 529494 280350
rect 528874 280226 529494 280294
rect 528874 280170 528970 280226
rect 529026 280170 529094 280226
rect 529150 280170 529218 280226
rect 529274 280170 529342 280226
rect 529398 280170 529494 280226
rect 528874 280102 529494 280170
rect 528874 280046 528970 280102
rect 529026 280046 529094 280102
rect 529150 280046 529218 280102
rect 529274 280046 529342 280102
rect 529398 280046 529494 280102
rect 528874 279978 529494 280046
rect 528874 279922 528970 279978
rect 529026 279922 529094 279978
rect 529150 279922 529218 279978
rect 529274 279922 529342 279978
rect 529398 279922 529494 279978
rect 528874 262350 529494 279922
rect 528874 262294 528970 262350
rect 529026 262294 529094 262350
rect 529150 262294 529218 262350
rect 529274 262294 529342 262350
rect 529398 262294 529494 262350
rect 528874 262226 529494 262294
rect 528874 262170 528970 262226
rect 529026 262170 529094 262226
rect 529150 262170 529218 262226
rect 529274 262170 529342 262226
rect 529398 262170 529494 262226
rect 528874 262102 529494 262170
rect 528874 262046 528970 262102
rect 529026 262046 529094 262102
rect 529150 262046 529218 262102
rect 529274 262046 529342 262102
rect 529398 262046 529494 262102
rect 528874 261978 529494 262046
rect 528874 261922 528970 261978
rect 529026 261922 529094 261978
rect 529150 261922 529218 261978
rect 529274 261922 529342 261978
rect 529398 261922 529494 261978
rect 528874 244350 529494 261922
rect 528874 244294 528970 244350
rect 529026 244294 529094 244350
rect 529150 244294 529218 244350
rect 529274 244294 529342 244350
rect 529398 244294 529494 244350
rect 528874 244226 529494 244294
rect 528874 244170 528970 244226
rect 529026 244170 529094 244226
rect 529150 244170 529218 244226
rect 529274 244170 529342 244226
rect 529398 244170 529494 244226
rect 528874 244102 529494 244170
rect 528874 244046 528970 244102
rect 529026 244046 529094 244102
rect 529150 244046 529218 244102
rect 529274 244046 529342 244102
rect 529398 244046 529494 244102
rect 528874 243978 529494 244046
rect 528874 243922 528970 243978
rect 529026 243922 529094 243978
rect 529150 243922 529218 243978
rect 529274 243922 529342 243978
rect 529398 243922 529494 243978
rect 510874 226294 510970 226350
rect 511026 226294 511094 226350
rect 511150 226294 511218 226350
rect 511274 226294 511342 226350
rect 511398 226294 511494 226350
rect 510874 226226 511494 226294
rect 510874 226170 510970 226226
rect 511026 226170 511094 226226
rect 511150 226170 511218 226226
rect 511274 226170 511342 226226
rect 511398 226170 511494 226226
rect 510874 226102 511494 226170
rect 510874 226046 510970 226102
rect 511026 226046 511094 226102
rect 511150 226046 511218 226102
rect 511274 226046 511342 226102
rect 511398 226046 511494 226102
rect 510874 225978 511494 226046
rect 510874 225922 510970 225978
rect 511026 225922 511094 225978
rect 511150 225922 511218 225978
rect 511274 225922 511342 225978
rect 511398 225922 511494 225978
rect 510874 217934 511494 225922
rect 525154 238350 525774 242964
rect 525154 238294 525250 238350
rect 525306 238294 525374 238350
rect 525430 238294 525498 238350
rect 525554 238294 525622 238350
rect 525678 238294 525774 238350
rect 525154 238226 525774 238294
rect 525154 238170 525250 238226
rect 525306 238170 525374 238226
rect 525430 238170 525498 238226
rect 525554 238170 525622 238226
rect 525678 238170 525774 238226
rect 525154 238102 525774 238170
rect 525154 238046 525250 238102
rect 525306 238046 525374 238102
rect 525430 238046 525498 238102
rect 525554 238046 525622 238102
rect 525678 238046 525774 238102
rect 525154 237978 525774 238046
rect 525154 237922 525250 237978
rect 525306 237922 525374 237978
rect 525430 237922 525498 237978
rect 525554 237922 525622 237978
rect 525678 237922 525774 237978
rect 525154 220350 525774 237922
rect 525154 220294 525250 220350
rect 525306 220294 525374 220350
rect 525430 220294 525498 220350
rect 525554 220294 525622 220350
rect 525678 220294 525774 220350
rect 525154 220226 525774 220294
rect 525154 220170 525250 220226
rect 525306 220170 525374 220226
rect 525430 220170 525498 220226
rect 525554 220170 525622 220226
rect 525678 220170 525774 220226
rect 525154 220102 525774 220170
rect 525154 220046 525250 220102
rect 525306 220046 525374 220102
rect 525430 220046 525498 220102
rect 525554 220046 525622 220102
rect 525678 220046 525774 220102
rect 525154 219978 525774 220046
rect 525154 219922 525250 219978
rect 525306 219922 525374 219978
rect 525430 219922 525498 219978
rect 525554 219922 525622 219978
rect 525678 219922 525774 219978
rect 525154 218572 525774 219922
rect 528874 226350 529494 243922
rect 528874 226294 528970 226350
rect 529026 226294 529094 226350
rect 529150 226294 529218 226350
rect 529274 226294 529342 226350
rect 529398 226294 529494 226350
rect 528874 226226 529494 226294
rect 528874 226170 528970 226226
rect 529026 226170 529094 226226
rect 529150 226170 529218 226226
rect 529274 226170 529342 226226
rect 529398 226170 529494 226226
rect 528874 226102 529494 226170
rect 528874 226046 528970 226102
rect 529026 226046 529094 226102
rect 529150 226046 529218 226102
rect 529274 226046 529342 226102
rect 529398 226046 529494 226102
rect 528874 225978 529494 226046
rect 528874 225922 528970 225978
rect 529026 225922 529094 225978
rect 529150 225922 529218 225978
rect 529274 225922 529342 225978
rect 529398 225922 529494 225978
rect 528874 217934 529494 225922
rect 543154 580350 543774 596784
rect 543154 580294 543250 580350
rect 543306 580294 543374 580350
rect 543430 580294 543498 580350
rect 543554 580294 543622 580350
rect 543678 580294 543774 580350
rect 543154 580226 543774 580294
rect 543154 580170 543250 580226
rect 543306 580170 543374 580226
rect 543430 580170 543498 580226
rect 543554 580170 543622 580226
rect 543678 580170 543774 580226
rect 543154 580102 543774 580170
rect 543154 580046 543250 580102
rect 543306 580046 543374 580102
rect 543430 580046 543498 580102
rect 543554 580046 543622 580102
rect 543678 580046 543774 580102
rect 543154 579978 543774 580046
rect 543154 579922 543250 579978
rect 543306 579922 543374 579978
rect 543430 579922 543498 579978
rect 543554 579922 543622 579978
rect 543678 579922 543774 579978
rect 543154 562350 543774 579922
rect 543154 562294 543250 562350
rect 543306 562294 543374 562350
rect 543430 562294 543498 562350
rect 543554 562294 543622 562350
rect 543678 562294 543774 562350
rect 543154 562226 543774 562294
rect 543154 562170 543250 562226
rect 543306 562170 543374 562226
rect 543430 562170 543498 562226
rect 543554 562170 543622 562226
rect 543678 562170 543774 562226
rect 543154 562102 543774 562170
rect 543154 562046 543250 562102
rect 543306 562046 543374 562102
rect 543430 562046 543498 562102
rect 543554 562046 543622 562102
rect 543678 562046 543774 562102
rect 543154 561978 543774 562046
rect 543154 561922 543250 561978
rect 543306 561922 543374 561978
rect 543430 561922 543498 561978
rect 543554 561922 543622 561978
rect 543678 561922 543774 561978
rect 543154 544350 543774 561922
rect 543154 544294 543250 544350
rect 543306 544294 543374 544350
rect 543430 544294 543498 544350
rect 543554 544294 543622 544350
rect 543678 544294 543774 544350
rect 543154 544226 543774 544294
rect 543154 544170 543250 544226
rect 543306 544170 543374 544226
rect 543430 544170 543498 544226
rect 543554 544170 543622 544226
rect 543678 544170 543774 544226
rect 543154 544102 543774 544170
rect 543154 544046 543250 544102
rect 543306 544046 543374 544102
rect 543430 544046 543498 544102
rect 543554 544046 543622 544102
rect 543678 544046 543774 544102
rect 543154 543978 543774 544046
rect 543154 543922 543250 543978
rect 543306 543922 543374 543978
rect 543430 543922 543498 543978
rect 543554 543922 543622 543978
rect 543678 543922 543774 543978
rect 543154 526350 543774 543922
rect 543154 526294 543250 526350
rect 543306 526294 543374 526350
rect 543430 526294 543498 526350
rect 543554 526294 543622 526350
rect 543678 526294 543774 526350
rect 543154 526226 543774 526294
rect 543154 526170 543250 526226
rect 543306 526170 543374 526226
rect 543430 526170 543498 526226
rect 543554 526170 543622 526226
rect 543678 526170 543774 526226
rect 543154 526102 543774 526170
rect 543154 526046 543250 526102
rect 543306 526046 543374 526102
rect 543430 526046 543498 526102
rect 543554 526046 543622 526102
rect 543678 526046 543774 526102
rect 543154 525978 543774 526046
rect 543154 525922 543250 525978
rect 543306 525922 543374 525978
rect 543430 525922 543498 525978
rect 543554 525922 543622 525978
rect 543678 525922 543774 525978
rect 543154 508350 543774 525922
rect 543154 508294 543250 508350
rect 543306 508294 543374 508350
rect 543430 508294 543498 508350
rect 543554 508294 543622 508350
rect 543678 508294 543774 508350
rect 543154 508226 543774 508294
rect 543154 508170 543250 508226
rect 543306 508170 543374 508226
rect 543430 508170 543498 508226
rect 543554 508170 543622 508226
rect 543678 508170 543774 508226
rect 543154 508102 543774 508170
rect 543154 508046 543250 508102
rect 543306 508046 543374 508102
rect 543430 508046 543498 508102
rect 543554 508046 543622 508102
rect 543678 508046 543774 508102
rect 543154 507978 543774 508046
rect 543154 507922 543250 507978
rect 543306 507922 543374 507978
rect 543430 507922 543498 507978
rect 543554 507922 543622 507978
rect 543678 507922 543774 507978
rect 543154 490350 543774 507922
rect 543154 490294 543250 490350
rect 543306 490294 543374 490350
rect 543430 490294 543498 490350
rect 543554 490294 543622 490350
rect 543678 490294 543774 490350
rect 543154 490226 543774 490294
rect 543154 490170 543250 490226
rect 543306 490170 543374 490226
rect 543430 490170 543498 490226
rect 543554 490170 543622 490226
rect 543678 490170 543774 490226
rect 543154 490102 543774 490170
rect 543154 490046 543250 490102
rect 543306 490046 543374 490102
rect 543430 490046 543498 490102
rect 543554 490046 543622 490102
rect 543678 490046 543774 490102
rect 543154 489978 543774 490046
rect 543154 489922 543250 489978
rect 543306 489922 543374 489978
rect 543430 489922 543498 489978
rect 543554 489922 543622 489978
rect 543678 489922 543774 489978
rect 543154 472350 543774 489922
rect 543154 472294 543250 472350
rect 543306 472294 543374 472350
rect 543430 472294 543498 472350
rect 543554 472294 543622 472350
rect 543678 472294 543774 472350
rect 543154 472226 543774 472294
rect 543154 472170 543250 472226
rect 543306 472170 543374 472226
rect 543430 472170 543498 472226
rect 543554 472170 543622 472226
rect 543678 472170 543774 472226
rect 543154 472102 543774 472170
rect 543154 472046 543250 472102
rect 543306 472046 543374 472102
rect 543430 472046 543498 472102
rect 543554 472046 543622 472102
rect 543678 472046 543774 472102
rect 543154 471978 543774 472046
rect 543154 471922 543250 471978
rect 543306 471922 543374 471978
rect 543430 471922 543498 471978
rect 543554 471922 543622 471978
rect 543678 471922 543774 471978
rect 543154 454350 543774 471922
rect 543154 454294 543250 454350
rect 543306 454294 543374 454350
rect 543430 454294 543498 454350
rect 543554 454294 543622 454350
rect 543678 454294 543774 454350
rect 543154 454226 543774 454294
rect 543154 454170 543250 454226
rect 543306 454170 543374 454226
rect 543430 454170 543498 454226
rect 543554 454170 543622 454226
rect 543678 454170 543774 454226
rect 543154 454102 543774 454170
rect 543154 454046 543250 454102
rect 543306 454046 543374 454102
rect 543430 454046 543498 454102
rect 543554 454046 543622 454102
rect 543678 454046 543774 454102
rect 543154 453978 543774 454046
rect 543154 453922 543250 453978
rect 543306 453922 543374 453978
rect 543430 453922 543498 453978
rect 543554 453922 543622 453978
rect 543678 453922 543774 453978
rect 543154 436350 543774 453922
rect 543154 436294 543250 436350
rect 543306 436294 543374 436350
rect 543430 436294 543498 436350
rect 543554 436294 543622 436350
rect 543678 436294 543774 436350
rect 543154 436226 543774 436294
rect 543154 436170 543250 436226
rect 543306 436170 543374 436226
rect 543430 436170 543498 436226
rect 543554 436170 543622 436226
rect 543678 436170 543774 436226
rect 543154 436102 543774 436170
rect 543154 436046 543250 436102
rect 543306 436046 543374 436102
rect 543430 436046 543498 436102
rect 543554 436046 543622 436102
rect 543678 436046 543774 436102
rect 543154 435978 543774 436046
rect 543154 435922 543250 435978
rect 543306 435922 543374 435978
rect 543430 435922 543498 435978
rect 543554 435922 543622 435978
rect 543678 435922 543774 435978
rect 543154 418350 543774 435922
rect 543154 418294 543250 418350
rect 543306 418294 543374 418350
rect 543430 418294 543498 418350
rect 543554 418294 543622 418350
rect 543678 418294 543774 418350
rect 543154 418226 543774 418294
rect 543154 418170 543250 418226
rect 543306 418170 543374 418226
rect 543430 418170 543498 418226
rect 543554 418170 543622 418226
rect 543678 418170 543774 418226
rect 543154 418102 543774 418170
rect 543154 418046 543250 418102
rect 543306 418046 543374 418102
rect 543430 418046 543498 418102
rect 543554 418046 543622 418102
rect 543678 418046 543774 418102
rect 543154 417978 543774 418046
rect 543154 417922 543250 417978
rect 543306 417922 543374 417978
rect 543430 417922 543498 417978
rect 543554 417922 543622 417978
rect 543678 417922 543774 417978
rect 543154 400350 543774 417922
rect 543154 400294 543250 400350
rect 543306 400294 543374 400350
rect 543430 400294 543498 400350
rect 543554 400294 543622 400350
rect 543678 400294 543774 400350
rect 543154 400226 543774 400294
rect 543154 400170 543250 400226
rect 543306 400170 543374 400226
rect 543430 400170 543498 400226
rect 543554 400170 543622 400226
rect 543678 400170 543774 400226
rect 543154 400102 543774 400170
rect 543154 400046 543250 400102
rect 543306 400046 543374 400102
rect 543430 400046 543498 400102
rect 543554 400046 543622 400102
rect 543678 400046 543774 400102
rect 543154 399978 543774 400046
rect 543154 399922 543250 399978
rect 543306 399922 543374 399978
rect 543430 399922 543498 399978
rect 543554 399922 543622 399978
rect 543678 399922 543774 399978
rect 543154 382350 543774 399922
rect 543154 382294 543250 382350
rect 543306 382294 543374 382350
rect 543430 382294 543498 382350
rect 543554 382294 543622 382350
rect 543678 382294 543774 382350
rect 543154 382226 543774 382294
rect 543154 382170 543250 382226
rect 543306 382170 543374 382226
rect 543430 382170 543498 382226
rect 543554 382170 543622 382226
rect 543678 382170 543774 382226
rect 543154 382102 543774 382170
rect 543154 382046 543250 382102
rect 543306 382046 543374 382102
rect 543430 382046 543498 382102
rect 543554 382046 543622 382102
rect 543678 382046 543774 382102
rect 543154 381978 543774 382046
rect 543154 381922 543250 381978
rect 543306 381922 543374 381978
rect 543430 381922 543498 381978
rect 543554 381922 543622 381978
rect 543678 381922 543774 381978
rect 543154 364350 543774 381922
rect 543154 364294 543250 364350
rect 543306 364294 543374 364350
rect 543430 364294 543498 364350
rect 543554 364294 543622 364350
rect 543678 364294 543774 364350
rect 543154 364226 543774 364294
rect 543154 364170 543250 364226
rect 543306 364170 543374 364226
rect 543430 364170 543498 364226
rect 543554 364170 543622 364226
rect 543678 364170 543774 364226
rect 543154 364102 543774 364170
rect 543154 364046 543250 364102
rect 543306 364046 543374 364102
rect 543430 364046 543498 364102
rect 543554 364046 543622 364102
rect 543678 364046 543774 364102
rect 543154 363978 543774 364046
rect 543154 363922 543250 363978
rect 543306 363922 543374 363978
rect 543430 363922 543498 363978
rect 543554 363922 543622 363978
rect 543678 363922 543774 363978
rect 543154 346350 543774 363922
rect 543154 346294 543250 346350
rect 543306 346294 543374 346350
rect 543430 346294 543498 346350
rect 543554 346294 543622 346350
rect 543678 346294 543774 346350
rect 543154 346226 543774 346294
rect 543154 346170 543250 346226
rect 543306 346170 543374 346226
rect 543430 346170 543498 346226
rect 543554 346170 543622 346226
rect 543678 346170 543774 346226
rect 543154 346102 543774 346170
rect 543154 346046 543250 346102
rect 543306 346046 543374 346102
rect 543430 346046 543498 346102
rect 543554 346046 543622 346102
rect 543678 346046 543774 346102
rect 543154 345978 543774 346046
rect 543154 345922 543250 345978
rect 543306 345922 543374 345978
rect 543430 345922 543498 345978
rect 543554 345922 543622 345978
rect 543678 345922 543774 345978
rect 543154 328350 543774 345922
rect 543154 328294 543250 328350
rect 543306 328294 543374 328350
rect 543430 328294 543498 328350
rect 543554 328294 543622 328350
rect 543678 328294 543774 328350
rect 543154 328226 543774 328294
rect 543154 328170 543250 328226
rect 543306 328170 543374 328226
rect 543430 328170 543498 328226
rect 543554 328170 543622 328226
rect 543678 328170 543774 328226
rect 543154 328102 543774 328170
rect 543154 328046 543250 328102
rect 543306 328046 543374 328102
rect 543430 328046 543498 328102
rect 543554 328046 543622 328102
rect 543678 328046 543774 328102
rect 543154 327978 543774 328046
rect 543154 327922 543250 327978
rect 543306 327922 543374 327978
rect 543430 327922 543498 327978
rect 543554 327922 543622 327978
rect 543678 327922 543774 327978
rect 543154 310350 543774 327922
rect 543154 310294 543250 310350
rect 543306 310294 543374 310350
rect 543430 310294 543498 310350
rect 543554 310294 543622 310350
rect 543678 310294 543774 310350
rect 543154 310226 543774 310294
rect 543154 310170 543250 310226
rect 543306 310170 543374 310226
rect 543430 310170 543498 310226
rect 543554 310170 543622 310226
rect 543678 310170 543774 310226
rect 543154 310102 543774 310170
rect 543154 310046 543250 310102
rect 543306 310046 543374 310102
rect 543430 310046 543498 310102
rect 543554 310046 543622 310102
rect 543678 310046 543774 310102
rect 543154 309978 543774 310046
rect 543154 309922 543250 309978
rect 543306 309922 543374 309978
rect 543430 309922 543498 309978
rect 543554 309922 543622 309978
rect 543678 309922 543774 309978
rect 543154 292350 543774 309922
rect 543154 292294 543250 292350
rect 543306 292294 543374 292350
rect 543430 292294 543498 292350
rect 543554 292294 543622 292350
rect 543678 292294 543774 292350
rect 543154 292226 543774 292294
rect 543154 292170 543250 292226
rect 543306 292170 543374 292226
rect 543430 292170 543498 292226
rect 543554 292170 543622 292226
rect 543678 292170 543774 292226
rect 543154 292102 543774 292170
rect 543154 292046 543250 292102
rect 543306 292046 543374 292102
rect 543430 292046 543498 292102
rect 543554 292046 543622 292102
rect 543678 292046 543774 292102
rect 543154 291978 543774 292046
rect 543154 291922 543250 291978
rect 543306 291922 543374 291978
rect 543430 291922 543498 291978
rect 543554 291922 543622 291978
rect 543678 291922 543774 291978
rect 543154 274350 543774 291922
rect 543154 274294 543250 274350
rect 543306 274294 543374 274350
rect 543430 274294 543498 274350
rect 543554 274294 543622 274350
rect 543678 274294 543774 274350
rect 543154 274226 543774 274294
rect 543154 274170 543250 274226
rect 543306 274170 543374 274226
rect 543430 274170 543498 274226
rect 543554 274170 543622 274226
rect 543678 274170 543774 274226
rect 543154 274102 543774 274170
rect 543154 274046 543250 274102
rect 543306 274046 543374 274102
rect 543430 274046 543498 274102
rect 543554 274046 543622 274102
rect 543678 274046 543774 274102
rect 543154 273978 543774 274046
rect 543154 273922 543250 273978
rect 543306 273922 543374 273978
rect 543430 273922 543498 273978
rect 543554 273922 543622 273978
rect 543678 273922 543774 273978
rect 543154 256350 543774 273922
rect 543154 256294 543250 256350
rect 543306 256294 543374 256350
rect 543430 256294 543498 256350
rect 543554 256294 543622 256350
rect 543678 256294 543774 256350
rect 543154 256226 543774 256294
rect 543154 256170 543250 256226
rect 543306 256170 543374 256226
rect 543430 256170 543498 256226
rect 543554 256170 543622 256226
rect 543678 256170 543774 256226
rect 543154 256102 543774 256170
rect 543154 256046 543250 256102
rect 543306 256046 543374 256102
rect 543430 256046 543498 256102
rect 543554 256046 543622 256102
rect 543678 256046 543774 256102
rect 543154 255978 543774 256046
rect 543154 255922 543250 255978
rect 543306 255922 543374 255978
rect 543430 255922 543498 255978
rect 543554 255922 543622 255978
rect 543678 255922 543774 255978
rect 543154 238350 543774 255922
rect 543154 238294 543250 238350
rect 543306 238294 543374 238350
rect 543430 238294 543498 238350
rect 543554 238294 543622 238350
rect 543678 238294 543774 238350
rect 543154 238226 543774 238294
rect 543154 238170 543250 238226
rect 543306 238170 543374 238226
rect 543430 238170 543498 238226
rect 543554 238170 543622 238226
rect 543678 238170 543774 238226
rect 543154 238102 543774 238170
rect 543154 238046 543250 238102
rect 543306 238046 543374 238102
rect 543430 238046 543498 238102
rect 543554 238046 543622 238102
rect 543678 238046 543774 238102
rect 543154 237978 543774 238046
rect 543154 237922 543250 237978
rect 543306 237922 543374 237978
rect 543430 237922 543498 237978
rect 543554 237922 543622 237978
rect 543678 237922 543774 237978
rect 543154 220350 543774 237922
rect 543154 220294 543250 220350
rect 543306 220294 543374 220350
rect 543430 220294 543498 220350
rect 543554 220294 543622 220350
rect 543678 220294 543774 220350
rect 543154 220226 543774 220294
rect 543154 220170 543250 220226
rect 543306 220170 543374 220226
rect 543430 220170 543498 220226
rect 543554 220170 543622 220226
rect 543678 220170 543774 220226
rect 543154 220102 543774 220170
rect 543154 220046 543250 220102
rect 543306 220046 543374 220102
rect 543430 220046 543498 220102
rect 543554 220046 543622 220102
rect 543678 220046 543774 220102
rect 543154 219978 543774 220046
rect 543154 219922 543250 219978
rect 543306 219922 543374 219978
rect 543430 219922 543498 219978
rect 543554 219922 543622 219978
rect 543678 219922 543774 219978
rect 543154 217934 543774 219922
rect 546874 598172 547494 598268
rect 546874 598116 546970 598172
rect 547026 598116 547094 598172
rect 547150 598116 547218 598172
rect 547274 598116 547342 598172
rect 547398 598116 547494 598172
rect 546874 598048 547494 598116
rect 546874 597992 546970 598048
rect 547026 597992 547094 598048
rect 547150 597992 547218 598048
rect 547274 597992 547342 598048
rect 547398 597992 547494 598048
rect 546874 597924 547494 597992
rect 546874 597868 546970 597924
rect 547026 597868 547094 597924
rect 547150 597868 547218 597924
rect 547274 597868 547342 597924
rect 547398 597868 547494 597924
rect 546874 597800 547494 597868
rect 546874 597744 546970 597800
rect 547026 597744 547094 597800
rect 547150 597744 547218 597800
rect 547274 597744 547342 597800
rect 547398 597744 547494 597800
rect 546874 586350 547494 597744
rect 546874 586294 546970 586350
rect 547026 586294 547094 586350
rect 547150 586294 547218 586350
rect 547274 586294 547342 586350
rect 547398 586294 547494 586350
rect 546874 586226 547494 586294
rect 546874 586170 546970 586226
rect 547026 586170 547094 586226
rect 547150 586170 547218 586226
rect 547274 586170 547342 586226
rect 547398 586170 547494 586226
rect 546874 586102 547494 586170
rect 546874 586046 546970 586102
rect 547026 586046 547094 586102
rect 547150 586046 547218 586102
rect 547274 586046 547342 586102
rect 547398 586046 547494 586102
rect 546874 585978 547494 586046
rect 546874 585922 546970 585978
rect 547026 585922 547094 585978
rect 547150 585922 547218 585978
rect 547274 585922 547342 585978
rect 547398 585922 547494 585978
rect 546874 568350 547494 585922
rect 546874 568294 546970 568350
rect 547026 568294 547094 568350
rect 547150 568294 547218 568350
rect 547274 568294 547342 568350
rect 547398 568294 547494 568350
rect 546874 568226 547494 568294
rect 546874 568170 546970 568226
rect 547026 568170 547094 568226
rect 547150 568170 547218 568226
rect 547274 568170 547342 568226
rect 547398 568170 547494 568226
rect 546874 568102 547494 568170
rect 546874 568046 546970 568102
rect 547026 568046 547094 568102
rect 547150 568046 547218 568102
rect 547274 568046 547342 568102
rect 547398 568046 547494 568102
rect 546874 567978 547494 568046
rect 546874 567922 546970 567978
rect 547026 567922 547094 567978
rect 547150 567922 547218 567978
rect 547274 567922 547342 567978
rect 547398 567922 547494 567978
rect 546874 550350 547494 567922
rect 546874 550294 546970 550350
rect 547026 550294 547094 550350
rect 547150 550294 547218 550350
rect 547274 550294 547342 550350
rect 547398 550294 547494 550350
rect 546874 550226 547494 550294
rect 546874 550170 546970 550226
rect 547026 550170 547094 550226
rect 547150 550170 547218 550226
rect 547274 550170 547342 550226
rect 547398 550170 547494 550226
rect 546874 550102 547494 550170
rect 546874 550046 546970 550102
rect 547026 550046 547094 550102
rect 547150 550046 547218 550102
rect 547274 550046 547342 550102
rect 547398 550046 547494 550102
rect 546874 549978 547494 550046
rect 546874 549922 546970 549978
rect 547026 549922 547094 549978
rect 547150 549922 547218 549978
rect 547274 549922 547342 549978
rect 547398 549922 547494 549978
rect 546874 532350 547494 549922
rect 546874 532294 546970 532350
rect 547026 532294 547094 532350
rect 547150 532294 547218 532350
rect 547274 532294 547342 532350
rect 547398 532294 547494 532350
rect 546874 532226 547494 532294
rect 546874 532170 546970 532226
rect 547026 532170 547094 532226
rect 547150 532170 547218 532226
rect 547274 532170 547342 532226
rect 547398 532170 547494 532226
rect 546874 532102 547494 532170
rect 546874 532046 546970 532102
rect 547026 532046 547094 532102
rect 547150 532046 547218 532102
rect 547274 532046 547342 532102
rect 547398 532046 547494 532102
rect 546874 531978 547494 532046
rect 546874 531922 546970 531978
rect 547026 531922 547094 531978
rect 547150 531922 547218 531978
rect 547274 531922 547342 531978
rect 547398 531922 547494 531978
rect 546874 514350 547494 531922
rect 546874 514294 546970 514350
rect 547026 514294 547094 514350
rect 547150 514294 547218 514350
rect 547274 514294 547342 514350
rect 547398 514294 547494 514350
rect 546874 514226 547494 514294
rect 546874 514170 546970 514226
rect 547026 514170 547094 514226
rect 547150 514170 547218 514226
rect 547274 514170 547342 514226
rect 547398 514170 547494 514226
rect 546874 514102 547494 514170
rect 546874 514046 546970 514102
rect 547026 514046 547094 514102
rect 547150 514046 547218 514102
rect 547274 514046 547342 514102
rect 547398 514046 547494 514102
rect 546874 513978 547494 514046
rect 546874 513922 546970 513978
rect 547026 513922 547094 513978
rect 547150 513922 547218 513978
rect 547274 513922 547342 513978
rect 547398 513922 547494 513978
rect 546874 496350 547494 513922
rect 546874 496294 546970 496350
rect 547026 496294 547094 496350
rect 547150 496294 547218 496350
rect 547274 496294 547342 496350
rect 547398 496294 547494 496350
rect 546874 496226 547494 496294
rect 546874 496170 546970 496226
rect 547026 496170 547094 496226
rect 547150 496170 547218 496226
rect 547274 496170 547342 496226
rect 547398 496170 547494 496226
rect 546874 496102 547494 496170
rect 546874 496046 546970 496102
rect 547026 496046 547094 496102
rect 547150 496046 547218 496102
rect 547274 496046 547342 496102
rect 547398 496046 547494 496102
rect 546874 495978 547494 496046
rect 546874 495922 546970 495978
rect 547026 495922 547094 495978
rect 547150 495922 547218 495978
rect 547274 495922 547342 495978
rect 547398 495922 547494 495978
rect 546874 478350 547494 495922
rect 561154 597212 561774 598268
rect 561154 597156 561250 597212
rect 561306 597156 561374 597212
rect 561430 597156 561498 597212
rect 561554 597156 561622 597212
rect 561678 597156 561774 597212
rect 561154 597088 561774 597156
rect 561154 597032 561250 597088
rect 561306 597032 561374 597088
rect 561430 597032 561498 597088
rect 561554 597032 561622 597088
rect 561678 597032 561774 597088
rect 561154 596964 561774 597032
rect 561154 596908 561250 596964
rect 561306 596908 561374 596964
rect 561430 596908 561498 596964
rect 561554 596908 561622 596964
rect 561678 596908 561774 596964
rect 561154 596840 561774 596908
rect 561154 596784 561250 596840
rect 561306 596784 561374 596840
rect 561430 596784 561498 596840
rect 561554 596784 561622 596840
rect 561678 596784 561774 596840
rect 561154 580350 561774 596784
rect 561154 580294 561250 580350
rect 561306 580294 561374 580350
rect 561430 580294 561498 580350
rect 561554 580294 561622 580350
rect 561678 580294 561774 580350
rect 561154 580226 561774 580294
rect 561154 580170 561250 580226
rect 561306 580170 561374 580226
rect 561430 580170 561498 580226
rect 561554 580170 561622 580226
rect 561678 580170 561774 580226
rect 561154 580102 561774 580170
rect 561154 580046 561250 580102
rect 561306 580046 561374 580102
rect 561430 580046 561498 580102
rect 561554 580046 561622 580102
rect 561678 580046 561774 580102
rect 561154 579978 561774 580046
rect 561154 579922 561250 579978
rect 561306 579922 561374 579978
rect 561430 579922 561498 579978
rect 561554 579922 561622 579978
rect 561678 579922 561774 579978
rect 561154 562350 561774 579922
rect 561154 562294 561250 562350
rect 561306 562294 561374 562350
rect 561430 562294 561498 562350
rect 561554 562294 561622 562350
rect 561678 562294 561774 562350
rect 561154 562226 561774 562294
rect 561154 562170 561250 562226
rect 561306 562170 561374 562226
rect 561430 562170 561498 562226
rect 561554 562170 561622 562226
rect 561678 562170 561774 562226
rect 561154 562102 561774 562170
rect 561154 562046 561250 562102
rect 561306 562046 561374 562102
rect 561430 562046 561498 562102
rect 561554 562046 561622 562102
rect 561678 562046 561774 562102
rect 561154 561978 561774 562046
rect 561154 561922 561250 561978
rect 561306 561922 561374 561978
rect 561430 561922 561498 561978
rect 561554 561922 561622 561978
rect 561678 561922 561774 561978
rect 561154 544350 561774 561922
rect 561154 544294 561250 544350
rect 561306 544294 561374 544350
rect 561430 544294 561498 544350
rect 561554 544294 561622 544350
rect 561678 544294 561774 544350
rect 561154 544226 561774 544294
rect 561154 544170 561250 544226
rect 561306 544170 561374 544226
rect 561430 544170 561498 544226
rect 561554 544170 561622 544226
rect 561678 544170 561774 544226
rect 561154 544102 561774 544170
rect 561154 544046 561250 544102
rect 561306 544046 561374 544102
rect 561430 544046 561498 544102
rect 561554 544046 561622 544102
rect 561678 544046 561774 544102
rect 561154 543978 561774 544046
rect 561154 543922 561250 543978
rect 561306 543922 561374 543978
rect 561430 543922 561498 543978
rect 561554 543922 561622 543978
rect 561678 543922 561774 543978
rect 561154 526350 561774 543922
rect 561154 526294 561250 526350
rect 561306 526294 561374 526350
rect 561430 526294 561498 526350
rect 561554 526294 561622 526350
rect 561678 526294 561774 526350
rect 561154 526226 561774 526294
rect 561154 526170 561250 526226
rect 561306 526170 561374 526226
rect 561430 526170 561498 526226
rect 561554 526170 561622 526226
rect 561678 526170 561774 526226
rect 561154 526102 561774 526170
rect 561154 526046 561250 526102
rect 561306 526046 561374 526102
rect 561430 526046 561498 526102
rect 561554 526046 561622 526102
rect 561678 526046 561774 526102
rect 561154 525978 561774 526046
rect 561154 525922 561250 525978
rect 561306 525922 561374 525978
rect 561430 525922 561498 525978
rect 561554 525922 561622 525978
rect 561678 525922 561774 525978
rect 561154 508350 561774 525922
rect 561154 508294 561250 508350
rect 561306 508294 561374 508350
rect 561430 508294 561498 508350
rect 561554 508294 561622 508350
rect 561678 508294 561774 508350
rect 561154 508226 561774 508294
rect 561154 508170 561250 508226
rect 561306 508170 561374 508226
rect 561430 508170 561498 508226
rect 561554 508170 561622 508226
rect 561678 508170 561774 508226
rect 561154 508102 561774 508170
rect 561154 508046 561250 508102
rect 561306 508046 561374 508102
rect 561430 508046 561498 508102
rect 561554 508046 561622 508102
rect 561678 508046 561774 508102
rect 561154 507978 561774 508046
rect 561154 507922 561250 507978
rect 561306 507922 561374 507978
rect 561430 507922 561498 507978
rect 561554 507922 561622 507978
rect 561678 507922 561774 507978
rect 561154 490350 561774 507922
rect 564874 598172 565494 598268
rect 564874 598116 564970 598172
rect 565026 598116 565094 598172
rect 565150 598116 565218 598172
rect 565274 598116 565342 598172
rect 565398 598116 565494 598172
rect 564874 598048 565494 598116
rect 564874 597992 564970 598048
rect 565026 597992 565094 598048
rect 565150 597992 565218 598048
rect 565274 597992 565342 598048
rect 565398 597992 565494 598048
rect 564874 597924 565494 597992
rect 564874 597868 564970 597924
rect 565026 597868 565094 597924
rect 565150 597868 565218 597924
rect 565274 597868 565342 597924
rect 565398 597868 565494 597924
rect 564874 597800 565494 597868
rect 564874 597744 564970 597800
rect 565026 597744 565094 597800
rect 565150 597744 565218 597800
rect 565274 597744 565342 597800
rect 565398 597744 565494 597800
rect 564874 586350 565494 597744
rect 564874 586294 564970 586350
rect 565026 586294 565094 586350
rect 565150 586294 565218 586350
rect 565274 586294 565342 586350
rect 565398 586294 565494 586350
rect 564874 586226 565494 586294
rect 564874 586170 564970 586226
rect 565026 586170 565094 586226
rect 565150 586170 565218 586226
rect 565274 586170 565342 586226
rect 565398 586170 565494 586226
rect 564874 586102 565494 586170
rect 564874 586046 564970 586102
rect 565026 586046 565094 586102
rect 565150 586046 565218 586102
rect 565274 586046 565342 586102
rect 565398 586046 565494 586102
rect 564874 585978 565494 586046
rect 564874 585922 564970 585978
rect 565026 585922 565094 585978
rect 565150 585922 565218 585978
rect 565274 585922 565342 585978
rect 565398 585922 565494 585978
rect 564874 568350 565494 585922
rect 564874 568294 564970 568350
rect 565026 568294 565094 568350
rect 565150 568294 565218 568350
rect 565274 568294 565342 568350
rect 565398 568294 565494 568350
rect 564874 568226 565494 568294
rect 564874 568170 564970 568226
rect 565026 568170 565094 568226
rect 565150 568170 565218 568226
rect 565274 568170 565342 568226
rect 565398 568170 565494 568226
rect 564874 568102 565494 568170
rect 564874 568046 564970 568102
rect 565026 568046 565094 568102
rect 565150 568046 565218 568102
rect 565274 568046 565342 568102
rect 565398 568046 565494 568102
rect 564874 567978 565494 568046
rect 564874 567922 564970 567978
rect 565026 567922 565094 567978
rect 565150 567922 565218 567978
rect 565274 567922 565342 567978
rect 565398 567922 565494 567978
rect 564874 550350 565494 567922
rect 564874 550294 564970 550350
rect 565026 550294 565094 550350
rect 565150 550294 565218 550350
rect 565274 550294 565342 550350
rect 565398 550294 565494 550350
rect 564874 550226 565494 550294
rect 564874 550170 564970 550226
rect 565026 550170 565094 550226
rect 565150 550170 565218 550226
rect 565274 550170 565342 550226
rect 565398 550170 565494 550226
rect 564874 550102 565494 550170
rect 564874 550046 564970 550102
rect 565026 550046 565094 550102
rect 565150 550046 565218 550102
rect 565274 550046 565342 550102
rect 565398 550046 565494 550102
rect 564874 549978 565494 550046
rect 564874 549922 564970 549978
rect 565026 549922 565094 549978
rect 565150 549922 565218 549978
rect 565274 549922 565342 549978
rect 565398 549922 565494 549978
rect 564874 532350 565494 549922
rect 564874 532294 564970 532350
rect 565026 532294 565094 532350
rect 565150 532294 565218 532350
rect 565274 532294 565342 532350
rect 565398 532294 565494 532350
rect 564874 532226 565494 532294
rect 564874 532170 564970 532226
rect 565026 532170 565094 532226
rect 565150 532170 565218 532226
rect 565274 532170 565342 532226
rect 565398 532170 565494 532226
rect 564874 532102 565494 532170
rect 564874 532046 564970 532102
rect 565026 532046 565094 532102
rect 565150 532046 565218 532102
rect 565274 532046 565342 532102
rect 565398 532046 565494 532102
rect 564874 531978 565494 532046
rect 564874 531922 564970 531978
rect 565026 531922 565094 531978
rect 565150 531922 565218 531978
rect 565274 531922 565342 531978
rect 565398 531922 565494 531978
rect 564874 514350 565494 531922
rect 564874 514294 564970 514350
rect 565026 514294 565094 514350
rect 565150 514294 565218 514350
rect 565274 514294 565342 514350
rect 565398 514294 565494 514350
rect 564874 514226 565494 514294
rect 564874 514170 564970 514226
rect 565026 514170 565094 514226
rect 565150 514170 565218 514226
rect 565274 514170 565342 514226
rect 565398 514170 565494 514226
rect 564874 514102 565494 514170
rect 564874 514046 564970 514102
rect 565026 514046 565094 514102
rect 565150 514046 565218 514102
rect 565274 514046 565342 514102
rect 565398 514046 565494 514102
rect 564874 513978 565494 514046
rect 564874 513922 564970 513978
rect 565026 513922 565094 513978
rect 565150 513922 565218 513978
rect 565274 513922 565342 513978
rect 565398 513922 565494 513978
rect 564874 500556 565494 513922
rect 579154 597212 579774 598268
rect 579154 597156 579250 597212
rect 579306 597156 579374 597212
rect 579430 597156 579498 597212
rect 579554 597156 579622 597212
rect 579678 597156 579774 597212
rect 579154 597088 579774 597156
rect 579154 597032 579250 597088
rect 579306 597032 579374 597088
rect 579430 597032 579498 597088
rect 579554 597032 579622 597088
rect 579678 597032 579774 597088
rect 579154 596964 579774 597032
rect 579154 596908 579250 596964
rect 579306 596908 579374 596964
rect 579430 596908 579498 596964
rect 579554 596908 579622 596964
rect 579678 596908 579774 596964
rect 579154 596840 579774 596908
rect 579154 596784 579250 596840
rect 579306 596784 579374 596840
rect 579430 596784 579498 596840
rect 579554 596784 579622 596840
rect 579678 596784 579774 596840
rect 579154 580350 579774 596784
rect 579154 580294 579250 580350
rect 579306 580294 579374 580350
rect 579430 580294 579498 580350
rect 579554 580294 579622 580350
rect 579678 580294 579774 580350
rect 579154 580226 579774 580294
rect 579154 580170 579250 580226
rect 579306 580170 579374 580226
rect 579430 580170 579498 580226
rect 579554 580170 579622 580226
rect 579678 580170 579774 580226
rect 579154 580102 579774 580170
rect 579154 580046 579250 580102
rect 579306 580046 579374 580102
rect 579430 580046 579498 580102
rect 579554 580046 579622 580102
rect 579678 580046 579774 580102
rect 579154 579978 579774 580046
rect 579154 579922 579250 579978
rect 579306 579922 579374 579978
rect 579430 579922 579498 579978
rect 579554 579922 579622 579978
rect 579678 579922 579774 579978
rect 579154 562350 579774 579922
rect 579154 562294 579250 562350
rect 579306 562294 579374 562350
rect 579430 562294 579498 562350
rect 579554 562294 579622 562350
rect 579678 562294 579774 562350
rect 579154 562226 579774 562294
rect 579154 562170 579250 562226
rect 579306 562170 579374 562226
rect 579430 562170 579498 562226
rect 579554 562170 579622 562226
rect 579678 562170 579774 562226
rect 579154 562102 579774 562170
rect 579154 562046 579250 562102
rect 579306 562046 579374 562102
rect 579430 562046 579498 562102
rect 579554 562046 579622 562102
rect 579678 562046 579774 562102
rect 579154 561978 579774 562046
rect 579154 561922 579250 561978
rect 579306 561922 579374 561978
rect 579430 561922 579498 561978
rect 579554 561922 579622 561978
rect 579678 561922 579774 561978
rect 579154 544350 579774 561922
rect 579154 544294 579250 544350
rect 579306 544294 579374 544350
rect 579430 544294 579498 544350
rect 579554 544294 579622 544350
rect 579678 544294 579774 544350
rect 579154 544226 579774 544294
rect 579154 544170 579250 544226
rect 579306 544170 579374 544226
rect 579430 544170 579498 544226
rect 579554 544170 579622 544226
rect 579678 544170 579774 544226
rect 579154 544102 579774 544170
rect 579154 544046 579250 544102
rect 579306 544046 579374 544102
rect 579430 544046 579498 544102
rect 579554 544046 579622 544102
rect 579678 544046 579774 544102
rect 579154 543978 579774 544046
rect 579154 543922 579250 543978
rect 579306 543922 579374 543978
rect 579430 543922 579498 543978
rect 579554 543922 579622 543978
rect 579678 543922 579774 543978
rect 579154 526350 579774 543922
rect 579154 526294 579250 526350
rect 579306 526294 579374 526350
rect 579430 526294 579498 526350
rect 579554 526294 579622 526350
rect 579678 526294 579774 526350
rect 579154 526226 579774 526294
rect 579154 526170 579250 526226
rect 579306 526170 579374 526226
rect 579430 526170 579498 526226
rect 579554 526170 579622 526226
rect 579678 526170 579774 526226
rect 579154 526102 579774 526170
rect 579154 526046 579250 526102
rect 579306 526046 579374 526102
rect 579430 526046 579498 526102
rect 579554 526046 579622 526102
rect 579678 526046 579774 526102
rect 579154 525978 579774 526046
rect 579154 525922 579250 525978
rect 579306 525922 579374 525978
rect 579430 525922 579498 525978
rect 579554 525922 579622 525978
rect 579678 525922 579774 525978
rect 579154 508350 579774 525922
rect 579154 508294 579250 508350
rect 579306 508294 579374 508350
rect 579430 508294 579498 508350
rect 579554 508294 579622 508350
rect 579678 508294 579774 508350
rect 579154 508226 579774 508294
rect 579154 508170 579250 508226
rect 579306 508170 579374 508226
rect 579430 508170 579498 508226
rect 579554 508170 579622 508226
rect 579678 508170 579774 508226
rect 579154 508102 579774 508170
rect 579154 508046 579250 508102
rect 579306 508046 579374 508102
rect 579430 508046 579498 508102
rect 579554 508046 579622 508102
rect 579678 508046 579774 508102
rect 579154 507978 579774 508046
rect 579154 507922 579250 507978
rect 579306 507922 579374 507978
rect 579430 507922 579498 507978
rect 579554 507922 579622 507978
rect 579678 507922 579774 507978
rect 567988 496350 568308 496384
rect 567988 496294 568058 496350
rect 568114 496294 568182 496350
rect 568238 496294 568308 496350
rect 567988 496226 568308 496294
rect 567988 496170 568058 496226
rect 568114 496170 568182 496226
rect 568238 496170 568308 496226
rect 567988 496102 568308 496170
rect 567988 496046 568058 496102
rect 568114 496046 568182 496102
rect 568238 496046 568308 496102
rect 567988 495978 568308 496046
rect 567988 495922 568058 495978
rect 568114 495922 568182 495978
rect 568238 495922 568308 495978
rect 567988 495888 568308 495922
rect 574792 496350 575112 496384
rect 574792 496294 574862 496350
rect 574918 496294 574986 496350
rect 575042 496294 575112 496350
rect 574792 496226 575112 496294
rect 574792 496170 574862 496226
rect 574918 496170 574986 496226
rect 575042 496170 575112 496226
rect 574792 496102 575112 496170
rect 574792 496046 574862 496102
rect 574918 496046 574986 496102
rect 575042 496046 575112 496102
rect 574792 495978 575112 496046
rect 574792 495922 574862 495978
rect 574918 495922 574986 495978
rect 575042 495922 575112 495978
rect 574792 495888 575112 495922
rect 561154 490294 561250 490350
rect 561306 490294 561374 490350
rect 561430 490294 561498 490350
rect 561554 490294 561622 490350
rect 561678 490294 561774 490350
rect 561154 490226 561774 490294
rect 561154 490170 561250 490226
rect 561306 490170 561374 490226
rect 561430 490170 561498 490226
rect 561554 490170 561622 490226
rect 561678 490170 561774 490226
rect 561154 490102 561774 490170
rect 561154 490046 561250 490102
rect 561306 490046 561374 490102
rect 561430 490046 561498 490102
rect 561554 490046 561622 490102
rect 561678 490046 561774 490102
rect 561154 489978 561774 490046
rect 561154 489922 561250 489978
rect 561306 489922 561374 489978
rect 561430 489922 561498 489978
rect 561554 489922 561622 489978
rect 561678 489922 561774 489978
rect 561154 487822 561774 489922
rect 564586 490350 564906 490384
rect 564586 490294 564656 490350
rect 564712 490294 564780 490350
rect 564836 490294 564906 490350
rect 564586 490226 564906 490294
rect 564586 490170 564656 490226
rect 564712 490170 564780 490226
rect 564836 490170 564906 490226
rect 564586 490102 564906 490170
rect 564586 490046 564656 490102
rect 564712 490046 564780 490102
rect 564836 490046 564906 490102
rect 564586 489978 564906 490046
rect 564586 489922 564656 489978
rect 564712 489922 564780 489978
rect 564836 489922 564906 489978
rect 564586 489888 564906 489922
rect 571390 490350 571710 490384
rect 571390 490294 571460 490350
rect 571516 490294 571584 490350
rect 571640 490294 571710 490350
rect 571390 490226 571710 490294
rect 571390 490170 571460 490226
rect 571516 490170 571584 490226
rect 571640 490170 571710 490226
rect 571390 490102 571710 490170
rect 571390 490046 571460 490102
rect 571516 490046 571584 490102
rect 571640 490046 571710 490102
rect 571390 489978 571710 490046
rect 571390 489922 571460 489978
rect 571516 489922 571584 489978
rect 571640 489922 571710 489978
rect 571390 489888 571710 489922
rect 578194 490350 578514 490384
rect 578194 490294 578264 490350
rect 578320 490294 578388 490350
rect 578444 490294 578514 490350
rect 578194 490226 578514 490294
rect 578194 490170 578264 490226
rect 578320 490170 578388 490226
rect 578444 490170 578514 490226
rect 578194 490102 578514 490170
rect 578194 490046 578264 490102
rect 578320 490046 578388 490102
rect 578444 490046 578514 490102
rect 578194 489978 578514 490046
rect 578194 489922 578264 489978
rect 578320 489922 578388 489978
rect 578444 489922 578514 489978
rect 578194 489888 578514 489922
rect 579154 490350 579774 507922
rect 582874 598172 583494 598268
rect 582874 598116 582970 598172
rect 583026 598116 583094 598172
rect 583150 598116 583218 598172
rect 583274 598116 583342 598172
rect 583398 598116 583494 598172
rect 582874 598048 583494 598116
rect 582874 597992 582970 598048
rect 583026 597992 583094 598048
rect 583150 597992 583218 598048
rect 583274 597992 583342 598048
rect 583398 597992 583494 598048
rect 582874 597924 583494 597992
rect 582874 597868 582970 597924
rect 583026 597868 583094 597924
rect 583150 597868 583218 597924
rect 583274 597868 583342 597924
rect 583398 597868 583494 597924
rect 582874 597800 583494 597868
rect 582874 597744 582970 597800
rect 583026 597744 583094 597800
rect 583150 597744 583218 597800
rect 583274 597744 583342 597800
rect 583398 597744 583494 597800
rect 582874 586350 583494 597744
rect 597360 598172 597980 598268
rect 597360 598116 597456 598172
rect 597512 598116 597580 598172
rect 597636 598116 597704 598172
rect 597760 598116 597828 598172
rect 597884 598116 597980 598172
rect 597360 598048 597980 598116
rect 597360 597992 597456 598048
rect 597512 597992 597580 598048
rect 597636 597992 597704 598048
rect 597760 597992 597828 598048
rect 597884 597992 597980 598048
rect 597360 597924 597980 597992
rect 597360 597868 597456 597924
rect 597512 597868 597580 597924
rect 597636 597868 597704 597924
rect 597760 597868 597828 597924
rect 597884 597868 597980 597924
rect 597360 597800 597980 597868
rect 597360 597744 597456 597800
rect 597512 597744 597580 597800
rect 597636 597744 597704 597800
rect 597760 597744 597828 597800
rect 597884 597744 597980 597800
rect 582874 586294 582970 586350
rect 583026 586294 583094 586350
rect 583150 586294 583218 586350
rect 583274 586294 583342 586350
rect 583398 586294 583494 586350
rect 582874 586226 583494 586294
rect 582874 586170 582970 586226
rect 583026 586170 583094 586226
rect 583150 586170 583218 586226
rect 583274 586170 583342 586226
rect 583398 586170 583494 586226
rect 582874 586102 583494 586170
rect 582874 586046 582970 586102
rect 583026 586046 583094 586102
rect 583150 586046 583218 586102
rect 583274 586046 583342 586102
rect 583398 586046 583494 586102
rect 582874 585978 583494 586046
rect 582874 585922 582970 585978
rect 583026 585922 583094 585978
rect 583150 585922 583218 585978
rect 583274 585922 583342 585978
rect 583398 585922 583494 585978
rect 582874 568350 583494 585922
rect 582874 568294 582970 568350
rect 583026 568294 583094 568350
rect 583150 568294 583218 568350
rect 583274 568294 583342 568350
rect 583398 568294 583494 568350
rect 582874 568226 583494 568294
rect 582874 568170 582970 568226
rect 583026 568170 583094 568226
rect 583150 568170 583218 568226
rect 583274 568170 583342 568226
rect 583398 568170 583494 568226
rect 582874 568102 583494 568170
rect 582874 568046 582970 568102
rect 583026 568046 583094 568102
rect 583150 568046 583218 568102
rect 583274 568046 583342 568102
rect 583398 568046 583494 568102
rect 582874 567978 583494 568046
rect 582874 567922 582970 567978
rect 583026 567922 583094 567978
rect 583150 567922 583218 567978
rect 583274 567922 583342 567978
rect 583398 567922 583494 567978
rect 582874 550350 583494 567922
rect 582874 550294 582970 550350
rect 583026 550294 583094 550350
rect 583150 550294 583218 550350
rect 583274 550294 583342 550350
rect 583398 550294 583494 550350
rect 582874 550226 583494 550294
rect 582874 550170 582970 550226
rect 583026 550170 583094 550226
rect 583150 550170 583218 550226
rect 583274 550170 583342 550226
rect 583398 550170 583494 550226
rect 582874 550102 583494 550170
rect 582874 550046 582970 550102
rect 583026 550046 583094 550102
rect 583150 550046 583218 550102
rect 583274 550046 583342 550102
rect 583398 550046 583494 550102
rect 582874 549978 583494 550046
rect 582874 549922 582970 549978
rect 583026 549922 583094 549978
rect 583150 549922 583218 549978
rect 583274 549922 583342 549978
rect 583398 549922 583494 549978
rect 582874 532350 583494 549922
rect 582874 532294 582970 532350
rect 583026 532294 583094 532350
rect 583150 532294 583218 532350
rect 583274 532294 583342 532350
rect 583398 532294 583494 532350
rect 582874 532226 583494 532294
rect 582874 532170 582970 532226
rect 583026 532170 583094 532226
rect 583150 532170 583218 532226
rect 583274 532170 583342 532226
rect 583398 532170 583494 532226
rect 582874 532102 583494 532170
rect 582874 532046 582970 532102
rect 583026 532046 583094 532102
rect 583150 532046 583218 532102
rect 583274 532046 583342 532102
rect 583398 532046 583494 532102
rect 582874 531978 583494 532046
rect 582874 531922 582970 531978
rect 583026 531922 583094 531978
rect 583150 531922 583218 531978
rect 583274 531922 583342 531978
rect 583398 531922 583494 531978
rect 582874 514350 583494 531922
rect 582874 514294 582970 514350
rect 583026 514294 583094 514350
rect 583150 514294 583218 514350
rect 583274 514294 583342 514350
rect 583398 514294 583494 514350
rect 582874 514226 583494 514294
rect 582874 514170 582970 514226
rect 583026 514170 583094 514226
rect 583150 514170 583218 514226
rect 583274 514170 583342 514226
rect 583398 514170 583494 514226
rect 582874 514102 583494 514170
rect 582874 514046 582970 514102
rect 583026 514046 583094 514102
rect 583150 514046 583218 514102
rect 583274 514046 583342 514102
rect 583398 514046 583494 514102
rect 582874 513978 583494 514046
rect 582874 513922 582970 513978
rect 583026 513922 583094 513978
rect 583150 513922 583218 513978
rect 583274 513922 583342 513978
rect 583398 513922 583494 513978
rect 581596 496350 581916 496384
rect 581596 496294 581666 496350
rect 581722 496294 581790 496350
rect 581846 496294 581916 496350
rect 581596 496226 581916 496294
rect 581596 496170 581666 496226
rect 581722 496170 581790 496226
rect 581846 496170 581916 496226
rect 581596 496102 581916 496170
rect 581596 496046 581666 496102
rect 581722 496046 581790 496102
rect 581846 496046 581916 496102
rect 581596 495978 581916 496046
rect 581596 495922 581666 495978
rect 581722 495922 581790 495978
rect 581846 495922 581916 495978
rect 581596 495888 581916 495922
rect 582874 496350 583494 513922
rect 596400 597212 597020 597308
rect 596400 597156 596496 597212
rect 596552 597156 596620 597212
rect 596676 597156 596744 597212
rect 596800 597156 596868 597212
rect 596924 597156 597020 597212
rect 596400 597088 597020 597156
rect 596400 597032 596496 597088
rect 596552 597032 596620 597088
rect 596676 597032 596744 597088
rect 596800 597032 596868 597088
rect 596924 597032 597020 597088
rect 596400 596964 597020 597032
rect 596400 596908 596496 596964
rect 596552 596908 596620 596964
rect 596676 596908 596744 596964
rect 596800 596908 596868 596964
rect 596924 596908 597020 596964
rect 596400 596840 597020 596908
rect 596400 596784 596496 596840
rect 596552 596784 596620 596840
rect 596676 596784 596744 596840
rect 596800 596784 596868 596840
rect 596924 596784 597020 596840
rect 596400 580350 597020 596784
rect 596400 580294 596496 580350
rect 596552 580294 596620 580350
rect 596676 580294 596744 580350
rect 596800 580294 596868 580350
rect 596924 580294 597020 580350
rect 596400 580226 597020 580294
rect 596400 580170 596496 580226
rect 596552 580170 596620 580226
rect 596676 580170 596744 580226
rect 596800 580170 596868 580226
rect 596924 580170 597020 580226
rect 596400 580102 597020 580170
rect 596400 580046 596496 580102
rect 596552 580046 596620 580102
rect 596676 580046 596744 580102
rect 596800 580046 596868 580102
rect 596924 580046 597020 580102
rect 596400 579978 597020 580046
rect 596400 579922 596496 579978
rect 596552 579922 596620 579978
rect 596676 579922 596744 579978
rect 596800 579922 596868 579978
rect 596924 579922 597020 579978
rect 596400 562350 597020 579922
rect 596400 562294 596496 562350
rect 596552 562294 596620 562350
rect 596676 562294 596744 562350
rect 596800 562294 596868 562350
rect 596924 562294 597020 562350
rect 596400 562226 597020 562294
rect 596400 562170 596496 562226
rect 596552 562170 596620 562226
rect 596676 562170 596744 562226
rect 596800 562170 596868 562226
rect 596924 562170 597020 562226
rect 596400 562102 597020 562170
rect 596400 562046 596496 562102
rect 596552 562046 596620 562102
rect 596676 562046 596744 562102
rect 596800 562046 596868 562102
rect 596924 562046 597020 562102
rect 596400 561978 597020 562046
rect 596400 561922 596496 561978
rect 596552 561922 596620 561978
rect 596676 561922 596744 561978
rect 596800 561922 596868 561978
rect 596924 561922 597020 561978
rect 596400 544350 597020 561922
rect 596400 544294 596496 544350
rect 596552 544294 596620 544350
rect 596676 544294 596744 544350
rect 596800 544294 596868 544350
rect 596924 544294 597020 544350
rect 596400 544226 597020 544294
rect 596400 544170 596496 544226
rect 596552 544170 596620 544226
rect 596676 544170 596744 544226
rect 596800 544170 596868 544226
rect 596924 544170 597020 544226
rect 596400 544102 597020 544170
rect 596400 544046 596496 544102
rect 596552 544046 596620 544102
rect 596676 544046 596744 544102
rect 596800 544046 596868 544102
rect 596924 544046 597020 544102
rect 596400 543978 597020 544046
rect 596400 543922 596496 543978
rect 596552 543922 596620 543978
rect 596676 543922 596744 543978
rect 596800 543922 596868 543978
rect 596924 543922 597020 543978
rect 596400 526350 597020 543922
rect 596400 526294 596496 526350
rect 596552 526294 596620 526350
rect 596676 526294 596744 526350
rect 596800 526294 596868 526350
rect 596924 526294 597020 526350
rect 596400 526226 597020 526294
rect 596400 526170 596496 526226
rect 596552 526170 596620 526226
rect 596676 526170 596744 526226
rect 596800 526170 596868 526226
rect 596924 526170 597020 526226
rect 596400 526102 597020 526170
rect 596400 526046 596496 526102
rect 596552 526046 596620 526102
rect 596676 526046 596744 526102
rect 596800 526046 596868 526102
rect 596924 526046 597020 526102
rect 596400 525978 597020 526046
rect 596400 525922 596496 525978
rect 596552 525922 596620 525978
rect 596676 525922 596744 525978
rect 596800 525922 596868 525978
rect 596924 525922 597020 525978
rect 596400 508350 597020 525922
rect 596400 508294 596496 508350
rect 596552 508294 596620 508350
rect 596676 508294 596744 508350
rect 596800 508294 596868 508350
rect 596924 508294 597020 508350
rect 596400 508226 597020 508294
rect 596400 508170 596496 508226
rect 596552 508170 596620 508226
rect 596676 508170 596744 508226
rect 596800 508170 596868 508226
rect 596924 508170 597020 508226
rect 596400 508102 597020 508170
rect 596400 508046 596496 508102
rect 596552 508046 596620 508102
rect 596676 508046 596744 508102
rect 596800 508046 596868 508102
rect 596924 508046 597020 508102
rect 596400 507978 597020 508046
rect 596400 507922 596496 507978
rect 596552 507922 596620 507978
rect 596676 507922 596744 507978
rect 596800 507922 596868 507978
rect 596924 507922 597020 507978
rect 582874 496294 582970 496350
rect 583026 496294 583094 496350
rect 583150 496294 583218 496350
rect 583274 496294 583342 496350
rect 583398 496294 583494 496350
rect 582874 496226 583494 496294
rect 582874 496170 582970 496226
rect 583026 496170 583094 496226
rect 583150 496170 583218 496226
rect 583274 496170 583342 496226
rect 583398 496170 583494 496226
rect 582874 496102 583494 496170
rect 582874 496046 582970 496102
rect 583026 496046 583094 496102
rect 583150 496046 583218 496102
rect 583274 496046 583342 496102
rect 583398 496046 583494 496102
rect 582874 495978 583494 496046
rect 582874 495922 582970 495978
rect 583026 495922 583094 495978
rect 583150 495922 583218 495978
rect 583274 495922 583342 495978
rect 583398 495922 583494 495978
rect 579154 490294 579250 490350
rect 579306 490294 579374 490350
rect 579430 490294 579498 490350
rect 579554 490294 579622 490350
rect 579678 490294 579774 490350
rect 579154 490226 579774 490294
rect 579154 490170 579250 490226
rect 579306 490170 579374 490226
rect 579430 490170 579498 490226
rect 579554 490170 579622 490226
rect 579678 490170 579774 490226
rect 579154 490102 579774 490170
rect 579154 490046 579250 490102
rect 579306 490046 579374 490102
rect 579430 490046 579498 490102
rect 579554 490046 579622 490102
rect 579678 490046 579774 490102
rect 579154 489978 579774 490046
rect 579154 489922 579250 489978
rect 579306 489922 579374 489978
rect 579430 489922 579498 489978
rect 579554 489922 579622 489978
rect 579678 489922 579774 489978
rect 579154 487822 579774 489922
rect 582874 487822 583494 495922
rect 588400 496350 588720 496384
rect 588400 496294 588470 496350
rect 588526 496294 588594 496350
rect 588650 496294 588720 496350
rect 588400 496226 588720 496294
rect 588400 496170 588470 496226
rect 588526 496170 588594 496226
rect 588650 496170 588720 496226
rect 588400 496102 588720 496170
rect 588400 496046 588470 496102
rect 588526 496046 588594 496102
rect 588650 496046 588720 496102
rect 588400 495978 588720 496046
rect 588400 495922 588470 495978
rect 588526 495922 588594 495978
rect 588650 495922 588720 495978
rect 588400 495888 588720 495922
rect 584998 490350 585318 490384
rect 584998 490294 585068 490350
rect 585124 490294 585192 490350
rect 585248 490294 585318 490350
rect 584998 490226 585318 490294
rect 584998 490170 585068 490226
rect 585124 490170 585192 490226
rect 585248 490170 585318 490226
rect 584998 490102 585318 490170
rect 584998 490046 585068 490102
rect 585124 490046 585192 490102
rect 585248 490046 585318 490102
rect 584998 489978 585318 490046
rect 584998 489922 585068 489978
rect 585124 489922 585192 489978
rect 585248 489922 585318 489978
rect 584998 489888 585318 489922
rect 596400 490350 597020 507922
rect 596400 490294 596496 490350
rect 596552 490294 596620 490350
rect 596676 490294 596744 490350
rect 596800 490294 596868 490350
rect 596924 490294 597020 490350
rect 596400 490226 597020 490294
rect 596400 490170 596496 490226
rect 596552 490170 596620 490226
rect 596676 490170 596744 490226
rect 596800 490170 596868 490226
rect 596924 490170 597020 490226
rect 596400 490102 597020 490170
rect 596400 490046 596496 490102
rect 596552 490046 596620 490102
rect 596676 490046 596744 490102
rect 596800 490046 596868 490102
rect 596924 490046 597020 490102
rect 596400 489978 597020 490046
rect 596400 489922 596496 489978
rect 596552 489922 596620 489978
rect 596676 489922 596744 489978
rect 596800 489922 596868 489978
rect 596924 489922 597020 489978
rect 546874 478294 546970 478350
rect 547026 478294 547094 478350
rect 547150 478294 547218 478350
rect 547274 478294 547342 478350
rect 547398 478294 547494 478350
rect 546874 478226 547494 478294
rect 546874 478170 546970 478226
rect 547026 478170 547094 478226
rect 547150 478170 547218 478226
rect 547274 478170 547342 478226
rect 547398 478170 547494 478226
rect 546874 478102 547494 478170
rect 546874 478046 546970 478102
rect 547026 478046 547094 478102
rect 547150 478046 547218 478102
rect 547274 478046 547342 478102
rect 547398 478046 547494 478102
rect 546874 477978 547494 478046
rect 546874 477922 546970 477978
rect 547026 477922 547094 477978
rect 547150 477922 547218 477978
rect 547274 477922 547342 477978
rect 547398 477922 547494 477978
rect 546874 460350 547494 477922
rect 567988 478350 568308 478384
rect 567988 478294 568058 478350
rect 568114 478294 568182 478350
rect 568238 478294 568308 478350
rect 567988 478226 568308 478294
rect 567988 478170 568058 478226
rect 568114 478170 568182 478226
rect 568238 478170 568308 478226
rect 567988 478102 568308 478170
rect 567988 478046 568058 478102
rect 568114 478046 568182 478102
rect 568238 478046 568308 478102
rect 567988 477978 568308 478046
rect 567988 477922 568058 477978
rect 568114 477922 568182 477978
rect 568238 477922 568308 477978
rect 567988 477888 568308 477922
rect 574792 478350 575112 478384
rect 574792 478294 574862 478350
rect 574918 478294 574986 478350
rect 575042 478294 575112 478350
rect 574792 478226 575112 478294
rect 574792 478170 574862 478226
rect 574918 478170 574986 478226
rect 575042 478170 575112 478226
rect 574792 478102 575112 478170
rect 574792 478046 574862 478102
rect 574918 478046 574986 478102
rect 575042 478046 575112 478102
rect 574792 477978 575112 478046
rect 574792 477922 574862 477978
rect 574918 477922 574986 477978
rect 575042 477922 575112 477978
rect 574792 477888 575112 477922
rect 581596 478350 581916 478384
rect 581596 478294 581666 478350
rect 581722 478294 581790 478350
rect 581846 478294 581916 478350
rect 581596 478226 581916 478294
rect 581596 478170 581666 478226
rect 581722 478170 581790 478226
rect 581846 478170 581916 478226
rect 581596 478102 581916 478170
rect 581596 478046 581666 478102
rect 581722 478046 581790 478102
rect 581846 478046 581916 478102
rect 581596 477978 581916 478046
rect 581596 477922 581666 477978
rect 581722 477922 581790 477978
rect 581846 477922 581916 477978
rect 581596 477888 581916 477922
rect 588400 478350 588720 478384
rect 588400 478294 588470 478350
rect 588526 478294 588594 478350
rect 588650 478294 588720 478350
rect 588400 478226 588720 478294
rect 588400 478170 588470 478226
rect 588526 478170 588594 478226
rect 588650 478170 588720 478226
rect 588400 478102 588720 478170
rect 588400 478046 588470 478102
rect 588526 478046 588594 478102
rect 588650 478046 588720 478102
rect 588400 477978 588720 478046
rect 588400 477922 588470 477978
rect 588526 477922 588594 477978
rect 588650 477922 588720 477978
rect 588400 477888 588720 477922
rect 564586 472350 564906 472384
rect 564586 472294 564656 472350
rect 564712 472294 564780 472350
rect 564836 472294 564906 472350
rect 564586 472226 564906 472294
rect 564586 472170 564656 472226
rect 564712 472170 564780 472226
rect 564836 472170 564906 472226
rect 564586 472102 564906 472170
rect 564586 472046 564656 472102
rect 564712 472046 564780 472102
rect 564836 472046 564906 472102
rect 564586 471978 564906 472046
rect 564586 471922 564656 471978
rect 564712 471922 564780 471978
rect 564836 471922 564906 471978
rect 564586 471888 564906 471922
rect 571390 472350 571710 472384
rect 571390 472294 571460 472350
rect 571516 472294 571584 472350
rect 571640 472294 571710 472350
rect 571390 472226 571710 472294
rect 571390 472170 571460 472226
rect 571516 472170 571584 472226
rect 571640 472170 571710 472226
rect 571390 472102 571710 472170
rect 571390 472046 571460 472102
rect 571516 472046 571584 472102
rect 571640 472046 571710 472102
rect 571390 471978 571710 472046
rect 571390 471922 571460 471978
rect 571516 471922 571584 471978
rect 571640 471922 571710 471978
rect 571390 471888 571710 471922
rect 578194 472350 578514 472384
rect 578194 472294 578264 472350
rect 578320 472294 578388 472350
rect 578444 472294 578514 472350
rect 578194 472226 578514 472294
rect 578194 472170 578264 472226
rect 578320 472170 578388 472226
rect 578444 472170 578514 472226
rect 578194 472102 578514 472170
rect 578194 472046 578264 472102
rect 578320 472046 578388 472102
rect 578444 472046 578514 472102
rect 578194 471978 578514 472046
rect 578194 471922 578264 471978
rect 578320 471922 578388 471978
rect 578444 471922 578514 471978
rect 578194 471888 578514 471922
rect 584998 472350 585318 472384
rect 584998 472294 585068 472350
rect 585124 472294 585192 472350
rect 585248 472294 585318 472350
rect 584998 472226 585318 472294
rect 584998 472170 585068 472226
rect 585124 472170 585192 472226
rect 585248 472170 585318 472226
rect 584998 472102 585318 472170
rect 584998 472046 585068 472102
rect 585124 472046 585192 472102
rect 585248 472046 585318 472102
rect 584998 471978 585318 472046
rect 584998 471922 585068 471978
rect 585124 471922 585192 471978
rect 585248 471922 585318 471978
rect 584998 471888 585318 471922
rect 596400 472350 597020 489922
rect 596400 472294 596496 472350
rect 596552 472294 596620 472350
rect 596676 472294 596744 472350
rect 596800 472294 596868 472350
rect 596924 472294 597020 472350
rect 596400 472226 597020 472294
rect 596400 472170 596496 472226
rect 596552 472170 596620 472226
rect 596676 472170 596744 472226
rect 596800 472170 596868 472226
rect 596924 472170 597020 472226
rect 596400 472102 597020 472170
rect 596400 472046 596496 472102
rect 596552 472046 596620 472102
rect 596676 472046 596744 472102
rect 596800 472046 596868 472102
rect 596924 472046 597020 472102
rect 596400 471978 597020 472046
rect 596400 471922 596496 471978
rect 596552 471922 596620 471978
rect 596676 471922 596744 471978
rect 596800 471922 596868 471978
rect 596924 471922 597020 471978
rect 560252 465444 560308 465454
rect 546874 460294 546970 460350
rect 547026 460294 547094 460350
rect 547150 460294 547218 460350
rect 547274 460294 547342 460350
rect 547398 460294 547494 460350
rect 546874 460226 547494 460294
rect 546874 460170 546970 460226
rect 547026 460170 547094 460226
rect 547150 460170 547218 460226
rect 547274 460170 547342 460226
rect 547398 460170 547494 460226
rect 546874 460102 547494 460170
rect 546874 460046 546970 460102
rect 547026 460046 547094 460102
rect 547150 460046 547218 460102
rect 547274 460046 547342 460102
rect 547398 460046 547494 460102
rect 546874 459978 547494 460046
rect 546874 459922 546970 459978
rect 547026 459922 547094 459978
rect 547150 459922 547218 459978
rect 547274 459922 547342 459978
rect 547398 459922 547494 459978
rect 546874 442350 547494 459922
rect 546874 442294 546970 442350
rect 547026 442294 547094 442350
rect 547150 442294 547218 442350
rect 547274 442294 547342 442350
rect 547398 442294 547494 442350
rect 546874 442226 547494 442294
rect 546874 442170 546970 442226
rect 547026 442170 547094 442226
rect 547150 442170 547218 442226
rect 547274 442170 547342 442226
rect 547398 442170 547494 442226
rect 546874 442102 547494 442170
rect 546874 442046 546970 442102
rect 547026 442046 547094 442102
rect 547150 442046 547218 442102
rect 547274 442046 547342 442102
rect 547398 442046 547494 442102
rect 546874 441978 547494 442046
rect 546874 441922 546970 441978
rect 547026 441922 547094 441978
rect 547150 441922 547218 441978
rect 547274 441922 547342 441978
rect 547398 441922 547494 441978
rect 546874 424350 547494 441922
rect 546874 424294 546970 424350
rect 547026 424294 547094 424350
rect 547150 424294 547218 424350
rect 547274 424294 547342 424350
rect 547398 424294 547494 424350
rect 546874 424226 547494 424294
rect 546874 424170 546970 424226
rect 547026 424170 547094 424226
rect 547150 424170 547218 424226
rect 547274 424170 547342 424226
rect 547398 424170 547494 424226
rect 546874 424102 547494 424170
rect 546874 424046 546970 424102
rect 547026 424046 547094 424102
rect 547150 424046 547218 424102
rect 547274 424046 547342 424102
rect 547398 424046 547494 424102
rect 546874 423978 547494 424046
rect 546874 423922 546970 423978
rect 547026 423922 547094 423978
rect 547150 423922 547218 423978
rect 547274 423922 547342 423978
rect 547398 423922 547494 423978
rect 546874 406350 547494 423922
rect 546874 406294 546970 406350
rect 547026 406294 547094 406350
rect 547150 406294 547218 406350
rect 547274 406294 547342 406350
rect 547398 406294 547494 406350
rect 546874 406226 547494 406294
rect 546874 406170 546970 406226
rect 547026 406170 547094 406226
rect 547150 406170 547218 406226
rect 547274 406170 547342 406226
rect 547398 406170 547494 406226
rect 546874 406102 547494 406170
rect 546874 406046 546970 406102
rect 547026 406046 547094 406102
rect 547150 406046 547218 406102
rect 547274 406046 547342 406102
rect 547398 406046 547494 406102
rect 546874 405978 547494 406046
rect 546874 405922 546970 405978
rect 547026 405922 547094 405978
rect 547150 405922 547218 405978
rect 547274 405922 547342 405978
rect 547398 405922 547494 405978
rect 546874 388350 547494 405922
rect 546874 388294 546970 388350
rect 547026 388294 547094 388350
rect 547150 388294 547218 388350
rect 547274 388294 547342 388350
rect 547398 388294 547494 388350
rect 546874 388226 547494 388294
rect 546874 388170 546970 388226
rect 547026 388170 547094 388226
rect 547150 388170 547218 388226
rect 547274 388170 547342 388226
rect 547398 388170 547494 388226
rect 546874 388102 547494 388170
rect 546874 388046 546970 388102
rect 547026 388046 547094 388102
rect 547150 388046 547218 388102
rect 547274 388046 547342 388102
rect 547398 388046 547494 388102
rect 546874 387978 547494 388046
rect 546874 387922 546970 387978
rect 547026 387922 547094 387978
rect 547150 387922 547218 387978
rect 547274 387922 547342 387978
rect 547398 387922 547494 387978
rect 546874 370350 547494 387922
rect 549276 462756 549332 462766
rect 546874 370294 546970 370350
rect 547026 370294 547094 370350
rect 547150 370294 547218 370350
rect 547274 370294 547342 370350
rect 547398 370294 547494 370350
rect 546874 370226 547494 370294
rect 546874 370170 546970 370226
rect 547026 370170 547094 370226
rect 547150 370170 547218 370226
rect 547274 370170 547342 370226
rect 547398 370170 547494 370226
rect 546874 370102 547494 370170
rect 546874 370046 546970 370102
rect 547026 370046 547094 370102
rect 547150 370046 547218 370102
rect 547274 370046 547342 370102
rect 547398 370046 547494 370102
rect 546874 369978 547494 370046
rect 546874 369922 546970 369978
rect 547026 369922 547094 369978
rect 547150 369922 547218 369978
rect 547274 369922 547342 369978
rect 547398 369922 547494 369978
rect 546874 352350 547494 369922
rect 546874 352294 546970 352350
rect 547026 352294 547094 352350
rect 547150 352294 547218 352350
rect 547274 352294 547342 352350
rect 547398 352294 547494 352350
rect 546874 352226 547494 352294
rect 546874 352170 546970 352226
rect 547026 352170 547094 352226
rect 547150 352170 547218 352226
rect 547274 352170 547342 352226
rect 547398 352170 547494 352226
rect 546874 352102 547494 352170
rect 546874 352046 546970 352102
rect 547026 352046 547094 352102
rect 547150 352046 547218 352102
rect 547274 352046 547342 352102
rect 547398 352046 547494 352102
rect 546874 351978 547494 352046
rect 546874 351922 546970 351978
rect 547026 351922 547094 351978
rect 547150 351922 547218 351978
rect 547274 351922 547342 351978
rect 547398 351922 547494 351978
rect 546874 334350 547494 351922
rect 546874 334294 546970 334350
rect 547026 334294 547094 334350
rect 547150 334294 547218 334350
rect 547274 334294 547342 334350
rect 547398 334294 547494 334350
rect 546874 334226 547494 334294
rect 546874 334170 546970 334226
rect 547026 334170 547094 334226
rect 547150 334170 547218 334226
rect 547274 334170 547342 334226
rect 547398 334170 547494 334226
rect 546874 334102 547494 334170
rect 546874 334046 546970 334102
rect 547026 334046 547094 334102
rect 547150 334046 547218 334102
rect 547274 334046 547342 334102
rect 547398 334046 547494 334102
rect 546874 333978 547494 334046
rect 546874 333922 546970 333978
rect 547026 333922 547094 333978
rect 547150 333922 547218 333978
rect 547274 333922 547342 333978
rect 547398 333922 547494 333978
rect 546874 316350 547494 333922
rect 546874 316294 546970 316350
rect 547026 316294 547094 316350
rect 547150 316294 547218 316350
rect 547274 316294 547342 316350
rect 547398 316294 547494 316350
rect 546874 316226 547494 316294
rect 546874 316170 546970 316226
rect 547026 316170 547094 316226
rect 547150 316170 547218 316226
rect 547274 316170 547342 316226
rect 547398 316170 547494 316226
rect 546874 316102 547494 316170
rect 546874 316046 546970 316102
rect 547026 316046 547094 316102
rect 547150 316046 547218 316102
rect 547274 316046 547342 316102
rect 547398 316046 547494 316102
rect 546874 315978 547494 316046
rect 546874 315922 546970 315978
rect 547026 315922 547094 315978
rect 547150 315922 547218 315978
rect 547274 315922 547342 315978
rect 547398 315922 547494 315978
rect 546874 298350 547494 315922
rect 546874 298294 546970 298350
rect 547026 298294 547094 298350
rect 547150 298294 547218 298350
rect 547274 298294 547342 298350
rect 547398 298294 547494 298350
rect 546874 298226 547494 298294
rect 546874 298170 546970 298226
rect 547026 298170 547094 298226
rect 547150 298170 547218 298226
rect 547274 298170 547342 298226
rect 547398 298170 547494 298226
rect 546874 298102 547494 298170
rect 546874 298046 546970 298102
rect 547026 298046 547094 298102
rect 547150 298046 547218 298102
rect 547274 298046 547342 298102
rect 547398 298046 547494 298102
rect 546874 297978 547494 298046
rect 546874 297922 546970 297978
rect 547026 297922 547094 297978
rect 547150 297922 547218 297978
rect 547274 297922 547342 297978
rect 547398 297922 547494 297978
rect 546874 280350 547494 297922
rect 546874 280294 546970 280350
rect 547026 280294 547094 280350
rect 547150 280294 547218 280350
rect 547274 280294 547342 280350
rect 547398 280294 547494 280350
rect 546874 280226 547494 280294
rect 546874 280170 546970 280226
rect 547026 280170 547094 280226
rect 547150 280170 547218 280226
rect 547274 280170 547342 280226
rect 547398 280170 547494 280226
rect 546874 280102 547494 280170
rect 546874 280046 546970 280102
rect 547026 280046 547094 280102
rect 547150 280046 547218 280102
rect 547274 280046 547342 280102
rect 547398 280046 547494 280102
rect 546874 279978 547494 280046
rect 546874 279922 546970 279978
rect 547026 279922 547094 279978
rect 547150 279922 547218 279978
rect 547274 279922 547342 279978
rect 547398 279922 547494 279978
rect 546874 262350 547494 279922
rect 546874 262294 546970 262350
rect 547026 262294 547094 262350
rect 547150 262294 547218 262350
rect 547274 262294 547342 262350
rect 547398 262294 547494 262350
rect 546874 262226 547494 262294
rect 546874 262170 546970 262226
rect 547026 262170 547094 262226
rect 547150 262170 547218 262226
rect 547274 262170 547342 262226
rect 547398 262170 547494 262226
rect 546874 262102 547494 262170
rect 546874 262046 546970 262102
rect 547026 262046 547094 262102
rect 547150 262046 547218 262102
rect 547274 262046 547342 262102
rect 547398 262046 547494 262102
rect 546874 261978 547494 262046
rect 546874 261922 546970 261978
rect 547026 261922 547094 261978
rect 547150 261922 547218 261978
rect 547274 261922 547342 261978
rect 547398 261922 547494 261978
rect 546874 244350 547494 261922
rect 546874 244294 546970 244350
rect 547026 244294 547094 244350
rect 547150 244294 547218 244350
rect 547274 244294 547342 244350
rect 547398 244294 547494 244350
rect 546874 244226 547494 244294
rect 546874 244170 546970 244226
rect 547026 244170 547094 244226
rect 547150 244170 547218 244226
rect 547274 244170 547342 244226
rect 547398 244170 547494 244226
rect 546874 244102 547494 244170
rect 546874 244046 546970 244102
rect 547026 244046 547094 244102
rect 547150 244046 547218 244102
rect 547274 244046 547342 244102
rect 547398 244046 547494 244102
rect 546874 243978 547494 244046
rect 546874 243922 546970 243978
rect 547026 243922 547094 243978
rect 547150 243922 547218 243978
rect 547274 243922 547342 243978
rect 547398 243922 547494 243978
rect 546874 226350 547494 243922
rect 546874 226294 546970 226350
rect 547026 226294 547094 226350
rect 547150 226294 547218 226350
rect 547274 226294 547342 226350
rect 547398 226294 547494 226350
rect 546874 226226 547494 226294
rect 546874 226170 546970 226226
rect 547026 226170 547094 226226
rect 547150 226170 547218 226226
rect 547274 226170 547342 226226
rect 547398 226170 547494 226226
rect 546874 226102 547494 226170
rect 546874 226046 546970 226102
rect 547026 226046 547094 226102
rect 547150 226046 547218 226102
rect 547274 226046 547342 226102
rect 547398 226046 547494 226102
rect 546874 225978 547494 226046
rect 546874 225922 546970 225978
rect 547026 225922 547094 225978
rect 547150 225922 547218 225978
rect 547274 225922 547342 225978
rect 547398 225922 547494 225978
rect 546874 217934 547494 225922
rect 549052 377300 549108 377310
rect 348874 208294 348970 208350
rect 349026 208294 349094 208350
rect 349150 208294 349218 208350
rect 349274 208294 349342 208350
rect 349398 208294 349494 208350
rect 348874 208226 349494 208294
rect 348874 208170 348970 208226
rect 349026 208170 349094 208226
rect 349150 208170 349218 208226
rect 349274 208170 349342 208226
rect 349398 208170 349494 208226
rect 348874 208102 349494 208170
rect 348874 208046 348970 208102
rect 349026 208046 349094 208102
rect 349150 208046 349218 208102
rect 349274 208046 349342 208102
rect 349398 208046 349494 208102
rect 348874 207978 349494 208046
rect 348874 207922 348970 207978
rect 349026 207922 349094 207978
rect 349150 207922 349218 207978
rect 349274 207922 349342 207978
rect 349398 207922 349494 207978
rect 348874 190350 349494 207922
rect 363988 208412 365228 208446
rect 363988 208356 364022 208412
rect 364078 208356 364146 208412
rect 364202 208356 364270 208412
rect 364326 208356 364394 208412
rect 364450 208356 364518 208412
rect 364574 208356 364642 208412
rect 364698 208356 364766 208412
rect 364822 208356 364890 208412
rect 364946 208356 365014 208412
rect 365070 208356 365138 208412
rect 365194 208356 365228 208412
rect 363988 208288 365228 208356
rect 363988 208232 364022 208288
rect 364078 208232 364146 208288
rect 364202 208232 364270 208288
rect 364326 208232 364394 208288
rect 364450 208232 364518 208288
rect 364574 208232 364642 208288
rect 364698 208232 364766 208288
rect 364822 208232 364890 208288
rect 364946 208232 365014 208288
rect 365070 208232 365138 208288
rect 365194 208232 365228 208288
rect 363988 208164 365228 208232
rect 363988 208108 364022 208164
rect 364078 208108 364146 208164
rect 364202 208108 364270 208164
rect 364326 208108 364394 208164
rect 364450 208108 364518 208164
rect 364574 208108 364642 208164
rect 364698 208108 364766 208164
rect 364822 208108 364890 208164
rect 364946 208108 365014 208164
rect 365070 208108 365138 208164
rect 365194 208108 365228 208164
rect 363988 208040 365228 208108
rect 363988 207984 364022 208040
rect 364078 207984 364146 208040
rect 364202 207984 364270 208040
rect 364326 207984 364394 208040
rect 364450 207984 364518 208040
rect 364574 207984 364642 208040
rect 364698 207984 364766 208040
rect 364822 207984 364890 208040
rect 364946 207984 365014 208040
rect 365070 207984 365138 208040
rect 365194 207984 365228 208040
rect 363988 207916 365228 207984
rect 363988 207860 364022 207916
rect 364078 207860 364146 207916
rect 364202 207860 364270 207916
rect 364326 207860 364394 207916
rect 364450 207860 364518 207916
rect 364574 207860 364642 207916
rect 364698 207860 364766 207916
rect 364822 207860 364890 207916
rect 364946 207860 365014 207916
rect 365070 207860 365138 207916
rect 365194 207860 365228 207916
rect 363988 207826 365228 207860
rect 383988 208412 385228 208446
rect 383988 208356 384022 208412
rect 384078 208356 384146 208412
rect 384202 208356 384270 208412
rect 384326 208356 384394 208412
rect 384450 208356 384518 208412
rect 384574 208356 384642 208412
rect 384698 208356 384766 208412
rect 384822 208356 384890 208412
rect 384946 208356 385014 208412
rect 385070 208356 385138 208412
rect 385194 208356 385228 208412
rect 383988 208288 385228 208356
rect 383988 208232 384022 208288
rect 384078 208232 384146 208288
rect 384202 208232 384270 208288
rect 384326 208232 384394 208288
rect 384450 208232 384518 208288
rect 384574 208232 384642 208288
rect 384698 208232 384766 208288
rect 384822 208232 384890 208288
rect 384946 208232 385014 208288
rect 385070 208232 385138 208288
rect 385194 208232 385228 208288
rect 383988 208164 385228 208232
rect 383988 208108 384022 208164
rect 384078 208108 384146 208164
rect 384202 208108 384270 208164
rect 384326 208108 384394 208164
rect 384450 208108 384518 208164
rect 384574 208108 384642 208164
rect 384698 208108 384766 208164
rect 384822 208108 384890 208164
rect 384946 208108 385014 208164
rect 385070 208108 385138 208164
rect 385194 208108 385228 208164
rect 383988 208040 385228 208108
rect 383988 207984 384022 208040
rect 384078 207984 384146 208040
rect 384202 207984 384270 208040
rect 384326 207984 384394 208040
rect 384450 207984 384518 208040
rect 384574 207984 384642 208040
rect 384698 207984 384766 208040
rect 384822 207984 384890 208040
rect 384946 207984 385014 208040
rect 385070 207984 385138 208040
rect 385194 207984 385228 208040
rect 383988 207916 385228 207984
rect 383988 207860 384022 207916
rect 384078 207860 384146 207916
rect 384202 207860 384270 207916
rect 384326 207860 384394 207916
rect 384450 207860 384518 207916
rect 384574 207860 384642 207916
rect 384698 207860 384766 207916
rect 384822 207860 384890 207916
rect 384946 207860 385014 207916
rect 385070 207860 385138 207916
rect 385194 207860 385228 207916
rect 383988 207826 385228 207860
rect 403988 208412 405228 208446
rect 403988 208356 404022 208412
rect 404078 208356 404146 208412
rect 404202 208356 404270 208412
rect 404326 208356 404394 208412
rect 404450 208356 404518 208412
rect 404574 208356 404642 208412
rect 404698 208356 404766 208412
rect 404822 208356 404890 208412
rect 404946 208356 405014 208412
rect 405070 208356 405138 208412
rect 405194 208356 405228 208412
rect 403988 208288 405228 208356
rect 403988 208232 404022 208288
rect 404078 208232 404146 208288
rect 404202 208232 404270 208288
rect 404326 208232 404394 208288
rect 404450 208232 404518 208288
rect 404574 208232 404642 208288
rect 404698 208232 404766 208288
rect 404822 208232 404890 208288
rect 404946 208232 405014 208288
rect 405070 208232 405138 208288
rect 405194 208232 405228 208288
rect 403988 208164 405228 208232
rect 403988 208108 404022 208164
rect 404078 208108 404146 208164
rect 404202 208108 404270 208164
rect 404326 208108 404394 208164
rect 404450 208108 404518 208164
rect 404574 208108 404642 208164
rect 404698 208108 404766 208164
rect 404822 208108 404890 208164
rect 404946 208108 405014 208164
rect 405070 208108 405138 208164
rect 405194 208108 405228 208164
rect 403988 208040 405228 208108
rect 403988 207984 404022 208040
rect 404078 207984 404146 208040
rect 404202 207984 404270 208040
rect 404326 207984 404394 208040
rect 404450 207984 404518 208040
rect 404574 207984 404642 208040
rect 404698 207984 404766 208040
rect 404822 207984 404890 208040
rect 404946 207984 405014 208040
rect 405070 207984 405138 208040
rect 405194 207984 405228 208040
rect 403988 207916 405228 207984
rect 403988 207860 404022 207916
rect 404078 207860 404146 207916
rect 404202 207860 404270 207916
rect 404326 207860 404394 207916
rect 404450 207860 404518 207916
rect 404574 207860 404642 207916
rect 404698 207860 404766 207916
rect 404822 207860 404890 207916
rect 404946 207860 405014 207916
rect 405070 207860 405138 207916
rect 405194 207860 405228 207916
rect 403988 207826 405228 207860
rect 423988 208412 425228 208446
rect 423988 208356 424022 208412
rect 424078 208356 424146 208412
rect 424202 208356 424270 208412
rect 424326 208356 424394 208412
rect 424450 208356 424518 208412
rect 424574 208356 424642 208412
rect 424698 208356 424766 208412
rect 424822 208356 424890 208412
rect 424946 208356 425014 208412
rect 425070 208356 425138 208412
rect 425194 208356 425228 208412
rect 423988 208288 425228 208356
rect 423988 208232 424022 208288
rect 424078 208232 424146 208288
rect 424202 208232 424270 208288
rect 424326 208232 424394 208288
rect 424450 208232 424518 208288
rect 424574 208232 424642 208288
rect 424698 208232 424766 208288
rect 424822 208232 424890 208288
rect 424946 208232 425014 208288
rect 425070 208232 425138 208288
rect 425194 208232 425228 208288
rect 423988 208164 425228 208232
rect 423988 208108 424022 208164
rect 424078 208108 424146 208164
rect 424202 208108 424270 208164
rect 424326 208108 424394 208164
rect 424450 208108 424518 208164
rect 424574 208108 424642 208164
rect 424698 208108 424766 208164
rect 424822 208108 424890 208164
rect 424946 208108 425014 208164
rect 425070 208108 425138 208164
rect 425194 208108 425228 208164
rect 423988 208040 425228 208108
rect 423988 207984 424022 208040
rect 424078 207984 424146 208040
rect 424202 207984 424270 208040
rect 424326 207984 424394 208040
rect 424450 207984 424518 208040
rect 424574 207984 424642 208040
rect 424698 207984 424766 208040
rect 424822 207984 424890 208040
rect 424946 207984 425014 208040
rect 425070 207984 425138 208040
rect 425194 207984 425228 208040
rect 423988 207916 425228 207984
rect 423988 207860 424022 207916
rect 424078 207860 424146 207916
rect 424202 207860 424270 207916
rect 424326 207860 424394 207916
rect 424450 207860 424518 207916
rect 424574 207860 424642 207916
rect 424698 207860 424766 207916
rect 424822 207860 424890 207916
rect 424946 207860 425014 207916
rect 425070 207860 425138 207916
rect 425194 207860 425228 207916
rect 423988 207826 425228 207860
rect 443988 208412 445228 208446
rect 443988 208356 444022 208412
rect 444078 208356 444146 208412
rect 444202 208356 444270 208412
rect 444326 208356 444394 208412
rect 444450 208356 444518 208412
rect 444574 208356 444642 208412
rect 444698 208356 444766 208412
rect 444822 208356 444890 208412
rect 444946 208356 445014 208412
rect 445070 208356 445138 208412
rect 445194 208356 445228 208412
rect 443988 208288 445228 208356
rect 443988 208232 444022 208288
rect 444078 208232 444146 208288
rect 444202 208232 444270 208288
rect 444326 208232 444394 208288
rect 444450 208232 444518 208288
rect 444574 208232 444642 208288
rect 444698 208232 444766 208288
rect 444822 208232 444890 208288
rect 444946 208232 445014 208288
rect 445070 208232 445138 208288
rect 445194 208232 445228 208288
rect 443988 208164 445228 208232
rect 443988 208108 444022 208164
rect 444078 208108 444146 208164
rect 444202 208108 444270 208164
rect 444326 208108 444394 208164
rect 444450 208108 444518 208164
rect 444574 208108 444642 208164
rect 444698 208108 444766 208164
rect 444822 208108 444890 208164
rect 444946 208108 445014 208164
rect 445070 208108 445138 208164
rect 445194 208108 445228 208164
rect 443988 208040 445228 208108
rect 443988 207984 444022 208040
rect 444078 207984 444146 208040
rect 444202 207984 444270 208040
rect 444326 207984 444394 208040
rect 444450 207984 444518 208040
rect 444574 207984 444642 208040
rect 444698 207984 444766 208040
rect 444822 207984 444890 208040
rect 444946 207984 445014 208040
rect 445070 207984 445138 208040
rect 445194 207984 445228 208040
rect 443988 207916 445228 207984
rect 443988 207860 444022 207916
rect 444078 207860 444146 207916
rect 444202 207860 444270 207916
rect 444326 207860 444394 207916
rect 444450 207860 444518 207916
rect 444574 207860 444642 207916
rect 444698 207860 444766 207916
rect 444822 207860 444890 207916
rect 444946 207860 445014 207916
rect 445070 207860 445138 207916
rect 445194 207860 445228 207916
rect 443988 207826 445228 207860
rect 463988 208412 465228 208446
rect 463988 208356 464022 208412
rect 464078 208356 464146 208412
rect 464202 208356 464270 208412
rect 464326 208356 464394 208412
rect 464450 208356 464518 208412
rect 464574 208356 464642 208412
rect 464698 208356 464766 208412
rect 464822 208356 464890 208412
rect 464946 208356 465014 208412
rect 465070 208356 465138 208412
rect 465194 208356 465228 208412
rect 463988 208288 465228 208356
rect 463988 208232 464022 208288
rect 464078 208232 464146 208288
rect 464202 208232 464270 208288
rect 464326 208232 464394 208288
rect 464450 208232 464518 208288
rect 464574 208232 464642 208288
rect 464698 208232 464766 208288
rect 464822 208232 464890 208288
rect 464946 208232 465014 208288
rect 465070 208232 465138 208288
rect 465194 208232 465228 208288
rect 463988 208164 465228 208232
rect 463988 208108 464022 208164
rect 464078 208108 464146 208164
rect 464202 208108 464270 208164
rect 464326 208108 464394 208164
rect 464450 208108 464518 208164
rect 464574 208108 464642 208164
rect 464698 208108 464766 208164
rect 464822 208108 464890 208164
rect 464946 208108 465014 208164
rect 465070 208108 465138 208164
rect 465194 208108 465228 208164
rect 463988 208040 465228 208108
rect 463988 207984 464022 208040
rect 464078 207984 464146 208040
rect 464202 207984 464270 208040
rect 464326 207984 464394 208040
rect 464450 207984 464518 208040
rect 464574 207984 464642 208040
rect 464698 207984 464766 208040
rect 464822 207984 464890 208040
rect 464946 207984 465014 208040
rect 465070 207984 465138 208040
rect 465194 207984 465228 208040
rect 463988 207916 465228 207984
rect 463988 207860 464022 207916
rect 464078 207860 464146 207916
rect 464202 207860 464270 207916
rect 464326 207860 464394 207916
rect 464450 207860 464518 207916
rect 464574 207860 464642 207916
rect 464698 207860 464766 207916
rect 464822 207860 464890 207916
rect 464946 207860 465014 207916
rect 465070 207860 465138 207916
rect 465194 207860 465228 207916
rect 463988 207826 465228 207860
rect 483988 208412 485228 208446
rect 483988 208356 484022 208412
rect 484078 208356 484146 208412
rect 484202 208356 484270 208412
rect 484326 208356 484394 208412
rect 484450 208356 484518 208412
rect 484574 208356 484642 208412
rect 484698 208356 484766 208412
rect 484822 208356 484890 208412
rect 484946 208356 485014 208412
rect 485070 208356 485138 208412
rect 485194 208356 485228 208412
rect 483988 208288 485228 208356
rect 483988 208232 484022 208288
rect 484078 208232 484146 208288
rect 484202 208232 484270 208288
rect 484326 208232 484394 208288
rect 484450 208232 484518 208288
rect 484574 208232 484642 208288
rect 484698 208232 484766 208288
rect 484822 208232 484890 208288
rect 484946 208232 485014 208288
rect 485070 208232 485138 208288
rect 485194 208232 485228 208288
rect 483988 208164 485228 208232
rect 483988 208108 484022 208164
rect 484078 208108 484146 208164
rect 484202 208108 484270 208164
rect 484326 208108 484394 208164
rect 484450 208108 484518 208164
rect 484574 208108 484642 208164
rect 484698 208108 484766 208164
rect 484822 208108 484890 208164
rect 484946 208108 485014 208164
rect 485070 208108 485138 208164
rect 485194 208108 485228 208164
rect 483988 208040 485228 208108
rect 483988 207984 484022 208040
rect 484078 207984 484146 208040
rect 484202 207984 484270 208040
rect 484326 207984 484394 208040
rect 484450 207984 484518 208040
rect 484574 207984 484642 208040
rect 484698 207984 484766 208040
rect 484822 207984 484890 208040
rect 484946 207984 485014 208040
rect 485070 207984 485138 208040
rect 485194 207984 485228 208040
rect 483988 207916 485228 207984
rect 483988 207860 484022 207916
rect 484078 207860 484146 207916
rect 484202 207860 484270 207916
rect 484326 207860 484394 207916
rect 484450 207860 484518 207916
rect 484574 207860 484642 207916
rect 484698 207860 484766 207916
rect 484822 207860 484890 207916
rect 484946 207860 485014 207916
rect 485070 207860 485138 207916
rect 485194 207860 485228 207916
rect 483988 207826 485228 207860
rect 503988 208412 505228 208446
rect 503988 208356 504022 208412
rect 504078 208356 504146 208412
rect 504202 208356 504270 208412
rect 504326 208356 504394 208412
rect 504450 208356 504518 208412
rect 504574 208356 504642 208412
rect 504698 208356 504766 208412
rect 504822 208356 504890 208412
rect 504946 208356 505014 208412
rect 505070 208356 505138 208412
rect 505194 208356 505228 208412
rect 503988 208288 505228 208356
rect 503988 208232 504022 208288
rect 504078 208232 504146 208288
rect 504202 208232 504270 208288
rect 504326 208232 504394 208288
rect 504450 208232 504518 208288
rect 504574 208232 504642 208288
rect 504698 208232 504766 208288
rect 504822 208232 504890 208288
rect 504946 208232 505014 208288
rect 505070 208232 505138 208288
rect 505194 208232 505228 208288
rect 503988 208164 505228 208232
rect 503988 208108 504022 208164
rect 504078 208108 504146 208164
rect 504202 208108 504270 208164
rect 504326 208108 504394 208164
rect 504450 208108 504518 208164
rect 504574 208108 504642 208164
rect 504698 208108 504766 208164
rect 504822 208108 504890 208164
rect 504946 208108 505014 208164
rect 505070 208108 505138 208164
rect 505194 208108 505228 208164
rect 503988 208040 505228 208108
rect 503988 207984 504022 208040
rect 504078 207984 504146 208040
rect 504202 207984 504270 208040
rect 504326 207984 504394 208040
rect 504450 207984 504518 208040
rect 504574 207984 504642 208040
rect 504698 207984 504766 208040
rect 504822 207984 504890 208040
rect 504946 207984 505014 208040
rect 505070 207984 505138 208040
rect 505194 207984 505228 208040
rect 503988 207916 505228 207984
rect 503988 207860 504022 207916
rect 504078 207860 504146 207916
rect 504202 207860 504270 207916
rect 504326 207860 504394 207916
rect 504450 207860 504518 207916
rect 504574 207860 504642 207916
rect 504698 207860 504766 207916
rect 504822 207860 504890 207916
rect 504946 207860 505014 207916
rect 505070 207860 505138 207916
rect 505194 207860 505228 207916
rect 503988 207826 505228 207860
rect 523988 208412 525228 208446
rect 523988 208356 524022 208412
rect 524078 208356 524146 208412
rect 524202 208356 524270 208412
rect 524326 208356 524394 208412
rect 524450 208356 524518 208412
rect 524574 208356 524642 208412
rect 524698 208356 524766 208412
rect 524822 208356 524890 208412
rect 524946 208356 525014 208412
rect 525070 208356 525138 208412
rect 525194 208356 525228 208412
rect 523988 208288 525228 208356
rect 523988 208232 524022 208288
rect 524078 208232 524146 208288
rect 524202 208232 524270 208288
rect 524326 208232 524394 208288
rect 524450 208232 524518 208288
rect 524574 208232 524642 208288
rect 524698 208232 524766 208288
rect 524822 208232 524890 208288
rect 524946 208232 525014 208288
rect 525070 208232 525138 208288
rect 525194 208232 525228 208288
rect 523988 208164 525228 208232
rect 523988 208108 524022 208164
rect 524078 208108 524146 208164
rect 524202 208108 524270 208164
rect 524326 208108 524394 208164
rect 524450 208108 524518 208164
rect 524574 208108 524642 208164
rect 524698 208108 524766 208164
rect 524822 208108 524890 208164
rect 524946 208108 525014 208164
rect 525070 208108 525138 208164
rect 525194 208108 525228 208164
rect 523988 208040 525228 208108
rect 523988 207984 524022 208040
rect 524078 207984 524146 208040
rect 524202 207984 524270 208040
rect 524326 207984 524394 208040
rect 524450 207984 524518 208040
rect 524574 207984 524642 208040
rect 524698 207984 524766 208040
rect 524822 207984 524890 208040
rect 524946 207984 525014 208040
rect 525070 207984 525138 208040
rect 525194 207984 525228 208040
rect 523988 207916 525228 207984
rect 523988 207860 524022 207916
rect 524078 207860 524146 207916
rect 524202 207860 524270 207916
rect 524326 207860 524394 207916
rect 524450 207860 524518 207916
rect 524574 207860 524642 207916
rect 524698 207860 524766 207916
rect 524822 207860 524890 207916
rect 524946 207860 525014 207916
rect 525070 207860 525138 207916
rect 525194 207860 525228 207916
rect 523988 207826 525228 207860
rect 543988 208412 545228 208446
rect 543988 208356 544022 208412
rect 544078 208356 544146 208412
rect 544202 208356 544270 208412
rect 544326 208356 544394 208412
rect 544450 208356 544518 208412
rect 544574 208356 544642 208412
rect 544698 208356 544766 208412
rect 544822 208356 544890 208412
rect 544946 208356 545014 208412
rect 545070 208356 545138 208412
rect 545194 208356 545228 208412
rect 543988 208288 545228 208356
rect 543988 208232 544022 208288
rect 544078 208232 544146 208288
rect 544202 208232 544270 208288
rect 544326 208232 544394 208288
rect 544450 208232 544518 208288
rect 544574 208232 544642 208288
rect 544698 208232 544766 208288
rect 544822 208232 544890 208288
rect 544946 208232 545014 208288
rect 545070 208232 545138 208288
rect 545194 208232 545228 208288
rect 543988 208164 545228 208232
rect 543988 208108 544022 208164
rect 544078 208108 544146 208164
rect 544202 208108 544270 208164
rect 544326 208108 544394 208164
rect 544450 208108 544518 208164
rect 544574 208108 544642 208164
rect 544698 208108 544766 208164
rect 544822 208108 544890 208164
rect 544946 208108 545014 208164
rect 545070 208108 545138 208164
rect 545194 208108 545228 208164
rect 543988 208040 545228 208108
rect 543988 207984 544022 208040
rect 544078 207984 544146 208040
rect 544202 207984 544270 208040
rect 544326 207984 544394 208040
rect 544450 207984 544518 208040
rect 544574 207984 544642 208040
rect 544698 207984 544766 208040
rect 544822 207984 544890 208040
rect 544946 207984 545014 208040
rect 545070 207984 545138 208040
rect 545194 207984 545228 208040
rect 543988 207916 545228 207984
rect 543988 207860 544022 207916
rect 544078 207860 544146 207916
rect 544202 207860 544270 207916
rect 544326 207860 544394 207916
rect 544450 207860 544518 207916
rect 544574 207860 544642 207916
rect 544698 207860 544766 207916
rect 544822 207860 544890 207916
rect 544946 207860 545014 207916
rect 545070 207860 545138 207916
rect 545194 207860 545228 207916
rect 543988 207826 545228 207860
rect 353988 202412 355228 202446
rect 353988 202356 354022 202412
rect 354078 202356 354146 202412
rect 354202 202356 354270 202412
rect 354326 202356 354394 202412
rect 354450 202356 354518 202412
rect 354574 202356 354642 202412
rect 354698 202356 354766 202412
rect 354822 202356 354890 202412
rect 354946 202356 355014 202412
rect 355070 202356 355138 202412
rect 355194 202356 355228 202412
rect 353988 202288 355228 202356
rect 353988 202232 354022 202288
rect 354078 202232 354146 202288
rect 354202 202232 354270 202288
rect 354326 202232 354394 202288
rect 354450 202232 354518 202288
rect 354574 202232 354642 202288
rect 354698 202232 354766 202288
rect 354822 202232 354890 202288
rect 354946 202232 355014 202288
rect 355070 202232 355138 202288
rect 355194 202232 355228 202288
rect 353988 202164 355228 202232
rect 353988 202108 354022 202164
rect 354078 202108 354146 202164
rect 354202 202108 354270 202164
rect 354326 202108 354394 202164
rect 354450 202108 354518 202164
rect 354574 202108 354642 202164
rect 354698 202108 354766 202164
rect 354822 202108 354890 202164
rect 354946 202108 355014 202164
rect 355070 202108 355138 202164
rect 355194 202108 355228 202164
rect 353988 202040 355228 202108
rect 353988 201984 354022 202040
rect 354078 201984 354146 202040
rect 354202 201984 354270 202040
rect 354326 201984 354394 202040
rect 354450 201984 354518 202040
rect 354574 201984 354642 202040
rect 354698 201984 354766 202040
rect 354822 201984 354890 202040
rect 354946 201984 355014 202040
rect 355070 201984 355138 202040
rect 355194 201984 355228 202040
rect 353988 201916 355228 201984
rect 353988 201860 354022 201916
rect 354078 201860 354146 201916
rect 354202 201860 354270 201916
rect 354326 201860 354394 201916
rect 354450 201860 354518 201916
rect 354574 201860 354642 201916
rect 354698 201860 354766 201916
rect 354822 201860 354890 201916
rect 354946 201860 355014 201916
rect 355070 201860 355138 201916
rect 355194 201860 355228 201916
rect 353988 201826 355228 201860
rect 373988 202412 375228 202446
rect 373988 202356 374022 202412
rect 374078 202356 374146 202412
rect 374202 202356 374270 202412
rect 374326 202356 374394 202412
rect 374450 202356 374518 202412
rect 374574 202356 374642 202412
rect 374698 202356 374766 202412
rect 374822 202356 374890 202412
rect 374946 202356 375014 202412
rect 375070 202356 375138 202412
rect 375194 202356 375228 202412
rect 373988 202288 375228 202356
rect 373988 202232 374022 202288
rect 374078 202232 374146 202288
rect 374202 202232 374270 202288
rect 374326 202232 374394 202288
rect 374450 202232 374518 202288
rect 374574 202232 374642 202288
rect 374698 202232 374766 202288
rect 374822 202232 374890 202288
rect 374946 202232 375014 202288
rect 375070 202232 375138 202288
rect 375194 202232 375228 202288
rect 373988 202164 375228 202232
rect 373988 202108 374022 202164
rect 374078 202108 374146 202164
rect 374202 202108 374270 202164
rect 374326 202108 374394 202164
rect 374450 202108 374518 202164
rect 374574 202108 374642 202164
rect 374698 202108 374766 202164
rect 374822 202108 374890 202164
rect 374946 202108 375014 202164
rect 375070 202108 375138 202164
rect 375194 202108 375228 202164
rect 373988 202040 375228 202108
rect 373988 201984 374022 202040
rect 374078 201984 374146 202040
rect 374202 201984 374270 202040
rect 374326 201984 374394 202040
rect 374450 201984 374518 202040
rect 374574 201984 374642 202040
rect 374698 201984 374766 202040
rect 374822 201984 374890 202040
rect 374946 201984 375014 202040
rect 375070 201984 375138 202040
rect 375194 201984 375228 202040
rect 373988 201916 375228 201984
rect 373988 201860 374022 201916
rect 374078 201860 374146 201916
rect 374202 201860 374270 201916
rect 374326 201860 374394 201916
rect 374450 201860 374518 201916
rect 374574 201860 374642 201916
rect 374698 201860 374766 201916
rect 374822 201860 374890 201916
rect 374946 201860 375014 201916
rect 375070 201860 375138 201916
rect 375194 201860 375228 201916
rect 373988 201826 375228 201860
rect 393988 202412 395228 202446
rect 393988 202356 394022 202412
rect 394078 202356 394146 202412
rect 394202 202356 394270 202412
rect 394326 202356 394394 202412
rect 394450 202356 394518 202412
rect 394574 202356 394642 202412
rect 394698 202356 394766 202412
rect 394822 202356 394890 202412
rect 394946 202356 395014 202412
rect 395070 202356 395138 202412
rect 395194 202356 395228 202412
rect 393988 202288 395228 202356
rect 393988 202232 394022 202288
rect 394078 202232 394146 202288
rect 394202 202232 394270 202288
rect 394326 202232 394394 202288
rect 394450 202232 394518 202288
rect 394574 202232 394642 202288
rect 394698 202232 394766 202288
rect 394822 202232 394890 202288
rect 394946 202232 395014 202288
rect 395070 202232 395138 202288
rect 395194 202232 395228 202288
rect 393988 202164 395228 202232
rect 393988 202108 394022 202164
rect 394078 202108 394146 202164
rect 394202 202108 394270 202164
rect 394326 202108 394394 202164
rect 394450 202108 394518 202164
rect 394574 202108 394642 202164
rect 394698 202108 394766 202164
rect 394822 202108 394890 202164
rect 394946 202108 395014 202164
rect 395070 202108 395138 202164
rect 395194 202108 395228 202164
rect 393988 202040 395228 202108
rect 393988 201984 394022 202040
rect 394078 201984 394146 202040
rect 394202 201984 394270 202040
rect 394326 201984 394394 202040
rect 394450 201984 394518 202040
rect 394574 201984 394642 202040
rect 394698 201984 394766 202040
rect 394822 201984 394890 202040
rect 394946 201984 395014 202040
rect 395070 201984 395138 202040
rect 395194 201984 395228 202040
rect 393988 201916 395228 201984
rect 393988 201860 394022 201916
rect 394078 201860 394146 201916
rect 394202 201860 394270 201916
rect 394326 201860 394394 201916
rect 394450 201860 394518 201916
rect 394574 201860 394642 201916
rect 394698 201860 394766 201916
rect 394822 201860 394890 201916
rect 394946 201860 395014 201916
rect 395070 201860 395138 201916
rect 395194 201860 395228 201916
rect 393988 201826 395228 201860
rect 413988 202412 415228 202446
rect 413988 202356 414022 202412
rect 414078 202356 414146 202412
rect 414202 202356 414270 202412
rect 414326 202356 414394 202412
rect 414450 202356 414518 202412
rect 414574 202356 414642 202412
rect 414698 202356 414766 202412
rect 414822 202356 414890 202412
rect 414946 202356 415014 202412
rect 415070 202356 415138 202412
rect 415194 202356 415228 202412
rect 413988 202288 415228 202356
rect 413988 202232 414022 202288
rect 414078 202232 414146 202288
rect 414202 202232 414270 202288
rect 414326 202232 414394 202288
rect 414450 202232 414518 202288
rect 414574 202232 414642 202288
rect 414698 202232 414766 202288
rect 414822 202232 414890 202288
rect 414946 202232 415014 202288
rect 415070 202232 415138 202288
rect 415194 202232 415228 202288
rect 413988 202164 415228 202232
rect 413988 202108 414022 202164
rect 414078 202108 414146 202164
rect 414202 202108 414270 202164
rect 414326 202108 414394 202164
rect 414450 202108 414518 202164
rect 414574 202108 414642 202164
rect 414698 202108 414766 202164
rect 414822 202108 414890 202164
rect 414946 202108 415014 202164
rect 415070 202108 415138 202164
rect 415194 202108 415228 202164
rect 413988 202040 415228 202108
rect 413988 201984 414022 202040
rect 414078 201984 414146 202040
rect 414202 201984 414270 202040
rect 414326 201984 414394 202040
rect 414450 201984 414518 202040
rect 414574 201984 414642 202040
rect 414698 201984 414766 202040
rect 414822 201984 414890 202040
rect 414946 201984 415014 202040
rect 415070 201984 415138 202040
rect 415194 201984 415228 202040
rect 413988 201916 415228 201984
rect 413988 201860 414022 201916
rect 414078 201860 414146 201916
rect 414202 201860 414270 201916
rect 414326 201860 414394 201916
rect 414450 201860 414518 201916
rect 414574 201860 414642 201916
rect 414698 201860 414766 201916
rect 414822 201860 414890 201916
rect 414946 201860 415014 201916
rect 415070 201860 415138 201916
rect 415194 201860 415228 201916
rect 413988 201826 415228 201860
rect 433988 202412 435228 202446
rect 433988 202356 434022 202412
rect 434078 202356 434146 202412
rect 434202 202356 434270 202412
rect 434326 202356 434394 202412
rect 434450 202356 434518 202412
rect 434574 202356 434642 202412
rect 434698 202356 434766 202412
rect 434822 202356 434890 202412
rect 434946 202356 435014 202412
rect 435070 202356 435138 202412
rect 435194 202356 435228 202412
rect 433988 202288 435228 202356
rect 433988 202232 434022 202288
rect 434078 202232 434146 202288
rect 434202 202232 434270 202288
rect 434326 202232 434394 202288
rect 434450 202232 434518 202288
rect 434574 202232 434642 202288
rect 434698 202232 434766 202288
rect 434822 202232 434890 202288
rect 434946 202232 435014 202288
rect 435070 202232 435138 202288
rect 435194 202232 435228 202288
rect 433988 202164 435228 202232
rect 433988 202108 434022 202164
rect 434078 202108 434146 202164
rect 434202 202108 434270 202164
rect 434326 202108 434394 202164
rect 434450 202108 434518 202164
rect 434574 202108 434642 202164
rect 434698 202108 434766 202164
rect 434822 202108 434890 202164
rect 434946 202108 435014 202164
rect 435070 202108 435138 202164
rect 435194 202108 435228 202164
rect 433988 202040 435228 202108
rect 433988 201984 434022 202040
rect 434078 201984 434146 202040
rect 434202 201984 434270 202040
rect 434326 201984 434394 202040
rect 434450 201984 434518 202040
rect 434574 201984 434642 202040
rect 434698 201984 434766 202040
rect 434822 201984 434890 202040
rect 434946 201984 435014 202040
rect 435070 201984 435138 202040
rect 435194 201984 435228 202040
rect 433988 201916 435228 201984
rect 433988 201860 434022 201916
rect 434078 201860 434146 201916
rect 434202 201860 434270 201916
rect 434326 201860 434394 201916
rect 434450 201860 434518 201916
rect 434574 201860 434642 201916
rect 434698 201860 434766 201916
rect 434822 201860 434890 201916
rect 434946 201860 435014 201916
rect 435070 201860 435138 201916
rect 435194 201860 435228 201916
rect 433988 201826 435228 201860
rect 453988 202412 455228 202446
rect 453988 202356 454022 202412
rect 454078 202356 454146 202412
rect 454202 202356 454270 202412
rect 454326 202356 454394 202412
rect 454450 202356 454518 202412
rect 454574 202356 454642 202412
rect 454698 202356 454766 202412
rect 454822 202356 454890 202412
rect 454946 202356 455014 202412
rect 455070 202356 455138 202412
rect 455194 202356 455228 202412
rect 453988 202288 455228 202356
rect 453988 202232 454022 202288
rect 454078 202232 454146 202288
rect 454202 202232 454270 202288
rect 454326 202232 454394 202288
rect 454450 202232 454518 202288
rect 454574 202232 454642 202288
rect 454698 202232 454766 202288
rect 454822 202232 454890 202288
rect 454946 202232 455014 202288
rect 455070 202232 455138 202288
rect 455194 202232 455228 202288
rect 453988 202164 455228 202232
rect 453988 202108 454022 202164
rect 454078 202108 454146 202164
rect 454202 202108 454270 202164
rect 454326 202108 454394 202164
rect 454450 202108 454518 202164
rect 454574 202108 454642 202164
rect 454698 202108 454766 202164
rect 454822 202108 454890 202164
rect 454946 202108 455014 202164
rect 455070 202108 455138 202164
rect 455194 202108 455228 202164
rect 453988 202040 455228 202108
rect 453988 201984 454022 202040
rect 454078 201984 454146 202040
rect 454202 201984 454270 202040
rect 454326 201984 454394 202040
rect 454450 201984 454518 202040
rect 454574 201984 454642 202040
rect 454698 201984 454766 202040
rect 454822 201984 454890 202040
rect 454946 201984 455014 202040
rect 455070 201984 455138 202040
rect 455194 201984 455228 202040
rect 453988 201916 455228 201984
rect 453988 201860 454022 201916
rect 454078 201860 454146 201916
rect 454202 201860 454270 201916
rect 454326 201860 454394 201916
rect 454450 201860 454518 201916
rect 454574 201860 454642 201916
rect 454698 201860 454766 201916
rect 454822 201860 454890 201916
rect 454946 201860 455014 201916
rect 455070 201860 455138 201916
rect 455194 201860 455228 201916
rect 453988 201826 455228 201860
rect 473988 202412 475228 202446
rect 473988 202356 474022 202412
rect 474078 202356 474146 202412
rect 474202 202356 474270 202412
rect 474326 202356 474394 202412
rect 474450 202356 474518 202412
rect 474574 202356 474642 202412
rect 474698 202356 474766 202412
rect 474822 202356 474890 202412
rect 474946 202356 475014 202412
rect 475070 202356 475138 202412
rect 475194 202356 475228 202412
rect 473988 202288 475228 202356
rect 473988 202232 474022 202288
rect 474078 202232 474146 202288
rect 474202 202232 474270 202288
rect 474326 202232 474394 202288
rect 474450 202232 474518 202288
rect 474574 202232 474642 202288
rect 474698 202232 474766 202288
rect 474822 202232 474890 202288
rect 474946 202232 475014 202288
rect 475070 202232 475138 202288
rect 475194 202232 475228 202288
rect 473988 202164 475228 202232
rect 473988 202108 474022 202164
rect 474078 202108 474146 202164
rect 474202 202108 474270 202164
rect 474326 202108 474394 202164
rect 474450 202108 474518 202164
rect 474574 202108 474642 202164
rect 474698 202108 474766 202164
rect 474822 202108 474890 202164
rect 474946 202108 475014 202164
rect 475070 202108 475138 202164
rect 475194 202108 475228 202164
rect 473988 202040 475228 202108
rect 473988 201984 474022 202040
rect 474078 201984 474146 202040
rect 474202 201984 474270 202040
rect 474326 201984 474394 202040
rect 474450 201984 474518 202040
rect 474574 201984 474642 202040
rect 474698 201984 474766 202040
rect 474822 201984 474890 202040
rect 474946 201984 475014 202040
rect 475070 201984 475138 202040
rect 475194 201984 475228 202040
rect 473988 201916 475228 201984
rect 473988 201860 474022 201916
rect 474078 201860 474146 201916
rect 474202 201860 474270 201916
rect 474326 201860 474394 201916
rect 474450 201860 474518 201916
rect 474574 201860 474642 201916
rect 474698 201860 474766 201916
rect 474822 201860 474890 201916
rect 474946 201860 475014 201916
rect 475070 201860 475138 201916
rect 475194 201860 475228 201916
rect 473988 201826 475228 201860
rect 493988 202412 495228 202446
rect 493988 202356 494022 202412
rect 494078 202356 494146 202412
rect 494202 202356 494270 202412
rect 494326 202356 494394 202412
rect 494450 202356 494518 202412
rect 494574 202356 494642 202412
rect 494698 202356 494766 202412
rect 494822 202356 494890 202412
rect 494946 202356 495014 202412
rect 495070 202356 495138 202412
rect 495194 202356 495228 202412
rect 493988 202288 495228 202356
rect 493988 202232 494022 202288
rect 494078 202232 494146 202288
rect 494202 202232 494270 202288
rect 494326 202232 494394 202288
rect 494450 202232 494518 202288
rect 494574 202232 494642 202288
rect 494698 202232 494766 202288
rect 494822 202232 494890 202288
rect 494946 202232 495014 202288
rect 495070 202232 495138 202288
rect 495194 202232 495228 202288
rect 493988 202164 495228 202232
rect 493988 202108 494022 202164
rect 494078 202108 494146 202164
rect 494202 202108 494270 202164
rect 494326 202108 494394 202164
rect 494450 202108 494518 202164
rect 494574 202108 494642 202164
rect 494698 202108 494766 202164
rect 494822 202108 494890 202164
rect 494946 202108 495014 202164
rect 495070 202108 495138 202164
rect 495194 202108 495228 202164
rect 493988 202040 495228 202108
rect 493988 201984 494022 202040
rect 494078 201984 494146 202040
rect 494202 201984 494270 202040
rect 494326 201984 494394 202040
rect 494450 201984 494518 202040
rect 494574 201984 494642 202040
rect 494698 201984 494766 202040
rect 494822 201984 494890 202040
rect 494946 201984 495014 202040
rect 495070 201984 495138 202040
rect 495194 201984 495228 202040
rect 493988 201916 495228 201984
rect 493988 201860 494022 201916
rect 494078 201860 494146 201916
rect 494202 201860 494270 201916
rect 494326 201860 494394 201916
rect 494450 201860 494518 201916
rect 494574 201860 494642 201916
rect 494698 201860 494766 201916
rect 494822 201860 494890 201916
rect 494946 201860 495014 201916
rect 495070 201860 495138 201916
rect 495194 201860 495228 201916
rect 493988 201826 495228 201860
rect 513988 202412 515228 202446
rect 513988 202356 514022 202412
rect 514078 202356 514146 202412
rect 514202 202356 514270 202412
rect 514326 202356 514394 202412
rect 514450 202356 514518 202412
rect 514574 202356 514642 202412
rect 514698 202356 514766 202412
rect 514822 202356 514890 202412
rect 514946 202356 515014 202412
rect 515070 202356 515138 202412
rect 515194 202356 515228 202412
rect 513988 202288 515228 202356
rect 513988 202232 514022 202288
rect 514078 202232 514146 202288
rect 514202 202232 514270 202288
rect 514326 202232 514394 202288
rect 514450 202232 514518 202288
rect 514574 202232 514642 202288
rect 514698 202232 514766 202288
rect 514822 202232 514890 202288
rect 514946 202232 515014 202288
rect 515070 202232 515138 202288
rect 515194 202232 515228 202288
rect 513988 202164 515228 202232
rect 513988 202108 514022 202164
rect 514078 202108 514146 202164
rect 514202 202108 514270 202164
rect 514326 202108 514394 202164
rect 514450 202108 514518 202164
rect 514574 202108 514642 202164
rect 514698 202108 514766 202164
rect 514822 202108 514890 202164
rect 514946 202108 515014 202164
rect 515070 202108 515138 202164
rect 515194 202108 515228 202164
rect 513988 202040 515228 202108
rect 513988 201984 514022 202040
rect 514078 201984 514146 202040
rect 514202 201984 514270 202040
rect 514326 201984 514394 202040
rect 514450 201984 514518 202040
rect 514574 201984 514642 202040
rect 514698 201984 514766 202040
rect 514822 201984 514890 202040
rect 514946 201984 515014 202040
rect 515070 201984 515138 202040
rect 515194 201984 515228 202040
rect 513988 201916 515228 201984
rect 513988 201860 514022 201916
rect 514078 201860 514146 201916
rect 514202 201860 514270 201916
rect 514326 201860 514394 201916
rect 514450 201860 514518 201916
rect 514574 201860 514642 201916
rect 514698 201860 514766 201916
rect 514822 201860 514890 201916
rect 514946 201860 515014 201916
rect 515070 201860 515138 201916
rect 515194 201860 515228 201916
rect 513988 201826 515228 201860
rect 533988 202412 535228 202446
rect 533988 202356 534022 202412
rect 534078 202356 534146 202412
rect 534202 202356 534270 202412
rect 534326 202356 534394 202412
rect 534450 202356 534518 202412
rect 534574 202356 534642 202412
rect 534698 202356 534766 202412
rect 534822 202356 534890 202412
rect 534946 202356 535014 202412
rect 535070 202356 535138 202412
rect 535194 202356 535228 202412
rect 533988 202288 535228 202356
rect 533988 202232 534022 202288
rect 534078 202232 534146 202288
rect 534202 202232 534270 202288
rect 534326 202232 534394 202288
rect 534450 202232 534518 202288
rect 534574 202232 534642 202288
rect 534698 202232 534766 202288
rect 534822 202232 534890 202288
rect 534946 202232 535014 202288
rect 535070 202232 535138 202288
rect 535194 202232 535228 202288
rect 533988 202164 535228 202232
rect 533988 202108 534022 202164
rect 534078 202108 534146 202164
rect 534202 202108 534270 202164
rect 534326 202108 534394 202164
rect 534450 202108 534518 202164
rect 534574 202108 534642 202164
rect 534698 202108 534766 202164
rect 534822 202108 534890 202164
rect 534946 202108 535014 202164
rect 535070 202108 535138 202164
rect 535194 202108 535228 202164
rect 533988 202040 535228 202108
rect 533988 201984 534022 202040
rect 534078 201984 534146 202040
rect 534202 201984 534270 202040
rect 534326 201984 534394 202040
rect 534450 201984 534518 202040
rect 534574 201984 534642 202040
rect 534698 201984 534766 202040
rect 534822 201984 534890 202040
rect 534946 201984 535014 202040
rect 535070 201984 535138 202040
rect 535194 201984 535228 202040
rect 533988 201916 535228 201984
rect 533988 201860 534022 201916
rect 534078 201860 534146 201916
rect 534202 201860 534270 201916
rect 534326 201860 534394 201916
rect 534450 201860 534518 201916
rect 534574 201860 534642 201916
rect 534698 201860 534766 201916
rect 534822 201860 534890 201916
rect 534946 201860 535014 201916
rect 535070 201860 535138 201916
rect 535194 201860 535228 201916
rect 533988 201826 535228 201860
rect 348874 190294 348970 190350
rect 349026 190294 349094 190350
rect 349150 190294 349218 190350
rect 349274 190294 349342 190350
rect 349398 190294 349494 190350
rect 348874 190226 349494 190294
rect 348874 190170 348970 190226
rect 349026 190170 349094 190226
rect 349150 190170 349218 190226
rect 349274 190170 349342 190226
rect 349398 190170 349494 190226
rect 348874 190102 349494 190170
rect 348874 190046 348970 190102
rect 349026 190046 349094 190102
rect 349150 190046 349218 190102
rect 349274 190046 349342 190102
rect 349398 190046 349494 190102
rect 348874 189978 349494 190046
rect 348874 189922 348970 189978
rect 349026 189922 349094 189978
rect 349150 189922 349218 189978
rect 349274 189922 349342 189978
rect 349398 189922 349494 189978
rect 347676 183652 347732 183662
rect 347564 178276 347620 178286
rect 347452 172900 347508 172910
rect 345154 166294 345250 166350
rect 345306 166294 345374 166350
rect 345430 166294 345498 166350
rect 345554 166294 345622 166350
rect 345678 166294 345774 166350
rect 345154 166226 345774 166294
rect 345154 166170 345250 166226
rect 345306 166170 345374 166226
rect 345430 166170 345498 166226
rect 345554 166170 345622 166226
rect 345678 166170 345774 166226
rect 345154 166102 345774 166170
rect 345154 166046 345250 166102
rect 345306 166046 345374 166102
rect 345430 166046 345498 166102
rect 345554 166046 345622 166102
rect 345678 166046 345774 166102
rect 345154 165978 345774 166046
rect 345154 165922 345250 165978
rect 345306 165922 345374 165978
rect 345430 165922 345498 165978
rect 345554 165922 345622 165978
rect 345678 165922 345774 165978
rect 345154 148350 345774 165922
rect 345154 148294 345250 148350
rect 345306 148294 345374 148350
rect 345430 148294 345498 148350
rect 345554 148294 345622 148350
rect 345678 148294 345774 148350
rect 345154 148226 345774 148294
rect 345154 148170 345250 148226
rect 345306 148170 345374 148226
rect 345430 148170 345498 148226
rect 345554 148170 345622 148226
rect 345678 148170 345774 148226
rect 345154 148102 345774 148170
rect 345154 148046 345250 148102
rect 345306 148046 345374 148102
rect 345430 148046 345498 148102
rect 345554 148046 345622 148102
rect 345678 148046 345774 148102
rect 345154 147978 345774 148046
rect 345154 147922 345250 147978
rect 345306 147922 345374 147978
rect 345430 147922 345498 147978
rect 345554 147922 345622 147978
rect 345678 147922 345774 147978
rect 345154 130350 345774 147922
rect 345154 130294 345250 130350
rect 345306 130294 345374 130350
rect 345430 130294 345498 130350
rect 345554 130294 345622 130350
rect 345678 130294 345774 130350
rect 345154 130226 345774 130294
rect 345154 130170 345250 130226
rect 345306 130170 345374 130226
rect 345430 130170 345498 130226
rect 345554 130170 345622 130226
rect 345678 130170 345774 130226
rect 345154 130102 345774 130170
rect 345154 130046 345250 130102
rect 345306 130046 345374 130102
rect 345430 130046 345498 130102
rect 345554 130046 345622 130102
rect 345678 130046 345774 130102
rect 345154 129978 345774 130046
rect 345154 129922 345250 129978
rect 345306 129922 345374 129978
rect 345430 129922 345498 129978
rect 345554 129922 345622 129978
rect 345678 129922 345774 129978
rect 345154 112350 345774 129922
rect 345154 112294 345250 112350
rect 345306 112294 345374 112350
rect 345430 112294 345498 112350
rect 345554 112294 345622 112350
rect 345678 112294 345774 112350
rect 345154 112226 345774 112294
rect 345154 112170 345250 112226
rect 345306 112170 345374 112226
rect 345430 112170 345498 112226
rect 345554 112170 345622 112226
rect 345678 112170 345774 112226
rect 345154 112102 345774 112170
rect 345154 112046 345250 112102
rect 345306 112046 345374 112102
rect 345430 112046 345498 112102
rect 345554 112046 345622 112102
rect 345678 112046 345774 112102
rect 345154 111978 345774 112046
rect 345154 111922 345250 111978
rect 345306 111922 345374 111978
rect 345430 111922 345498 111978
rect 345554 111922 345622 111978
rect 345678 111922 345774 111978
rect 345154 94350 345774 111922
rect 346892 167524 346948 167534
rect 345154 94294 345250 94350
rect 345306 94294 345374 94350
rect 345430 94294 345498 94350
rect 345554 94294 345622 94350
rect 345678 94294 345774 94350
rect 345154 94226 345774 94294
rect 345154 94170 345250 94226
rect 345306 94170 345374 94226
rect 345430 94170 345498 94226
rect 345554 94170 345622 94226
rect 345678 94170 345774 94226
rect 345154 94102 345774 94170
rect 345154 94046 345250 94102
rect 345306 94046 345374 94102
rect 345430 94046 345498 94102
rect 345554 94046 345622 94102
rect 345678 94046 345774 94102
rect 345154 93978 345774 94046
rect 345154 93922 345250 93978
rect 345306 93922 345374 93978
rect 345430 93922 345498 93978
rect 345554 93922 345622 93978
rect 345678 93922 345774 93978
rect 345154 76350 345774 93922
rect 345154 76294 345250 76350
rect 345306 76294 345374 76350
rect 345430 76294 345498 76350
rect 345554 76294 345622 76350
rect 345678 76294 345774 76350
rect 345154 76226 345774 76294
rect 345154 76170 345250 76226
rect 345306 76170 345374 76226
rect 345430 76170 345498 76226
rect 345554 76170 345622 76226
rect 345678 76170 345774 76226
rect 345154 76102 345774 76170
rect 345154 76046 345250 76102
rect 345306 76046 345374 76102
rect 345430 76046 345498 76102
rect 345554 76046 345622 76102
rect 345678 76046 345774 76102
rect 345154 75978 345774 76046
rect 345154 75922 345250 75978
rect 345306 75922 345374 75978
rect 345430 75922 345498 75978
rect 345554 75922 345622 75978
rect 345678 75922 345774 75978
rect 345154 58350 345774 75922
rect 345154 58294 345250 58350
rect 345306 58294 345374 58350
rect 345430 58294 345498 58350
rect 345554 58294 345622 58350
rect 345678 58294 345774 58350
rect 345154 58226 345774 58294
rect 345154 58170 345250 58226
rect 345306 58170 345374 58226
rect 345430 58170 345498 58226
rect 345554 58170 345622 58226
rect 345678 58170 345774 58226
rect 345154 58102 345774 58170
rect 345154 58046 345250 58102
rect 345306 58046 345374 58102
rect 345430 58046 345498 58102
rect 345554 58046 345622 58102
rect 345678 58046 345774 58102
rect 345154 57978 345774 58046
rect 345154 57922 345250 57978
rect 345306 57922 345374 57978
rect 345430 57922 345498 57978
rect 345554 57922 345622 57978
rect 345678 57922 345774 57978
rect 343980 55412 344036 55422
rect 330874 46294 330970 46350
rect 331026 46294 331094 46350
rect 331150 46294 331218 46350
rect 331274 46294 331342 46350
rect 331398 46294 331494 46350
rect 330874 46226 331494 46294
rect 330874 46170 330970 46226
rect 331026 46170 331094 46226
rect 331150 46170 331218 46226
rect 331274 46170 331342 46226
rect 331398 46170 331494 46226
rect 330874 46102 331494 46170
rect 330874 46046 330970 46102
rect 331026 46046 331094 46102
rect 331150 46046 331218 46102
rect 331274 46046 331342 46102
rect 331398 46046 331494 46102
rect 330874 45978 331494 46046
rect 330874 45922 330970 45978
rect 331026 45922 331094 45978
rect 331150 45922 331218 45978
rect 331274 45922 331342 45978
rect 331398 45922 331494 45978
rect 330874 28350 331494 45922
rect 343532 47348 343588 47358
rect 343532 36596 343588 47292
rect 343532 36530 343588 36540
rect 343980 36484 344036 55356
rect 343980 36418 344036 36428
rect 345154 40350 345774 57922
rect 345154 40294 345250 40350
rect 345306 40294 345374 40350
rect 345430 40294 345498 40350
rect 345554 40294 345622 40350
rect 345678 40294 345774 40350
rect 345154 40226 345774 40294
rect 345154 40170 345250 40226
rect 345306 40170 345374 40226
rect 345430 40170 345498 40226
rect 345554 40170 345622 40226
rect 345678 40170 345774 40226
rect 345154 40102 345774 40170
rect 345154 40046 345250 40102
rect 345306 40046 345374 40102
rect 345430 40046 345498 40102
rect 345554 40046 345622 40102
rect 345678 40046 345774 40102
rect 345154 39978 345774 40046
rect 345154 39922 345250 39978
rect 345306 39922 345374 39978
rect 345430 39922 345498 39978
rect 345554 39922 345622 39978
rect 345678 39922 345774 39978
rect 330874 28294 330970 28350
rect 331026 28294 331094 28350
rect 331150 28294 331218 28350
rect 331274 28294 331342 28350
rect 331398 28294 331494 28350
rect 330874 28226 331494 28294
rect 330874 28170 330970 28226
rect 331026 28170 331094 28226
rect 331150 28170 331218 28226
rect 331274 28170 331342 28226
rect 331398 28170 331494 28226
rect 330874 28102 331494 28170
rect 330874 28046 330970 28102
rect 331026 28046 331094 28102
rect 331150 28046 331218 28102
rect 331274 28046 331342 28102
rect 331398 28046 331494 28102
rect 330874 27978 331494 28046
rect 330874 27922 330970 27978
rect 331026 27922 331094 27978
rect 331150 27922 331218 27978
rect 331274 27922 331342 27978
rect 331398 27922 331494 27978
rect 330874 10350 331494 27922
rect 330874 10294 330970 10350
rect 331026 10294 331094 10350
rect 331150 10294 331218 10350
rect 331274 10294 331342 10350
rect 331398 10294 331494 10350
rect 330874 10226 331494 10294
rect 330874 10170 330970 10226
rect 331026 10170 331094 10226
rect 331150 10170 331218 10226
rect 331274 10170 331342 10226
rect 331398 10170 331494 10226
rect 330874 10102 331494 10170
rect 330874 10046 330970 10102
rect 331026 10046 331094 10102
rect 331150 10046 331218 10102
rect 331274 10046 331342 10102
rect 331398 10046 331494 10102
rect 330874 9978 331494 10046
rect 330874 9922 330970 9978
rect 331026 9922 331094 9978
rect 331150 9922 331218 9978
rect 331274 9922 331342 9978
rect 331398 9922 331494 9978
rect 330874 -1120 331494 9922
rect 330874 -1176 330970 -1120
rect 331026 -1176 331094 -1120
rect 331150 -1176 331218 -1120
rect 331274 -1176 331342 -1120
rect 331398 -1176 331494 -1120
rect 330874 -1244 331494 -1176
rect 330874 -1300 330970 -1244
rect 331026 -1300 331094 -1244
rect 331150 -1300 331218 -1244
rect 331274 -1300 331342 -1244
rect 331398 -1300 331494 -1244
rect 330874 -1368 331494 -1300
rect 330874 -1424 330970 -1368
rect 331026 -1424 331094 -1368
rect 331150 -1424 331218 -1368
rect 331274 -1424 331342 -1368
rect 331398 -1424 331494 -1368
rect 330874 -1492 331494 -1424
rect 330874 -1548 330970 -1492
rect 331026 -1548 331094 -1492
rect 331150 -1548 331218 -1492
rect 331274 -1548 331342 -1492
rect 331398 -1548 331494 -1492
rect 330874 -1644 331494 -1548
rect 345154 22350 345774 39922
rect 346780 103012 346836 103022
rect 346780 42778 346836 102956
rect 346108 28532 346164 28542
rect 346108 28196 346164 28476
rect 346108 28130 346164 28140
rect 346780 26404 346836 42722
rect 346892 27860 346948 167468
rect 347340 162148 347396 162158
rect 347228 124516 347284 124526
rect 347116 119140 347172 119150
rect 347004 113764 347060 113774
rect 347004 39508 347060 113708
rect 347004 39442 347060 39452
rect 346892 27794 346948 27804
rect 347004 38278 347060 38286
rect 347116 38278 347172 119084
rect 347004 38276 347172 38278
rect 347060 38222 347172 38276
rect 346780 26338 346836 26348
rect 347004 24500 347060 38220
rect 347228 36932 347284 124460
rect 347228 31948 347284 36876
rect 347116 31892 347284 31948
rect 347116 26292 347172 31892
rect 347340 27412 347396 162092
rect 347452 28420 347508 172844
rect 347452 28354 347508 28364
rect 347564 28308 347620 178220
rect 347676 28532 347732 183596
rect 347676 28466 347732 28476
rect 348874 172350 349494 189922
rect 348874 172294 348970 172350
rect 349026 172294 349094 172350
rect 349150 172294 349218 172350
rect 349274 172294 349342 172350
rect 349398 172294 349494 172350
rect 348874 172226 349494 172294
rect 348874 172170 348970 172226
rect 349026 172170 349094 172226
rect 349150 172170 349218 172226
rect 349274 172170 349342 172226
rect 349398 172170 349494 172226
rect 348874 172102 349494 172170
rect 348874 172046 348970 172102
rect 349026 172046 349094 172102
rect 349150 172046 349218 172102
rect 349274 172046 349342 172102
rect 349398 172046 349494 172102
rect 348874 171978 349494 172046
rect 348874 171922 348970 171978
rect 349026 171922 349094 171978
rect 349150 171922 349218 171978
rect 349274 171922 349342 171978
rect 349398 171922 349494 171978
rect 348874 154350 349494 171922
rect 348874 154294 348970 154350
rect 349026 154294 349094 154350
rect 349150 154294 349218 154350
rect 349274 154294 349342 154350
rect 349398 154294 349494 154350
rect 348874 154226 349494 154294
rect 348874 154170 348970 154226
rect 349026 154170 349094 154226
rect 349150 154170 349218 154226
rect 349274 154170 349342 154226
rect 349398 154170 349494 154226
rect 348874 154102 349494 154170
rect 348874 154046 348970 154102
rect 349026 154046 349094 154102
rect 349150 154046 349218 154102
rect 349274 154046 349342 154102
rect 349398 154046 349494 154102
rect 348874 153978 349494 154046
rect 348874 153922 348970 153978
rect 349026 153922 349094 153978
rect 349150 153922 349218 153978
rect 349274 153922 349342 153978
rect 349398 153922 349494 153978
rect 348874 136350 349494 153922
rect 348874 136294 348970 136350
rect 349026 136294 349094 136350
rect 349150 136294 349218 136350
rect 349274 136294 349342 136350
rect 349398 136294 349494 136350
rect 348874 136226 349494 136294
rect 348874 136170 348970 136226
rect 349026 136170 349094 136226
rect 349150 136170 349218 136226
rect 349274 136170 349342 136226
rect 349398 136170 349494 136226
rect 348874 136102 349494 136170
rect 348874 136046 348970 136102
rect 349026 136046 349094 136102
rect 349150 136046 349218 136102
rect 349274 136046 349342 136102
rect 349398 136046 349494 136102
rect 348874 135978 349494 136046
rect 348874 135922 348970 135978
rect 349026 135922 349094 135978
rect 349150 135922 349218 135978
rect 349274 135922 349342 135978
rect 349398 135922 349494 135978
rect 348874 118350 349494 135922
rect 348874 118294 348970 118350
rect 349026 118294 349094 118350
rect 349150 118294 349218 118350
rect 349274 118294 349342 118350
rect 349398 118294 349494 118350
rect 348874 118226 349494 118294
rect 348874 118170 348970 118226
rect 349026 118170 349094 118226
rect 349150 118170 349218 118226
rect 349274 118170 349342 118226
rect 349398 118170 349494 118226
rect 348874 118102 349494 118170
rect 348874 118046 348970 118102
rect 349026 118046 349094 118102
rect 349150 118046 349218 118102
rect 349274 118046 349342 118102
rect 349398 118046 349494 118102
rect 348874 117978 349494 118046
rect 348874 117922 348970 117978
rect 349026 117922 349094 117978
rect 349150 117922 349218 117978
rect 349274 117922 349342 117978
rect 349398 117922 349494 117978
rect 348874 100350 349494 117922
rect 348874 100294 348970 100350
rect 349026 100294 349094 100350
rect 349150 100294 349218 100350
rect 349274 100294 349342 100350
rect 349398 100294 349494 100350
rect 348874 100226 349494 100294
rect 348874 100170 348970 100226
rect 349026 100170 349094 100226
rect 349150 100170 349218 100226
rect 349274 100170 349342 100226
rect 349398 100170 349494 100226
rect 348874 100102 349494 100170
rect 348874 100046 348970 100102
rect 349026 100046 349094 100102
rect 349150 100046 349218 100102
rect 349274 100046 349342 100102
rect 349398 100046 349494 100102
rect 348874 99978 349494 100046
rect 348874 99922 348970 99978
rect 349026 99922 349094 99978
rect 349150 99922 349218 99978
rect 349274 99922 349342 99978
rect 349398 99922 349494 99978
rect 348874 82350 349494 99922
rect 348874 82294 348970 82350
rect 349026 82294 349094 82350
rect 349150 82294 349218 82350
rect 349274 82294 349342 82350
rect 349398 82294 349494 82350
rect 348874 82226 349494 82294
rect 348874 82170 348970 82226
rect 349026 82170 349094 82226
rect 349150 82170 349218 82226
rect 349274 82170 349342 82226
rect 349398 82170 349494 82226
rect 348874 82102 349494 82170
rect 348874 82046 348970 82102
rect 349026 82046 349094 82102
rect 349150 82046 349218 82102
rect 349274 82046 349342 82102
rect 349398 82046 349494 82102
rect 348874 81978 349494 82046
rect 348874 81922 348970 81978
rect 349026 81922 349094 81978
rect 349150 81922 349218 81978
rect 349274 81922 349342 81978
rect 349398 81922 349494 81978
rect 348874 64350 349494 81922
rect 348874 64294 348970 64350
rect 349026 64294 349094 64350
rect 349150 64294 349218 64350
rect 349274 64294 349342 64350
rect 349398 64294 349494 64350
rect 348874 64226 349494 64294
rect 348874 64170 348970 64226
rect 349026 64170 349094 64226
rect 349150 64170 349218 64226
rect 349274 64170 349342 64226
rect 349398 64170 349494 64226
rect 348874 64102 349494 64170
rect 348874 64046 348970 64102
rect 349026 64046 349094 64102
rect 349150 64046 349218 64102
rect 349274 64046 349342 64102
rect 349398 64046 349494 64102
rect 348874 63978 349494 64046
rect 348874 63922 348970 63978
rect 349026 63922 349094 63978
rect 349150 63922 349218 63978
rect 349274 63922 349342 63978
rect 349398 63922 349494 63978
rect 348874 46350 349494 63922
rect 349916 65604 349972 65614
rect 349916 55468 349972 65548
rect 548940 59878 548996 59888
rect 548940 55468 548996 59822
rect 349916 55412 350308 55468
rect 348874 46294 348970 46350
rect 349026 46294 349094 46350
rect 349150 46294 349218 46350
rect 349274 46294 349342 46350
rect 349398 46294 349494 46350
rect 348874 46226 349494 46294
rect 348874 46170 348970 46226
rect 349026 46170 349094 46226
rect 349150 46170 349218 46226
rect 349274 46170 349342 46226
rect 349398 46170 349494 46226
rect 348874 46102 349494 46170
rect 348874 46046 348970 46102
rect 349026 46046 349094 46102
rect 349150 46046 349218 46102
rect 349274 46046 349342 46102
rect 349398 46046 349494 46102
rect 348874 45978 349494 46046
rect 348874 45922 348970 45978
rect 349026 45922 349094 45978
rect 349150 45922 349218 45978
rect 349274 45922 349342 45978
rect 349398 45922 349494 45978
rect 347564 28242 347620 28252
rect 348874 28350 349494 45922
rect 350140 51380 350196 51390
rect 349916 45444 349972 45454
rect 349580 45332 349636 45342
rect 349580 36372 349636 45276
rect 349580 36306 349636 36316
rect 348874 28294 348970 28350
rect 349026 28294 349094 28350
rect 349150 28294 349218 28350
rect 349274 28294 349342 28350
rect 349398 28294 349494 28350
rect 347340 27346 347396 27356
rect 348874 28226 349494 28294
rect 348874 28170 348970 28226
rect 349026 28170 349094 28226
rect 349150 28170 349218 28226
rect 349274 28170 349342 28226
rect 349398 28170 349494 28226
rect 348874 28102 349494 28170
rect 348874 28046 348970 28102
rect 349026 28046 349094 28102
rect 349150 28046 349218 28102
rect 349274 28046 349342 28102
rect 349398 28046 349494 28102
rect 348874 27978 349494 28046
rect 348874 27922 348970 27978
rect 349026 27922 349094 27978
rect 349150 27922 349218 27978
rect 349274 27922 349342 27978
rect 349398 27922 349494 27978
rect 347116 26226 347172 26236
rect 347004 24434 347060 24444
rect 345154 22294 345250 22350
rect 345306 22294 345374 22350
rect 345430 22294 345498 22350
rect 345554 22294 345622 22350
rect 345678 22294 345774 22350
rect 345154 22226 345774 22294
rect 345154 22170 345250 22226
rect 345306 22170 345374 22226
rect 345430 22170 345498 22226
rect 345554 22170 345622 22226
rect 345678 22170 345774 22226
rect 345154 22102 345774 22170
rect 345154 22046 345250 22102
rect 345306 22046 345374 22102
rect 345430 22046 345498 22102
rect 345554 22046 345622 22102
rect 345678 22046 345774 22102
rect 345154 21978 345774 22046
rect 345154 21922 345250 21978
rect 345306 21922 345374 21978
rect 345430 21922 345498 21978
rect 345554 21922 345622 21978
rect 345678 21922 345774 21978
rect 345154 4350 345774 21922
rect 345154 4294 345250 4350
rect 345306 4294 345374 4350
rect 345430 4294 345498 4350
rect 345554 4294 345622 4350
rect 345678 4294 345774 4350
rect 345154 4226 345774 4294
rect 345154 4170 345250 4226
rect 345306 4170 345374 4226
rect 345430 4170 345498 4226
rect 345554 4170 345622 4226
rect 345678 4170 345774 4226
rect 345154 4102 345774 4170
rect 345154 4046 345250 4102
rect 345306 4046 345374 4102
rect 345430 4046 345498 4102
rect 345554 4046 345622 4102
rect 345678 4046 345774 4102
rect 345154 3978 345774 4046
rect 345154 3922 345250 3978
rect 345306 3922 345374 3978
rect 345430 3922 345498 3978
rect 345554 3922 345622 3978
rect 345678 3922 345774 3978
rect 345154 -160 345774 3922
rect 345154 -216 345250 -160
rect 345306 -216 345374 -160
rect 345430 -216 345498 -160
rect 345554 -216 345622 -160
rect 345678 -216 345774 -160
rect 345154 -284 345774 -216
rect 345154 -340 345250 -284
rect 345306 -340 345374 -284
rect 345430 -340 345498 -284
rect 345554 -340 345622 -284
rect 345678 -340 345774 -284
rect 345154 -408 345774 -340
rect 345154 -464 345250 -408
rect 345306 -464 345374 -408
rect 345430 -464 345498 -408
rect 345554 -464 345622 -408
rect 345678 -464 345774 -408
rect 345154 -532 345774 -464
rect 345154 -588 345250 -532
rect 345306 -588 345374 -532
rect 345430 -588 345498 -532
rect 345554 -588 345622 -532
rect 345678 -588 345774 -532
rect 345154 -1644 345774 -588
rect 348874 10350 349494 27922
rect 349916 34916 349972 45388
rect 350140 35252 350196 51324
rect 350140 35186 350196 35196
rect 349916 24612 349972 34860
rect 350252 25138 350308 55412
rect 548828 55412 548996 55468
rect 548716 54658 548772 54668
rect 548492 54602 548716 54658
rect 350588 53396 350644 53406
rect 350476 52052 350532 52062
rect 350252 25072 350308 25082
rect 350364 48468 350420 48478
rect 350364 33572 350420 48412
rect 349916 24546 349972 24556
rect 350364 20916 350420 33516
rect 350364 20850 350420 20860
rect 350476 21700 350532 51996
rect 350588 35028 350644 53340
rect 525308 43138 525364 43148
rect 516460 42958 516516 42968
rect 525308 42958 525364 43082
rect 496300 41524 496356 41534
rect 436268 41338 436324 41348
rect 363154 40350 363774 41266
rect 363154 40294 363250 40350
rect 363306 40294 363374 40350
rect 363430 40294 363498 40350
rect 363554 40294 363622 40350
rect 363678 40294 363774 40350
rect 363154 40226 363774 40294
rect 363154 40170 363250 40226
rect 363306 40170 363374 40226
rect 363430 40170 363498 40226
rect 363554 40170 363622 40226
rect 363678 40170 363774 40226
rect 363154 40102 363774 40170
rect 363154 40046 363250 40102
rect 363306 40046 363374 40102
rect 363430 40046 363498 40102
rect 363554 40046 363622 40102
rect 363678 40046 363774 40102
rect 363154 39978 363774 40046
rect 363154 39922 363250 39978
rect 363306 39922 363374 39978
rect 363430 39922 363498 39978
rect 363554 39922 363622 39978
rect 363678 39922 363774 39978
rect 354508 37738 354564 37754
rect 354508 37650 354564 37660
rect 362908 37044 362964 37054
rect 362908 36950 362964 36962
rect 350588 34962 350644 34972
rect 350476 17556 350532 21644
rect 350476 17490 350532 17500
rect 363154 22350 363774 39922
rect 363154 22294 363250 22350
rect 363306 22294 363374 22350
rect 363430 22294 363498 22350
rect 363554 22294 363622 22350
rect 363678 22294 363774 22350
rect 363154 22226 363774 22294
rect 363154 22170 363250 22226
rect 363306 22170 363374 22226
rect 363430 22170 363498 22226
rect 363554 22170 363622 22226
rect 363678 22170 363774 22226
rect 363154 22102 363774 22170
rect 363154 22046 363250 22102
rect 363306 22046 363374 22102
rect 363430 22046 363498 22102
rect 363554 22046 363622 22102
rect 363678 22046 363774 22102
rect 363154 21978 363774 22046
rect 363154 21922 363250 21978
rect 363306 21922 363374 21978
rect 363430 21922 363498 21978
rect 363554 21922 363622 21978
rect 363678 21922 363774 21978
rect 348874 10294 348970 10350
rect 349026 10294 349094 10350
rect 349150 10294 349218 10350
rect 349274 10294 349342 10350
rect 349398 10294 349494 10350
rect 348874 10226 349494 10294
rect 348874 10170 348970 10226
rect 349026 10170 349094 10226
rect 349150 10170 349218 10226
rect 349274 10170 349342 10226
rect 349398 10170 349494 10226
rect 348874 10102 349494 10170
rect 348874 10046 348970 10102
rect 349026 10046 349094 10102
rect 349150 10046 349218 10102
rect 349274 10046 349342 10102
rect 349398 10046 349494 10102
rect 348874 9978 349494 10046
rect 348874 9922 348970 9978
rect 349026 9922 349094 9978
rect 349150 9922 349218 9978
rect 349274 9922 349342 9978
rect 349398 9922 349494 9978
rect 348874 -1120 349494 9922
rect 348874 -1176 348970 -1120
rect 349026 -1176 349094 -1120
rect 349150 -1176 349218 -1120
rect 349274 -1176 349342 -1120
rect 349398 -1176 349494 -1120
rect 348874 -1244 349494 -1176
rect 348874 -1300 348970 -1244
rect 349026 -1300 349094 -1244
rect 349150 -1300 349218 -1244
rect 349274 -1300 349342 -1244
rect 349398 -1300 349494 -1244
rect 348874 -1368 349494 -1300
rect 348874 -1424 348970 -1368
rect 349026 -1424 349094 -1368
rect 349150 -1424 349218 -1368
rect 349274 -1424 349342 -1368
rect 349398 -1424 349494 -1368
rect 348874 -1492 349494 -1424
rect 348874 -1548 348970 -1492
rect 349026 -1548 349094 -1492
rect 349150 -1548 349218 -1492
rect 349274 -1548 349342 -1492
rect 349398 -1548 349494 -1492
rect 348874 -1644 349494 -1548
rect 363154 4350 363774 21922
rect 363154 4294 363250 4350
rect 363306 4294 363374 4350
rect 363430 4294 363498 4350
rect 363554 4294 363622 4350
rect 363678 4294 363774 4350
rect 363154 4226 363774 4294
rect 363154 4170 363250 4226
rect 363306 4170 363374 4226
rect 363430 4170 363498 4226
rect 363554 4170 363622 4226
rect 363678 4170 363774 4226
rect 363154 4102 363774 4170
rect 363154 4046 363250 4102
rect 363306 4046 363374 4102
rect 363430 4046 363498 4102
rect 363554 4046 363622 4102
rect 363678 4046 363774 4102
rect 363154 3978 363774 4046
rect 363154 3922 363250 3978
rect 363306 3922 363374 3978
rect 363430 3922 363498 3978
rect 363554 3922 363622 3978
rect 363678 3922 363774 3978
rect 363154 -160 363774 3922
rect 363154 -216 363250 -160
rect 363306 -216 363374 -160
rect 363430 -216 363498 -160
rect 363554 -216 363622 -160
rect 363678 -216 363774 -160
rect 363154 -284 363774 -216
rect 363154 -340 363250 -284
rect 363306 -340 363374 -284
rect 363430 -340 363498 -284
rect 363554 -340 363622 -284
rect 363678 -340 363774 -284
rect 363154 -408 363774 -340
rect 363154 -464 363250 -408
rect 363306 -464 363374 -408
rect 363430 -464 363498 -408
rect 363554 -464 363622 -408
rect 363678 -464 363774 -408
rect 363154 -532 363774 -464
rect 363154 -588 363250 -532
rect 363306 -588 363374 -532
rect 363430 -588 363498 -532
rect 363554 -588 363622 -532
rect 363678 -588 363774 -532
rect 363154 -1644 363774 -588
rect 366874 28350 367494 41266
rect 381154 40350 381774 41266
rect 381154 40294 381250 40350
rect 381306 40294 381374 40350
rect 381430 40294 381498 40350
rect 381554 40294 381622 40350
rect 381678 40294 381774 40350
rect 381154 40226 381774 40294
rect 381154 40170 381250 40226
rect 381306 40170 381374 40226
rect 381430 40170 381498 40226
rect 381554 40170 381622 40226
rect 381678 40170 381774 40226
rect 381154 40102 381774 40170
rect 381154 40046 381250 40102
rect 381306 40046 381374 40102
rect 381430 40046 381498 40102
rect 381554 40046 381622 40102
rect 381678 40046 381774 40102
rect 381154 39978 381774 40046
rect 381154 39922 381250 39978
rect 381306 39922 381374 39978
rect 381430 39922 381498 39978
rect 381554 39922 381622 39978
rect 381678 39922 381774 39978
rect 366874 28294 366970 28350
rect 367026 28294 367094 28350
rect 367150 28294 367218 28350
rect 367274 28294 367342 28350
rect 367398 28294 367494 28350
rect 366874 28226 367494 28294
rect 366874 28170 366970 28226
rect 367026 28170 367094 28226
rect 367150 28170 367218 28226
rect 367274 28170 367342 28226
rect 367398 28170 367494 28226
rect 366874 28102 367494 28170
rect 366874 28046 366970 28102
rect 367026 28046 367094 28102
rect 367150 28046 367218 28102
rect 367274 28046 367342 28102
rect 367398 28046 367494 28102
rect 366874 27978 367494 28046
rect 366874 27922 366970 27978
rect 367026 27922 367094 27978
rect 367150 27922 367218 27978
rect 367274 27922 367342 27978
rect 367398 27922 367494 27978
rect 366874 10350 367494 27922
rect 371308 28644 371364 28654
rect 371308 24958 371364 28588
rect 371308 24892 371364 24902
rect 366874 10294 366970 10350
rect 367026 10294 367094 10350
rect 367150 10294 367218 10350
rect 367274 10294 367342 10350
rect 367398 10294 367494 10350
rect 366874 10226 367494 10294
rect 366874 10170 366970 10226
rect 367026 10170 367094 10226
rect 367150 10170 367218 10226
rect 367274 10170 367342 10226
rect 367398 10170 367494 10226
rect 366874 10102 367494 10170
rect 366874 10046 366970 10102
rect 367026 10046 367094 10102
rect 367150 10046 367218 10102
rect 367274 10046 367342 10102
rect 367398 10046 367494 10102
rect 366874 9978 367494 10046
rect 366874 9922 366970 9978
rect 367026 9922 367094 9978
rect 367150 9922 367218 9978
rect 367274 9922 367342 9978
rect 367398 9922 367494 9978
rect 366874 -1120 367494 9922
rect 366874 -1176 366970 -1120
rect 367026 -1176 367094 -1120
rect 367150 -1176 367218 -1120
rect 367274 -1176 367342 -1120
rect 367398 -1176 367494 -1120
rect 366874 -1244 367494 -1176
rect 366874 -1300 366970 -1244
rect 367026 -1300 367094 -1244
rect 367150 -1300 367218 -1244
rect 367274 -1300 367342 -1244
rect 367398 -1300 367494 -1244
rect 366874 -1368 367494 -1300
rect 366874 -1424 366970 -1368
rect 367026 -1424 367094 -1368
rect 367150 -1424 367218 -1368
rect 367274 -1424 367342 -1368
rect 367398 -1424 367494 -1368
rect 366874 -1492 367494 -1424
rect 366874 -1548 366970 -1492
rect 367026 -1548 367094 -1492
rect 367150 -1548 367218 -1492
rect 367274 -1548 367342 -1492
rect 367398 -1548 367494 -1492
rect 366874 -1644 367494 -1548
rect 381154 22350 381774 39922
rect 383852 37044 383908 37054
rect 383852 24418 383908 36988
rect 383852 24352 383908 24362
rect 384874 28350 385494 40964
rect 399154 40350 399774 41266
rect 399154 40294 399250 40350
rect 399306 40294 399374 40350
rect 399430 40294 399498 40350
rect 399554 40294 399622 40350
rect 399678 40294 399774 40350
rect 399154 40226 399774 40294
rect 399154 40170 399250 40226
rect 399306 40170 399374 40226
rect 399430 40170 399498 40226
rect 399554 40170 399622 40226
rect 399678 40170 399774 40226
rect 399154 40102 399774 40170
rect 399154 40046 399250 40102
rect 399306 40046 399374 40102
rect 399430 40046 399498 40102
rect 399554 40046 399622 40102
rect 399678 40046 399774 40102
rect 399154 39978 399774 40046
rect 399154 39922 399250 39978
rect 399306 39922 399374 39978
rect 399430 39922 399498 39978
rect 399554 39922 399622 39978
rect 399678 39922 399774 39978
rect 394828 29652 394884 29662
rect 394828 29558 394884 29582
rect 384874 28294 384970 28350
rect 385026 28294 385094 28350
rect 385150 28294 385218 28350
rect 385274 28294 385342 28350
rect 385398 28294 385494 28350
rect 384874 28226 385494 28294
rect 384874 28170 384970 28226
rect 385026 28170 385094 28226
rect 385150 28170 385218 28226
rect 385274 28170 385342 28226
rect 385398 28170 385494 28226
rect 384874 28102 385494 28170
rect 384874 28046 384970 28102
rect 385026 28046 385094 28102
rect 385150 28046 385218 28102
rect 385274 28046 385342 28102
rect 385398 28046 385494 28102
rect 384874 27978 385494 28046
rect 384874 27922 384970 27978
rect 385026 27922 385094 27978
rect 385150 27922 385218 27978
rect 385274 27922 385342 27978
rect 385398 27922 385494 27978
rect 381154 22294 381250 22350
rect 381306 22294 381374 22350
rect 381430 22294 381498 22350
rect 381554 22294 381622 22350
rect 381678 22294 381774 22350
rect 381154 22226 381774 22294
rect 381154 22170 381250 22226
rect 381306 22170 381374 22226
rect 381430 22170 381498 22226
rect 381554 22170 381622 22226
rect 381678 22170 381774 22226
rect 381154 22102 381774 22170
rect 381154 22046 381250 22102
rect 381306 22046 381374 22102
rect 381430 22046 381498 22102
rect 381554 22046 381622 22102
rect 381678 22046 381774 22102
rect 381154 21978 381774 22046
rect 381154 21922 381250 21978
rect 381306 21922 381374 21978
rect 381430 21922 381498 21978
rect 381554 21922 381622 21978
rect 381678 21922 381774 21978
rect 381154 4350 381774 21922
rect 381154 4294 381250 4350
rect 381306 4294 381374 4350
rect 381430 4294 381498 4350
rect 381554 4294 381622 4350
rect 381678 4294 381774 4350
rect 381154 4226 381774 4294
rect 381154 4170 381250 4226
rect 381306 4170 381374 4226
rect 381430 4170 381498 4226
rect 381554 4170 381622 4226
rect 381678 4170 381774 4226
rect 381154 4102 381774 4170
rect 381154 4046 381250 4102
rect 381306 4046 381374 4102
rect 381430 4046 381498 4102
rect 381554 4046 381622 4102
rect 381678 4046 381774 4102
rect 381154 3978 381774 4046
rect 381154 3922 381250 3978
rect 381306 3922 381374 3978
rect 381430 3922 381498 3978
rect 381554 3922 381622 3978
rect 381678 3922 381774 3978
rect 381154 -160 381774 3922
rect 381154 -216 381250 -160
rect 381306 -216 381374 -160
rect 381430 -216 381498 -160
rect 381554 -216 381622 -160
rect 381678 -216 381774 -160
rect 381154 -284 381774 -216
rect 381154 -340 381250 -284
rect 381306 -340 381374 -284
rect 381430 -340 381498 -284
rect 381554 -340 381622 -284
rect 381678 -340 381774 -284
rect 381154 -408 381774 -340
rect 381154 -464 381250 -408
rect 381306 -464 381374 -408
rect 381430 -464 381498 -408
rect 381554 -464 381622 -408
rect 381678 -464 381774 -408
rect 381154 -532 381774 -464
rect 381154 -588 381250 -532
rect 381306 -588 381374 -532
rect 381430 -588 381498 -532
rect 381554 -588 381622 -532
rect 381678 -588 381774 -532
rect 381154 -1644 381774 -588
rect 384874 10350 385494 27922
rect 384874 10294 384970 10350
rect 385026 10294 385094 10350
rect 385150 10294 385218 10350
rect 385274 10294 385342 10350
rect 385398 10294 385494 10350
rect 384874 10226 385494 10294
rect 384874 10170 384970 10226
rect 385026 10170 385094 10226
rect 385150 10170 385218 10226
rect 385274 10170 385342 10226
rect 385398 10170 385494 10226
rect 384874 10102 385494 10170
rect 384874 10046 384970 10102
rect 385026 10046 385094 10102
rect 385150 10046 385218 10102
rect 385274 10046 385342 10102
rect 385398 10046 385494 10102
rect 384874 9978 385494 10046
rect 384874 9922 384970 9978
rect 385026 9922 385094 9978
rect 385150 9922 385218 9978
rect 385274 9922 385342 9978
rect 385398 9922 385494 9978
rect 384874 -1120 385494 9922
rect 384874 -1176 384970 -1120
rect 385026 -1176 385094 -1120
rect 385150 -1176 385218 -1120
rect 385274 -1176 385342 -1120
rect 385398 -1176 385494 -1120
rect 384874 -1244 385494 -1176
rect 384874 -1300 384970 -1244
rect 385026 -1300 385094 -1244
rect 385150 -1300 385218 -1244
rect 385274 -1300 385342 -1244
rect 385398 -1300 385494 -1244
rect 384874 -1368 385494 -1300
rect 384874 -1424 384970 -1368
rect 385026 -1424 385094 -1368
rect 385150 -1424 385218 -1368
rect 385274 -1424 385342 -1368
rect 385398 -1424 385494 -1368
rect 384874 -1492 385494 -1424
rect 384874 -1548 384970 -1492
rect 385026 -1548 385094 -1492
rect 385150 -1548 385218 -1492
rect 385274 -1548 385342 -1492
rect 385398 -1548 385494 -1492
rect 384874 -1644 385494 -1548
rect 399154 22350 399774 39922
rect 399154 22294 399250 22350
rect 399306 22294 399374 22350
rect 399430 22294 399498 22350
rect 399554 22294 399622 22350
rect 399678 22294 399774 22350
rect 399154 22226 399774 22294
rect 399154 22170 399250 22226
rect 399306 22170 399374 22226
rect 399430 22170 399498 22226
rect 399554 22170 399622 22226
rect 399678 22170 399774 22226
rect 399154 22102 399774 22170
rect 399154 22046 399250 22102
rect 399306 22046 399374 22102
rect 399430 22046 399498 22102
rect 399554 22046 399622 22102
rect 399678 22046 399774 22102
rect 399154 21978 399774 22046
rect 399154 21922 399250 21978
rect 399306 21922 399374 21978
rect 399430 21922 399498 21978
rect 399554 21922 399622 21978
rect 399678 21922 399774 21978
rect 399154 4350 399774 21922
rect 399154 4294 399250 4350
rect 399306 4294 399374 4350
rect 399430 4294 399498 4350
rect 399554 4294 399622 4350
rect 399678 4294 399774 4350
rect 399154 4226 399774 4294
rect 399154 4170 399250 4226
rect 399306 4170 399374 4226
rect 399430 4170 399498 4226
rect 399554 4170 399622 4226
rect 399678 4170 399774 4226
rect 399154 4102 399774 4170
rect 399154 4046 399250 4102
rect 399306 4046 399374 4102
rect 399430 4046 399498 4102
rect 399554 4046 399622 4102
rect 399678 4046 399774 4102
rect 399154 3978 399774 4046
rect 399154 3922 399250 3978
rect 399306 3922 399374 3978
rect 399430 3922 399498 3978
rect 399554 3922 399622 3978
rect 399678 3922 399774 3978
rect 399154 -160 399774 3922
rect 399154 -216 399250 -160
rect 399306 -216 399374 -160
rect 399430 -216 399498 -160
rect 399554 -216 399622 -160
rect 399678 -216 399774 -160
rect 399154 -284 399774 -216
rect 399154 -340 399250 -284
rect 399306 -340 399374 -284
rect 399430 -340 399498 -284
rect 399554 -340 399622 -284
rect 399678 -340 399774 -284
rect 399154 -408 399774 -340
rect 399154 -464 399250 -408
rect 399306 -464 399374 -408
rect 399430 -464 399498 -408
rect 399554 -464 399622 -408
rect 399678 -464 399774 -408
rect 399154 -532 399774 -464
rect 399154 -588 399250 -532
rect 399306 -588 399374 -532
rect 399430 -588 399498 -532
rect 399554 -588 399622 -532
rect 399678 -588 399774 -532
rect 399154 -1644 399774 -588
rect 402874 28350 403494 41266
rect 402874 28294 402970 28350
rect 403026 28294 403094 28350
rect 403150 28294 403218 28350
rect 403274 28294 403342 28350
rect 403398 28294 403494 28350
rect 402874 28226 403494 28294
rect 402874 28170 402970 28226
rect 403026 28170 403094 28226
rect 403150 28170 403218 28226
rect 403274 28170 403342 28226
rect 403398 28170 403494 28226
rect 402874 28102 403494 28170
rect 402874 28046 402970 28102
rect 403026 28046 403094 28102
rect 403150 28046 403218 28102
rect 403274 28046 403342 28102
rect 403398 28046 403494 28102
rect 402874 27978 403494 28046
rect 402874 27922 402970 27978
rect 403026 27922 403094 27978
rect 403150 27922 403218 27978
rect 403274 27922 403342 27978
rect 403398 27922 403494 27978
rect 402874 10350 403494 27922
rect 402874 10294 402970 10350
rect 403026 10294 403094 10350
rect 403150 10294 403218 10350
rect 403274 10294 403342 10350
rect 403398 10294 403494 10350
rect 402874 10226 403494 10294
rect 402874 10170 402970 10226
rect 403026 10170 403094 10226
rect 403150 10170 403218 10226
rect 403274 10170 403342 10226
rect 403398 10170 403494 10226
rect 402874 10102 403494 10170
rect 402874 10046 402970 10102
rect 403026 10046 403094 10102
rect 403150 10046 403218 10102
rect 403274 10046 403342 10102
rect 403398 10046 403494 10102
rect 402874 9978 403494 10046
rect 402874 9922 402970 9978
rect 403026 9922 403094 9978
rect 403150 9922 403218 9978
rect 403274 9922 403342 9978
rect 403398 9922 403494 9978
rect 402874 -1120 403494 9922
rect 402874 -1176 402970 -1120
rect 403026 -1176 403094 -1120
rect 403150 -1176 403218 -1120
rect 403274 -1176 403342 -1120
rect 403398 -1176 403494 -1120
rect 402874 -1244 403494 -1176
rect 402874 -1300 402970 -1244
rect 403026 -1300 403094 -1244
rect 403150 -1300 403218 -1244
rect 403274 -1300 403342 -1244
rect 403398 -1300 403494 -1244
rect 402874 -1368 403494 -1300
rect 402874 -1424 402970 -1368
rect 403026 -1424 403094 -1368
rect 403150 -1424 403218 -1368
rect 403274 -1424 403342 -1368
rect 403398 -1424 403494 -1368
rect 402874 -1492 403494 -1424
rect 402874 -1548 402970 -1492
rect 403026 -1548 403094 -1492
rect 403150 -1548 403218 -1492
rect 403274 -1548 403342 -1492
rect 403398 -1548 403494 -1492
rect 402874 -1644 403494 -1548
rect 417154 40350 417774 41266
rect 417154 40294 417250 40350
rect 417306 40294 417374 40350
rect 417430 40294 417498 40350
rect 417554 40294 417622 40350
rect 417678 40294 417774 40350
rect 417154 40226 417774 40294
rect 417154 40170 417250 40226
rect 417306 40170 417374 40226
rect 417430 40170 417498 40226
rect 417554 40170 417622 40226
rect 417678 40170 417774 40226
rect 417154 40102 417774 40170
rect 417154 40046 417250 40102
rect 417306 40046 417374 40102
rect 417430 40046 417498 40102
rect 417554 40046 417622 40102
rect 417678 40046 417774 40102
rect 417154 39978 417774 40046
rect 417154 39922 417250 39978
rect 417306 39922 417374 39978
rect 417430 39922 417498 39978
rect 417554 39922 417622 39978
rect 417678 39922 417774 39978
rect 417154 22350 417774 39922
rect 419692 39732 419748 39756
rect 418348 39718 418404 39728
rect 418348 34498 418404 39662
rect 419692 39652 419748 39662
rect 418348 34432 418404 34442
rect 417154 22294 417250 22350
rect 417306 22294 417374 22350
rect 417430 22294 417498 22350
rect 417554 22294 417622 22350
rect 417678 22294 417774 22350
rect 417154 22226 417774 22294
rect 417154 22170 417250 22226
rect 417306 22170 417374 22226
rect 417430 22170 417498 22226
rect 417554 22170 417622 22226
rect 417678 22170 417774 22226
rect 417154 22102 417774 22170
rect 417154 22046 417250 22102
rect 417306 22046 417374 22102
rect 417430 22046 417498 22102
rect 417554 22046 417622 22102
rect 417678 22046 417774 22102
rect 417154 21978 417774 22046
rect 417154 21922 417250 21978
rect 417306 21922 417374 21978
rect 417430 21922 417498 21978
rect 417554 21922 417622 21978
rect 417678 21922 417774 21978
rect 417154 4350 417774 21922
rect 417154 4294 417250 4350
rect 417306 4294 417374 4350
rect 417430 4294 417498 4350
rect 417554 4294 417622 4350
rect 417678 4294 417774 4350
rect 417154 4226 417774 4294
rect 417154 4170 417250 4226
rect 417306 4170 417374 4226
rect 417430 4170 417498 4226
rect 417554 4170 417622 4226
rect 417678 4170 417774 4226
rect 417154 4102 417774 4170
rect 417154 4046 417250 4102
rect 417306 4046 417374 4102
rect 417430 4046 417498 4102
rect 417554 4046 417622 4102
rect 417678 4046 417774 4102
rect 417154 3978 417774 4046
rect 417154 3922 417250 3978
rect 417306 3922 417374 3978
rect 417430 3922 417498 3978
rect 417554 3922 417622 3978
rect 417678 3922 417774 3978
rect 417154 -160 417774 3922
rect 417154 -216 417250 -160
rect 417306 -216 417374 -160
rect 417430 -216 417498 -160
rect 417554 -216 417622 -160
rect 417678 -216 417774 -160
rect 417154 -284 417774 -216
rect 417154 -340 417250 -284
rect 417306 -340 417374 -284
rect 417430 -340 417498 -284
rect 417554 -340 417622 -284
rect 417678 -340 417774 -284
rect 417154 -408 417774 -340
rect 417154 -464 417250 -408
rect 417306 -464 417374 -408
rect 417430 -464 417498 -408
rect 417554 -464 417622 -408
rect 417678 -464 417774 -408
rect 417154 -532 417774 -464
rect 417154 -588 417250 -532
rect 417306 -588 417374 -532
rect 417430 -588 417498 -532
rect 417554 -588 417622 -532
rect 417678 -588 417774 -532
rect 417154 -1644 417774 -588
rect 420874 28350 421494 41266
rect 431788 41158 431844 41168
rect 431788 40740 431844 41102
rect 423388 35364 423444 35374
rect 423388 35218 423444 35308
rect 423388 35152 423444 35162
rect 431788 29458 431844 40684
rect 431788 29392 431844 29402
rect 435154 40350 435774 40964
rect 436268 40516 436324 41282
rect 483868 41300 483924 41310
rect 436268 40450 436324 40460
rect 435154 40294 435250 40350
rect 435306 40294 435374 40350
rect 435430 40294 435498 40350
rect 435554 40294 435622 40350
rect 435678 40294 435774 40350
rect 435154 40226 435774 40294
rect 435154 40170 435250 40226
rect 435306 40170 435374 40226
rect 435430 40170 435498 40226
rect 435554 40170 435622 40226
rect 435678 40170 435774 40226
rect 435154 40102 435774 40170
rect 435154 40046 435250 40102
rect 435306 40046 435374 40102
rect 435430 40046 435498 40102
rect 435554 40046 435622 40102
rect 435678 40046 435774 40102
rect 435154 39978 435774 40046
rect 435154 39922 435250 39978
rect 435306 39922 435374 39978
rect 435430 39922 435498 39978
rect 435554 39922 435622 39978
rect 435678 39922 435774 39978
rect 420874 28294 420970 28350
rect 421026 28294 421094 28350
rect 421150 28294 421218 28350
rect 421274 28294 421342 28350
rect 421398 28294 421494 28350
rect 420874 28226 421494 28294
rect 420874 28170 420970 28226
rect 421026 28170 421094 28226
rect 421150 28170 421218 28226
rect 421274 28170 421342 28226
rect 421398 28170 421494 28226
rect 420874 28102 421494 28170
rect 420874 28046 420970 28102
rect 421026 28046 421094 28102
rect 421150 28046 421218 28102
rect 421274 28046 421342 28102
rect 421398 28046 421494 28102
rect 420874 27978 421494 28046
rect 420874 27922 420970 27978
rect 421026 27922 421094 27978
rect 421150 27922 421218 27978
rect 421274 27922 421342 27978
rect 421398 27922 421494 27978
rect 420874 10350 421494 27922
rect 420874 10294 420970 10350
rect 421026 10294 421094 10350
rect 421150 10294 421218 10350
rect 421274 10294 421342 10350
rect 421398 10294 421494 10350
rect 420874 10226 421494 10294
rect 420874 10170 420970 10226
rect 421026 10170 421094 10226
rect 421150 10170 421218 10226
rect 421274 10170 421342 10226
rect 421398 10170 421494 10226
rect 420874 10102 421494 10170
rect 420874 10046 420970 10102
rect 421026 10046 421094 10102
rect 421150 10046 421218 10102
rect 421274 10046 421342 10102
rect 421398 10046 421494 10102
rect 420874 9978 421494 10046
rect 420874 9922 420970 9978
rect 421026 9922 421094 9978
rect 421150 9922 421218 9978
rect 421274 9922 421342 9978
rect 421398 9922 421494 9978
rect 420874 -1120 421494 9922
rect 420874 -1176 420970 -1120
rect 421026 -1176 421094 -1120
rect 421150 -1176 421218 -1120
rect 421274 -1176 421342 -1120
rect 421398 -1176 421494 -1120
rect 420874 -1244 421494 -1176
rect 420874 -1300 420970 -1244
rect 421026 -1300 421094 -1244
rect 421150 -1300 421218 -1244
rect 421274 -1300 421342 -1244
rect 421398 -1300 421494 -1244
rect 420874 -1368 421494 -1300
rect 420874 -1424 420970 -1368
rect 421026 -1424 421094 -1368
rect 421150 -1424 421218 -1368
rect 421274 -1424 421342 -1368
rect 421398 -1424 421494 -1368
rect 420874 -1492 421494 -1424
rect 420874 -1548 420970 -1492
rect 421026 -1548 421094 -1492
rect 421150 -1548 421218 -1492
rect 421274 -1548 421342 -1492
rect 421398 -1548 421494 -1492
rect 420874 -1644 421494 -1548
rect 435154 22350 435774 39922
rect 437612 39284 437668 39294
rect 437612 34804 437668 39228
rect 437612 34738 437668 34748
rect 435154 22294 435250 22350
rect 435306 22294 435374 22350
rect 435430 22294 435498 22350
rect 435554 22294 435622 22350
rect 435678 22294 435774 22350
rect 435154 22226 435774 22294
rect 435154 22170 435250 22226
rect 435306 22170 435374 22226
rect 435430 22170 435498 22226
rect 435554 22170 435622 22226
rect 435678 22170 435774 22226
rect 435154 22102 435774 22170
rect 435154 22046 435250 22102
rect 435306 22046 435374 22102
rect 435430 22046 435498 22102
rect 435554 22046 435622 22102
rect 435678 22046 435774 22102
rect 435154 21978 435774 22046
rect 435154 21922 435250 21978
rect 435306 21922 435374 21978
rect 435430 21922 435498 21978
rect 435554 21922 435622 21978
rect 435678 21922 435774 21978
rect 435154 4350 435774 21922
rect 435154 4294 435250 4350
rect 435306 4294 435374 4350
rect 435430 4294 435498 4350
rect 435554 4294 435622 4350
rect 435678 4294 435774 4350
rect 435154 4226 435774 4294
rect 435154 4170 435250 4226
rect 435306 4170 435374 4226
rect 435430 4170 435498 4226
rect 435554 4170 435622 4226
rect 435678 4170 435774 4226
rect 435154 4102 435774 4170
rect 435154 4046 435250 4102
rect 435306 4046 435374 4102
rect 435430 4046 435498 4102
rect 435554 4046 435622 4102
rect 435678 4046 435774 4102
rect 435154 3978 435774 4046
rect 435154 3922 435250 3978
rect 435306 3922 435374 3978
rect 435430 3922 435498 3978
rect 435554 3922 435622 3978
rect 435678 3922 435774 3978
rect 435154 -160 435774 3922
rect 435154 -216 435250 -160
rect 435306 -216 435374 -160
rect 435430 -216 435498 -160
rect 435554 -216 435622 -160
rect 435678 -216 435774 -160
rect 435154 -284 435774 -216
rect 435154 -340 435250 -284
rect 435306 -340 435374 -284
rect 435430 -340 435498 -284
rect 435554 -340 435622 -284
rect 435678 -340 435774 -284
rect 435154 -408 435774 -340
rect 435154 -464 435250 -408
rect 435306 -464 435374 -408
rect 435430 -464 435498 -408
rect 435554 -464 435622 -408
rect 435678 -464 435774 -408
rect 435154 -532 435774 -464
rect 435154 -588 435250 -532
rect 435306 -588 435374 -532
rect 435430 -588 435498 -532
rect 435554 -588 435622 -532
rect 435678 -588 435774 -532
rect 435154 -1644 435774 -588
rect 438874 28350 439494 41266
rect 453154 40350 453774 41266
rect 453154 40294 453250 40350
rect 453306 40294 453374 40350
rect 453430 40294 453498 40350
rect 453554 40294 453622 40350
rect 453678 40294 453774 40350
rect 453154 40226 453774 40294
rect 453154 40170 453250 40226
rect 453306 40170 453374 40226
rect 453430 40170 453498 40226
rect 453554 40170 453622 40226
rect 453678 40170 453774 40226
rect 453154 40102 453774 40170
rect 453154 40046 453250 40102
rect 453306 40046 453374 40102
rect 453430 40046 453498 40102
rect 453554 40046 453622 40102
rect 453678 40046 453774 40102
rect 453154 39978 453774 40046
rect 453154 39922 453250 39978
rect 453306 39922 453374 39978
rect 453430 39922 453498 39978
rect 453554 39922 453622 39978
rect 453678 39922 453774 39978
rect 451948 39538 452004 39548
rect 451948 39442 452004 39452
rect 438874 28294 438970 28350
rect 439026 28294 439094 28350
rect 439150 28294 439218 28350
rect 439274 28294 439342 28350
rect 439398 28294 439494 28350
rect 438874 28226 439494 28294
rect 438874 28170 438970 28226
rect 439026 28170 439094 28226
rect 439150 28170 439218 28226
rect 439274 28170 439342 28226
rect 439398 28170 439494 28226
rect 438874 28102 439494 28170
rect 438874 28046 438970 28102
rect 439026 28046 439094 28102
rect 439150 28046 439218 28102
rect 439274 28046 439342 28102
rect 439398 28046 439494 28102
rect 438874 27978 439494 28046
rect 438874 27922 438970 27978
rect 439026 27922 439094 27978
rect 439150 27922 439218 27978
rect 439274 27922 439342 27978
rect 439398 27922 439494 27978
rect 438874 10350 439494 27922
rect 438874 10294 438970 10350
rect 439026 10294 439094 10350
rect 439150 10294 439218 10350
rect 439274 10294 439342 10350
rect 439398 10294 439494 10350
rect 438874 10226 439494 10294
rect 438874 10170 438970 10226
rect 439026 10170 439094 10226
rect 439150 10170 439218 10226
rect 439274 10170 439342 10226
rect 439398 10170 439494 10226
rect 438874 10102 439494 10170
rect 438874 10046 438970 10102
rect 439026 10046 439094 10102
rect 439150 10046 439218 10102
rect 439274 10046 439342 10102
rect 439398 10046 439494 10102
rect 438874 9978 439494 10046
rect 438874 9922 438970 9978
rect 439026 9922 439094 9978
rect 439150 9922 439218 9978
rect 439274 9922 439342 9978
rect 439398 9922 439494 9978
rect 438874 -1120 439494 9922
rect 438874 -1176 438970 -1120
rect 439026 -1176 439094 -1120
rect 439150 -1176 439218 -1120
rect 439274 -1176 439342 -1120
rect 439398 -1176 439494 -1120
rect 438874 -1244 439494 -1176
rect 438874 -1300 438970 -1244
rect 439026 -1300 439094 -1244
rect 439150 -1300 439218 -1244
rect 439274 -1300 439342 -1244
rect 439398 -1300 439494 -1244
rect 438874 -1368 439494 -1300
rect 438874 -1424 438970 -1368
rect 439026 -1424 439094 -1368
rect 439150 -1424 439218 -1368
rect 439274 -1424 439342 -1368
rect 439398 -1424 439494 -1368
rect 438874 -1492 439494 -1424
rect 438874 -1548 438970 -1492
rect 439026 -1548 439094 -1492
rect 439150 -1548 439218 -1492
rect 439274 -1548 439342 -1492
rect 439398 -1548 439494 -1492
rect 438874 -1644 439494 -1548
rect 453154 22350 453774 39922
rect 453154 22294 453250 22350
rect 453306 22294 453374 22350
rect 453430 22294 453498 22350
rect 453554 22294 453622 22350
rect 453678 22294 453774 22350
rect 453154 22226 453774 22294
rect 453154 22170 453250 22226
rect 453306 22170 453374 22226
rect 453430 22170 453498 22226
rect 453554 22170 453622 22226
rect 453678 22170 453774 22226
rect 453154 22102 453774 22170
rect 453154 22046 453250 22102
rect 453306 22046 453374 22102
rect 453430 22046 453498 22102
rect 453554 22046 453622 22102
rect 453678 22046 453774 22102
rect 453154 21978 453774 22046
rect 453154 21922 453250 21978
rect 453306 21922 453374 21978
rect 453430 21922 453498 21978
rect 453554 21922 453622 21978
rect 453678 21922 453774 21978
rect 453154 4350 453774 21922
rect 453154 4294 453250 4350
rect 453306 4294 453374 4350
rect 453430 4294 453498 4350
rect 453554 4294 453622 4350
rect 453678 4294 453774 4350
rect 453154 4226 453774 4294
rect 453154 4170 453250 4226
rect 453306 4170 453374 4226
rect 453430 4170 453498 4226
rect 453554 4170 453622 4226
rect 453678 4170 453774 4226
rect 453154 4102 453774 4170
rect 453154 4046 453250 4102
rect 453306 4046 453374 4102
rect 453430 4046 453498 4102
rect 453554 4046 453622 4102
rect 453678 4046 453774 4102
rect 453154 3978 453774 4046
rect 453154 3922 453250 3978
rect 453306 3922 453374 3978
rect 453430 3922 453498 3978
rect 453554 3922 453622 3978
rect 453678 3922 453774 3978
rect 453154 -160 453774 3922
rect 453154 -216 453250 -160
rect 453306 -216 453374 -160
rect 453430 -216 453498 -160
rect 453554 -216 453622 -160
rect 453678 -216 453774 -160
rect 453154 -284 453774 -216
rect 453154 -340 453250 -284
rect 453306 -340 453374 -284
rect 453430 -340 453498 -284
rect 453554 -340 453622 -284
rect 453678 -340 453774 -284
rect 453154 -408 453774 -340
rect 453154 -464 453250 -408
rect 453306 -464 453374 -408
rect 453430 -464 453498 -408
rect 453554 -464 453622 -408
rect 453678 -464 453774 -408
rect 453154 -532 453774 -464
rect 453154 -588 453250 -532
rect 453306 -588 453374 -532
rect 453430 -588 453498 -532
rect 453554 -588 453622 -532
rect 453678 -588 453774 -532
rect 453154 -1644 453774 -588
rect 456874 28350 457494 41266
rect 461132 40404 461188 40414
rect 460012 39396 460068 39406
rect 460012 39292 460068 39302
rect 461132 34692 461188 40348
rect 471154 40350 471774 41266
rect 480172 41188 480228 41198
rect 471154 40294 471250 40350
rect 471306 40294 471374 40350
rect 471430 40294 471498 40350
rect 471554 40294 471622 40350
rect 471678 40294 471774 40350
rect 471154 40226 471774 40294
rect 471154 40170 471250 40226
rect 471306 40170 471374 40226
rect 471430 40170 471498 40226
rect 471554 40170 471622 40226
rect 471678 40170 471774 40226
rect 471154 40102 471774 40170
rect 471154 40046 471250 40102
rect 471306 40046 471374 40102
rect 471430 40046 471498 40102
rect 471554 40046 471622 40102
rect 471678 40046 471774 40102
rect 471154 39978 471774 40046
rect 471154 39922 471250 39978
rect 471306 39922 471374 39978
rect 471430 39922 471498 39978
rect 471554 39922 471622 39978
rect 471678 39922 471774 39978
rect 461132 34626 461188 34636
rect 463708 37380 463764 37390
rect 463708 31798 463764 37324
rect 463708 31732 463764 31742
rect 456874 28294 456970 28350
rect 457026 28294 457094 28350
rect 457150 28294 457218 28350
rect 457274 28294 457342 28350
rect 457398 28294 457494 28350
rect 456874 28226 457494 28294
rect 456874 28170 456970 28226
rect 457026 28170 457094 28226
rect 457150 28170 457218 28226
rect 457274 28170 457342 28226
rect 457398 28170 457494 28226
rect 456874 28102 457494 28170
rect 456874 28046 456970 28102
rect 457026 28046 457094 28102
rect 457150 28046 457218 28102
rect 457274 28046 457342 28102
rect 457398 28046 457494 28102
rect 456874 27978 457494 28046
rect 456874 27922 456970 27978
rect 457026 27922 457094 27978
rect 457150 27922 457218 27978
rect 457274 27922 457342 27978
rect 457398 27922 457494 27978
rect 456874 10350 457494 27922
rect 456874 10294 456970 10350
rect 457026 10294 457094 10350
rect 457150 10294 457218 10350
rect 457274 10294 457342 10350
rect 457398 10294 457494 10350
rect 456874 10226 457494 10294
rect 456874 10170 456970 10226
rect 457026 10170 457094 10226
rect 457150 10170 457218 10226
rect 457274 10170 457342 10226
rect 457398 10170 457494 10226
rect 456874 10102 457494 10170
rect 456874 10046 456970 10102
rect 457026 10046 457094 10102
rect 457150 10046 457218 10102
rect 457274 10046 457342 10102
rect 457398 10046 457494 10102
rect 456874 9978 457494 10046
rect 456874 9922 456970 9978
rect 457026 9922 457094 9978
rect 457150 9922 457218 9978
rect 457274 9922 457342 9978
rect 457398 9922 457494 9978
rect 456874 -1120 457494 9922
rect 456874 -1176 456970 -1120
rect 457026 -1176 457094 -1120
rect 457150 -1176 457218 -1120
rect 457274 -1176 457342 -1120
rect 457398 -1176 457494 -1120
rect 456874 -1244 457494 -1176
rect 456874 -1300 456970 -1244
rect 457026 -1300 457094 -1244
rect 457150 -1300 457218 -1244
rect 457274 -1300 457342 -1244
rect 457398 -1300 457494 -1244
rect 456874 -1368 457494 -1300
rect 456874 -1424 456970 -1368
rect 457026 -1424 457094 -1368
rect 457150 -1424 457218 -1368
rect 457274 -1424 457342 -1368
rect 457398 -1424 457494 -1368
rect 456874 -1492 457494 -1424
rect 456874 -1548 456970 -1492
rect 457026 -1548 457094 -1492
rect 457150 -1548 457218 -1492
rect 457274 -1548 457342 -1492
rect 457398 -1548 457494 -1492
rect 456874 -1644 457494 -1548
rect 471154 22350 471774 39922
rect 471154 22294 471250 22350
rect 471306 22294 471374 22350
rect 471430 22294 471498 22350
rect 471554 22294 471622 22350
rect 471678 22294 471774 22350
rect 471154 22226 471774 22294
rect 471154 22170 471250 22226
rect 471306 22170 471374 22226
rect 471430 22170 471498 22226
rect 471554 22170 471622 22226
rect 471678 22170 471774 22226
rect 471154 22102 471774 22170
rect 471154 22046 471250 22102
rect 471306 22046 471374 22102
rect 471430 22046 471498 22102
rect 471554 22046 471622 22102
rect 471678 22046 471774 22102
rect 471154 21978 471774 22046
rect 471154 21922 471250 21978
rect 471306 21922 471374 21978
rect 471430 21922 471498 21978
rect 471554 21922 471622 21978
rect 471678 21922 471774 21978
rect 471154 4350 471774 21922
rect 471154 4294 471250 4350
rect 471306 4294 471374 4350
rect 471430 4294 471498 4350
rect 471554 4294 471622 4350
rect 471678 4294 471774 4350
rect 471154 4226 471774 4294
rect 471154 4170 471250 4226
rect 471306 4170 471374 4226
rect 471430 4170 471498 4226
rect 471554 4170 471622 4226
rect 471678 4170 471774 4226
rect 471154 4102 471774 4170
rect 471154 4046 471250 4102
rect 471306 4046 471374 4102
rect 471430 4046 471498 4102
rect 471554 4046 471622 4102
rect 471678 4046 471774 4102
rect 471154 3978 471774 4046
rect 471154 3922 471250 3978
rect 471306 3922 471374 3978
rect 471430 3922 471498 3978
rect 471554 3922 471622 3978
rect 471678 3922 471774 3978
rect 471154 -160 471774 3922
rect 471154 -216 471250 -160
rect 471306 -216 471374 -160
rect 471430 -216 471498 -160
rect 471554 -216 471622 -160
rect 471678 -216 471774 -160
rect 471154 -284 471774 -216
rect 471154 -340 471250 -284
rect 471306 -340 471374 -284
rect 471430 -340 471498 -284
rect 471554 -340 471622 -284
rect 471678 -340 471774 -284
rect 471154 -408 471774 -340
rect 471154 -464 471250 -408
rect 471306 -464 471374 -408
rect 471430 -464 471498 -408
rect 471554 -464 471622 -408
rect 471678 -464 471774 -408
rect 471154 -532 471774 -464
rect 471154 -588 471250 -532
rect 471306 -588 471374 -532
rect 471430 -588 471498 -532
rect 471554 -588 471622 -532
rect 471678 -588 471774 -532
rect 471154 -1644 471774 -588
rect 474874 28350 475494 40964
rect 480172 39732 480228 41132
rect 480172 39666 480228 39676
rect 483868 39732 483924 41244
rect 483868 39666 483924 39676
rect 488236 41300 488292 41310
rect 488236 39732 488292 41244
rect 488236 39666 488292 39676
rect 489154 40350 489774 41266
rect 489154 40294 489250 40350
rect 489306 40294 489374 40350
rect 489430 40294 489498 40350
rect 489554 40294 489622 40350
rect 489678 40294 489774 40350
rect 489154 40226 489774 40294
rect 489154 40170 489250 40226
rect 489306 40170 489374 40226
rect 489430 40170 489498 40226
rect 489554 40170 489622 40226
rect 489678 40170 489774 40226
rect 489154 40102 489774 40170
rect 489154 40046 489250 40102
rect 489306 40046 489374 40102
rect 489430 40046 489498 40102
rect 489554 40046 489622 40102
rect 489678 40046 489774 40102
rect 489154 39978 489774 40046
rect 489154 39922 489250 39978
rect 489306 39922 489374 39978
rect 489430 39922 489498 39978
rect 489554 39922 489622 39978
rect 489678 39922 489774 39978
rect 478828 37716 478884 37726
rect 478828 31618 478884 37660
rect 478828 31552 478884 31562
rect 483868 37716 483924 37726
rect 483868 31438 483924 37660
rect 483868 31372 483924 31382
rect 487228 37716 487284 37726
rect 487228 31258 487284 37660
rect 487228 31192 487284 31202
rect 474874 28294 474970 28350
rect 475026 28294 475094 28350
rect 475150 28294 475218 28350
rect 475274 28294 475342 28350
rect 475398 28294 475494 28350
rect 474874 28226 475494 28294
rect 474874 28170 474970 28226
rect 475026 28170 475094 28226
rect 475150 28170 475218 28226
rect 475274 28170 475342 28226
rect 475398 28170 475494 28226
rect 474874 28102 475494 28170
rect 474874 28046 474970 28102
rect 475026 28046 475094 28102
rect 475150 28046 475218 28102
rect 475274 28046 475342 28102
rect 475398 28046 475494 28102
rect 474874 27978 475494 28046
rect 474874 27922 474970 27978
rect 475026 27922 475094 27978
rect 475150 27922 475218 27978
rect 475274 27922 475342 27978
rect 475398 27922 475494 27978
rect 474874 10350 475494 27922
rect 474874 10294 474970 10350
rect 475026 10294 475094 10350
rect 475150 10294 475218 10350
rect 475274 10294 475342 10350
rect 475398 10294 475494 10350
rect 474874 10226 475494 10294
rect 474874 10170 474970 10226
rect 475026 10170 475094 10226
rect 475150 10170 475218 10226
rect 475274 10170 475342 10226
rect 475398 10170 475494 10226
rect 474874 10102 475494 10170
rect 474874 10046 474970 10102
rect 475026 10046 475094 10102
rect 475150 10046 475218 10102
rect 475274 10046 475342 10102
rect 475398 10046 475494 10102
rect 474874 9978 475494 10046
rect 474874 9922 474970 9978
rect 475026 9922 475094 9978
rect 475150 9922 475218 9978
rect 475274 9922 475342 9978
rect 475398 9922 475494 9978
rect 474874 -1120 475494 9922
rect 474874 -1176 474970 -1120
rect 475026 -1176 475094 -1120
rect 475150 -1176 475218 -1120
rect 475274 -1176 475342 -1120
rect 475398 -1176 475494 -1120
rect 474874 -1244 475494 -1176
rect 474874 -1300 474970 -1244
rect 475026 -1300 475094 -1244
rect 475150 -1300 475218 -1244
rect 475274 -1300 475342 -1244
rect 475398 -1300 475494 -1244
rect 474874 -1368 475494 -1300
rect 474874 -1424 474970 -1368
rect 475026 -1424 475094 -1368
rect 475150 -1424 475218 -1368
rect 475274 -1424 475342 -1368
rect 475398 -1424 475494 -1368
rect 474874 -1492 475494 -1424
rect 474874 -1548 474970 -1492
rect 475026 -1548 475094 -1492
rect 475150 -1548 475218 -1492
rect 475274 -1548 475342 -1492
rect 475398 -1548 475494 -1492
rect 474874 -1644 475494 -1548
rect 489154 22350 489774 39922
rect 489154 22294 489250 22350
rect 489306 22294 489374 22350
rect 489430 22294 489498 22350
rect 489554 22294 489622 22350
rect 489678 22294 489774 22350
rect 489154 22226 489774 22294
rect 489154 22170 489250 22226
rect 489306 22170 489374 22226
rect 489430 22170 489498 22226
rect 489554 22170 489622 22226
rect 489678 22170 489774 22226
rect 489154 22102 489774 22170
rect 489154 22046 489250 22102
rect 489306 22046 489374 22102
rect 489430 22046 489498 22102
rect 489554 22046 489622 22102
rect 489678 22046 489774 22102
rect 489154 21978 489774 22046
rect 489154 21922 489250 21978
rect 489306 21922 489374 21978
rect 489430 21922 489498 21978
rect 489554 21922 489622 21978
rect 489678 21922 489774 21978
rect 489154 4350 489774 21922
rect 489154 4294 489250 4350
rect 489306 4294 489374 4350
rect 489430 4294 489498 4350
rect 489554 4294 489622 4350
rect 489678 4294 489774 4350
rect 489154 4226 489774 4294
rect 489154 4170 489250 4226
rect 489306 4170 489374 4226
rect 489430 4170 489498 4226
rect 489554 4170 489622 4226
rect 489678 4170 489774 4226
rect 489154 4102 489774 4170
rect 489154 4046 489250 4102
rect 489306 4046 489374 4102
rect 489430 4046 489498 4102
rect 489554 4046 489622 4102
rect 489678 4046 489774 4102
rect 489154 3978 489774 4046
rect 489154 3922 489250 3978
rect 489306 3922 489374 3978
rect 489430 3922 489498 3978
rect 489554 3922 489622 3978
rect 489678 3922 489774 3978
rect 489154 -160 489774 3922
rect 489154 -216 489250 -160
rect 489306 -216 489374 -160
rect 489430 -216 489498 -160
rect 489554 -216 489622 -160
rect 489678 -216 489774 -160
rect 489154 -284 489774 -216
rect 489154 -340 489250 -284
rect 489306 -340 489374 -284
rect 489430 -340 489498 -284
rect 489554 -340 489622 -284
rect 489678 -340 489774 -284
rect 489154 -408 489774 -340
rect 489154 -464 489250 -408
rect 489306 -464 489374 -408
rect 489430 -464 489498 -408
rect 489554 -464 489622 -408
rect 489678 -464 489774 -408
rect 489154 -532 489774 -464
rect 489154 -588 489250 -532
rect 489306 -588 489374 -532
rect 489430 -588 489498 -532
rect 489554 -588 489622 -532
rect 489678 -588 489774 -532
rect 489154 -1644 489774 -588
rect 492874 28350 493494 41266
rect 496300 39732 496356 41468
rect 496300 39666 496356 39676
rect 507154 40350 507774 41266
rect 507154 40294 507250 40350
rect 507306 40294 507374 40350
rect 507430 40294 507498 40350
rect 507554 40294 507622 40350
rect 507678 40294 507774 40350
rect 507154 40226 507774 40294
rect 507154 40170 507250 40226
rect 507306 40170 507374 40226
rect 507430 40170 507498 40226
rect 507554 40170 507622 40226
rect 507678 40170 507774 40226
rect 507154 40102 507774 40170
rect 507154 40046 507250 40102
rect 507306 40046 507374 40102
rect 507430 40046 507498 40102
rect 507554 40046 507622 40102
rect 507678 40046 507774 40102
rect 507154 39978 507774 40046
rect 507154 39922 507250 39978
rect 507306 39922 507374 39978
rect 507430 39922 507498 39978
rect 507554 39922 507622 39978
rect 507678 39922 507774 39978
rect 500332 37044 500388 37054
rect 500332 29818 500388 36988
rect 504812 37044 504868 37054
rect 504812 31078 504868 36988
rect 504812 31012 504868 31022
rect 500332 29752 500388 29762
rect 492874 28294 492970 28350
rect 493026 28294 493094 28350
rect 493150 28294 493218 28350
rect 493274 28294 493342 28350
rect 493398 28294 493494 28350
rect 492874 28226 493494 28294
rect 492874 28170 492970 28226
rect 493026 28170 493094 28226
rect 493150 28170 493218 28226
rect 493274 28170 493342 28226
rect 493398 28170 493494 28226
rect 492874 28102 493494 28170
rect 492874 28046 492970 28102
rect 493026 28046 493094 28102
rect 493150 28046 493218 28102
rect 493274 28046 493342 28102
rect 493398 28046 493494 28102
rect 492874 27978 493494 28046
rect 492874 27922 492970 27978
rect 493026 27922 493094 27978
rect 493150 27922 493218 27978
rect 493274 27922 493342 27978
rect 493398 27922 493494 27978
rect 492874 10350 493494 27922
rect 492874 10294 492970 10350
rect 493026 10294 493094 10350
rect 493150 10294 493218 10350
rect 493274 10294 493342 10350
rect 493398 10294 493494 10350
rect 492874 10226 493494 10294
rect 492874 10170 492970 10226
rect 493026 10170 493094 10226
rect 493150 10170 493218 10226
rect 493274 10170 493342 10226
rect 493398 10170 493494 10226
rect 492874 10102 493494 10170
rect 492874 10046 492970 10102
rect 493026 10046 493094 10102
rect 493150 10046 493218 10102
rect 493274 10046 493342 10102
rect 493398 10046 493494 10102
rect 492874 9978 493494 10046
rect 492874 9922 492970 9978
rect 493026 9922 493094 9978
rect 493150 9922 493218 9978
rect 493274 9922 493342 9978
rect 493398 9922 493494 9978
rect 492874 -1120 493494 9922
rect 492874 -1176 492970 -1120
rect 493026 -1176 493094 -1120
rect 493150 -1176 493218 -1120
rect 493274 -1176 493342 -1120
rect 493398 -1176 493494 -1120
rect 492874 -1244 493494 -1176
rect 492874 -1300 492970 -1244
rect 493026 -1300 493094 -1244
rect 493150 -1300 493218 -1244
rect 493274 -1300 493342 -1244
rect 493398 -1300 493494 -1244
rect 492874 -1368 493494 -1300
rect 492874 -1424 492970 -1368
rect 493026 -1424 493094 -1368
rect 493150 -1424 493218 -1368
rect 493274 -1424 493342 -1368
rect 493398 -1424 493494 -1368
rect 492874 -1492 493494 -1424
rect 492874 -1548 492970 -1492
rect 493026 -1548 493094 -1492
rect 493150 -1548 493218 -1492
rect 493274 -1548 493342 -1492
rect 493398 -1548 493494 -1492
rect 492874 -1644 493494 -1548
rect 507154 22350 507774 39922
rect 507154 22294 507250 22350
rect 507306 22294 507374 22350
rect 507430 22294 507498 22350
rect 507554 22294 507622 22350
rect 507678 22294 507774 22350
rect 507154 22226 507774 22294
rect 507154 22170 507250 22226
rect 507306 22170 507374 22226
rect 507430 22170 507498 22226
rect 507554 22170 507622 22226
rect 507678 22170 507774 22226
rect 507154 22102 507774 22170
rect 507154 22046 507250 22102
rect 507306 22046 507374 22102
rect 507430 22046 507498 22102
rect 507554 22046 507622 22102
rect 507678 22046 507774 22102
rect 507154 21978 507774 22046
rect 507154 21922 507250 21978
rect 507306 21922 507374 21978
rect 507430 21922 507498 21978
rect 507554 21922 507622 21978
rect 507678 21922 507774 21978
rect 507154 4350 507774 21922
rect 507154 4294 507250 4350
rect 507306 4294 507374 4350
rect 507430 4294 507498 4350
rect 507554 4294 507622 4350
rect 507678 4294 507774 4350
rect 507154 4226 507774 4294
rect 507154 4170 507250 4226
rect 507306 4170 507374 4226
rect 507430 4170 507498 4226
rect 507554 4170 507622 4226
rect 507678 4170 507774 4226
rect 507154 4102 507774 4170
rect 507154 4046 507250 4102
rect 507306 4046 507374 4102
rect 507430 4046 507498 4102
rect 507554 4046 507622 4102
rect 507678 4046 507774 4102
rect 507154 3978 507774 4046
rect 507154 3922 507250 3978
rect 507306 3922 507374 3978
rect 507430 3922 507498 3978
rect 507554 3922 507622 3978
rect 507678 3922 507774 3978
rect 507154 -160 507774 3922
rect 507154 -216 507250 -160
rect 507306 -216 507374 -160
rect 507430 -216 507498 -160
rect 507554 -216 507622 -160
rect 507678 -216 507774 -160
rect 507154 -284 507774 -216
rect 507154 -340 507250 -284
rect 507306 -340 507374 -284
rect 507430 -340 507498 -284
rect 507554 -340 507622 -284
rect 507678 -340 507774 -284
rect 507154 -408 507774 -340
rect 507154 -464 507250 -408
rect 507306 -464 507374 -408
rect 507430 -464 507498 -408
rect 507554 -464 507622 -408
rect 507678 -464 507774 -408
rect 507154 -532 507774 -464
rect 507154 -588 507250 -532
rect 507306 -588 507374 -532
rect 507430 -588 507498 -532
rect 507554 -588 507622 -532
rect 507678 -588 507774 -532
rect 507154 -1644 507774 -588
rect 510874 28350 511494 41266
rect 516460 39732 516516 42902
rect 512428 37044 512484 37054
rect 512428 33238 512484 36988
rect 512428 33172 512484 33182
rect 516460 29998 516516 39676
rect 524972 42902 525364 42958
rect 524524 38612 524580 38622
rect 519148 34580 519204 34590
rect 519148 30178 519204 34524
rect 524524 33058 524580 38556
rect 524972 38612 525028 42902
rect 532700 41518 532756 41528
rect 524972 38546 525028 38556
rect 525154 40350 525774 40964
rect 525154 40294 525250 40350
rect 525306 40294 525374 40350
rect 525430 40294 525498 40350
rect 525554 40294 525622 40350
rect 525678 40294 525774 40350
rect 525154 40226 525774 40294
rect 525154 40170 525250 40226
rect 525306 40170 525374 40226
rect 525430 40170 525498 40226
rect 525554 40170 525622 40226
rect 525678 40170 525774 40226
rect 525154 40102 525774 40170
rect 525154 40046 525250 40102
rect 525306 40046 525374 40102
rect 525430 40046 525498 40102
rect 525554 40046 525622 40102
rect 525678 40046 525774 40102
rect 525154 39978 525774 40046
rect 525154 39922 525250 39978
rect 525306 39922 525374 39978
rect 525430 39922 525498 39978
rect 525554 39922 525622 39978
rect 525678 39922 525774 39978
rect 524524 32992 524580 33002
rect 519148 30112 519204 30122
rect 516460 29932 516516 29942
rect 510874 28294 510970 28350
rect 511026 28294 511094 28350
rect 511150 28294 511218 28350
rect 511274 28294 511342 28350
rect 511398 28294 511494 28350
rect 510874 28226 511494 28294
rect 510874 28170 510970 28226
rect 511026 28170 511094 28226
rect 511150 28170 511218 28226
rect 511274 28170 511342 28226
rect 511398 28170 511494 28226
rect 510874 28102 511494 28170
rect 510874 28046 510970 28102
rect 511026 28046 511094 28102
rect 511150 28046 511218 28102
rect 511274 28046 511342 28102
rect 511398 28046 511494 28102
rect 510874 27978 511494 28046
rect 510874 27922 510970 27978
rect 511026 27922 511094 27978
rect 511150 27922 511218 27978
rect 511274 27922 511342 27978
rect 511398 27922 511494 27978
rect 510874 10350 511494 27922
rect 510874 10294 510970 10350
rect 511026 10294 511094 10350
rect 511150 10294 511218 10350
rect 511274 10294 511342 10350
rect 511398 10294 511494 10350
rect 510874 10226 511494 10294
rect 510874 10170 510970 10226
rect 511026 10170 511094 10226
rect 511150 10170 511218 10226
rect 511274 10170 511342 10226
rect 511398 10170 511494 10226
rect 510874 10102 511494 10170
rect 510874 10046 510970 10102
rect 511026 10046 511094 10102
rect 511150 10046 511218 10102
rect 511274 10046 511342 10102
rect 511398 10046 511494 10102
rect 510874 9978 511494 10046
rect 510874 9922 510970 9978
rect 511026 9922 511094 9978
rect 511150 9922 511218 9978
rect 511274 9922 511342 9978
rect 511398 9922 511494 9978
rect 510874 -1120 511494 9922
rect 510874 -1176 510970 -1120
rect 511026 -1176 511094 -1120
rect 511150 -1176 511218 -1120
rect 511274 -1176 511342 -1120
rect 511398 -1176 511494 -1120
rect 510874 -1244 511494 -1176
rect 510874 -1300 510970 -1244
rect 511026 -1300 511094 -1244
rect 511150 -1300 511218 -1244
rect 511274 -1300 511342 -1244
rect 511398 -1300 511494 -1244
rect 510874 -1368 511494 -1300
rect 510874 -1424 510970 -1368
rect 511026 -1424 511094 -1368
rect 511150 -1424 511218 -1368
rect 511274 -1424 511342 -1368
rect 511398 -1424 511494 -1368
rect 510874 -1492 511494 -1424
rect 510874 -1548 510970 -1492
rect 511026 -1548 511094 -1492
rect 511150 -1548 511218 -1492
rect 511274 -1548 511342 -1492
rect 511398 -1548 511494 -1492
rect 510874 -1644 511494 -1548
rect 525154 22350 525774 39922
rect 528556 37044 528612 37054
rect 528556 34468 528612 36988
rect 528556 32878 528612 34412
rect 528556 32812 528612 32822
rect 525154 22294 525250 22350
rect 525306 22294 525374 22350
rect 525430 22294 525498 22350
rect 525554 22294 525622 22350
rect 525678 22294 525774 22350
rect 525154 22226 525774 22294
rect 525154 22170 525250 22226
rect 525306 22170 525374 22226
rect 525430 22170 525498 22226
rect 525554 22170 525622 22226
rect 525678 22170 525774 22226
rect 525154 22102 525774 22170
rect 525154 22046 525250 22102
rect 525306 22046 525374 22102
rect 525430 22046 525498 22102
rect 525554 22046 525622 22102
rect 525678 22046 525774 22102
rect 525154 21978 525774 22046
rect 525154 21922 525250 21978
rect 525306 21922 525374 21978
rect 525430 21922 525498 21978
rect 525554 21922 525622 21978
rect 525678 21922 525774 21978
rect 525154 4350 525774 21922
rect 525154 4294 525250 4350
rect 525306 4294 525374 4350
rect 525430 4294 525498 4350
rect 525554 4294 525622 4350
rect 525678 4294 525774 4350
rect 525154 4226 525774 4294
rect 525154 4170 525250 4226
rect 525306 4170 525374 4226
rect 525430 4170 525498 4226
rect 525554 4170 525622 4226
rect 525678 4170 525774 4226
rect 525154 4102 525774 4170
rect 525154 4046 525250 4102
rect 525306 4046 525374 4102
rect 525430 4046 525498 4102
rect 525554 4046 525622 4102
rect 525678 4046 525774 4102
rect 525154 3978 525774 4046
rect 525154 3922 525250 3978
rect 525306 3922 525374 3978
rect 525430 3922 525498 3978
rect 525554 3922 525622 3978
rect 525678 3922 525774 3978
rect 525154 -160 525774 3922
rect 525154 -216 525250 -160
rect 525306 -216 525374 -160
rect 525430 -216 525498 -160
rect 525554 -216 525622 -160
rect 525678 -216 525774 -160
rect 525154 -284 525774 -216
rect 525154 -340 525250 -284
rect 525306 -340 525374 -284
rect 525430 -340 525498 -284
rect 525554 -340 525622 -284
rect 525678 -340 525774 -284
rect 525154 -408 525774 -340
rect 525154 -464 525250 -408
rect 525306 -464 525374 -408
rect 525430 -464 525498 -408
rect 525554 -464 525622 -408
rect 525678 -464 525774 -408
rect 525154 -532 525774 -464
rect 525154 -588 525250 -532
rect 525306 -588 525374 -532
rect 525430 -588 525498 -532
rect 525554 -588 525622 -532
rect 525678 -588 525774 -532
rect 525154 -1644 525774 -588
rect 528874 28350 529494 41266
rect 532700 39732 532756 41462
rect 532700 39666 532756 39676
rect 543154 40350 543774 41266
rect 543154 40294 543250 40350
rect 543306 40294 543374 40350
rect 543430 40294 543498 40350
rect 543554 40294 543622 40350
rect 543678 40294 543774 40350
rect 543154 40226 543774 40294
rect 543154 40170 543250 40226
rect 543306 40170 543374 40226
rect 543430 40170 543498 40226
rect 543554 40170 543622 40226
rect 543678 40170 543774 40226
rect 543154 40102 543774 40170
rect 543154 40046 543250 40102
rect 543306 40046 543374 40102
rect 543430 40046 543498 40102
rect 543554 40046 543622 40102
rect 543678 40046 543774 40102
rect 543154 39978 543774 40046
rect 543154 39922 543250 39978
rect 543306 39922 543374 39978
rect 543430 39922 543498 39978
rect 543554 39922 543622 39978
rect 543678 39922 543774 39978
rect 532588 38052 532644 38062
rect 532588 32698 532644 37996
rect 532588 32632 532644 32642
rect 528874 28294 528970 28350
rect 529026 28294 529094 28350
rect 529150 28294 529218 28350
rect 529274 28294 529342 28350
rect 529398 28294 529494 28350
rect 528874 28226 529494 28294
rect 528874 28170 528970 28226
rect 529026 28170 529094 28226
rect 529150 28170 529218 28226
rect 529274 28170 529342 28226
rect 529398 28170 529494 28226
rect 528874 28102 529494 28170
rect 528874 28046 528970 28102
rect 529026 28046 529094 28102
rect 529150 28046 529218 28102
rect 529274 28046 529342 28102
rect 529398 28046 529494 28102
rect 528874 27978 529494 28046
rect 528874 27922 528970 27978
rect 529026 27922 529094 27978
rect 529150 27922 529218 27978
rect 529274 27922 529342 27978
rect 529398 27922 529494 27978
rect 528874 10350 529494 27922
rect 528874 10294 528970 10350
rect 529026 10294 529094 10350
rect 529150 10294 529218 10350
rect 529274 10294 529342 10350
rect 529398 10294 529494 10350
rect 528874 10226 529494 10294
rect 528874 10170 528970 10226
rect 529026 10170 529094 10226
rect 529150 10170 529218 10226
rect 529274 10170 529342 10226
rect 529398 10170 529494 10226
rect 528874 10102 529494 10170
rect 528874 10046 528970 10102
rect 529026 10046 529094 10102
rect 529150 10046 529218 10102
rect 529274 10046 529342 10102
rect 529398 10046 529494 10102
rect 528874 9978 529494 10046
rect 528874 9922 528970 9978
rect 529026 9922 529094 9978
rect 529150 9922 529218 9978
rect 529274 9922 529342 9978
rect 529398 9922 529494 9978
rect 528874 -1120 529494 9922
rect 528874 -1176 528970 -1120
rect 529026 -1176 529094 -1120
rect 529150 -1176 529218 -1120
rect 529274 -1176 529342 -1120
rect 529398 -1176 529494 -1120
rect 528874 -1244 529494 -1176
rect 528874 -1300 528970 -1244
rect 529026 -1300 529094 -1244
rect 529150 -1300 529218 -1244
rect 529274 -1300 529342 -1244
rect 529398 -1300 529494 -1244
rect 528874 -1368 529494 -1300
rect 528874 -1424 528970 -1368
rect 529026 -1424 529094 -1368
rect 529150 -1424 529218 -1368
rect 529274 -1424 529342 -1368
rect 529398 -1424 529494 -1368
rect 528874 -1492 529494 -1424
rect 528874 -1548 528970 -1492
rect 529026 -1548 529094 -1492
rect 529150 -1548 529218 -1492
rect 529274 -1548 529342 -1492
rect 529398 -1548 529494 -1492
rect 528874 -1644 529494 -1548
rect 543154 22350 543774 39922
rect 546028 37940 546084 37956
rect 546028 37852 546084 37862
rect 543154 22294 543250 22350
rect 543306 22294 543374 22350
rect 543430 22294 543498 22350
rect 543554 22294 543622 22350
rect 543678 22294 543774 22350
rect 543154 22226 543774 22294
rect 543154 22170 543250 22226
rect 543306 22170 543374 22226
rect 543430 22170 543498 22226
rect 543554 22170 543622 22226
rect 543678 22170 543774 22226
rect 543154 22102 543774 22170
rect 543154 22046 543250 22102
rect 543306 22046 543374 22102
rect 543430 22046 543498 22102
rect 543554 22046 543622 22102
rect 543678 22046 543774 22102
rect 543154 21978 543774 22046
rect 543154 21922 543250 21978
rect 543306 21922 543374 21978
rect 543430 21922 543498 21978
rect 543554 21922 543622 21978
rect 543678 21922 543774 21978
rect 543154 4350 543774 21922
rect 543154 4294 543250 4350
rect 543306 4294 543374 4350
rect 543430 4294 543498 4350
rect 543554 4294 543622 4350
rect 543678 4294 543774 4350
rect 543154 4226 543774 4294
rect 543154 4170 543250 4226
rect 543306 4170 543374 4226
rect 543430 4170 543498 4226
rect 543554 4170 543622 4226
rect 543678 4170 543774 4226
rect 543154 4102 543774 4170
rect 543154 4046 543250 4102
rect 543306 4046 543374 4102
rect 543430 4046 543498 4102
rect 543554 4046 543622 4102
rect 543678 4046 543774 4102
rect 543154 3978 543774 4046
rect 543154 3922 543250 3978
rect 543306 3922 543374 3978
rect 543430 3922 543498 3978
rect 543554 3922 543622 3978
rect 543678 3922 543774 3978
rect 543154 -160 543774 3922
rect 543154 -216 543250 -160
rect 543306 -216 543374 -160
rect 543430 -216 543498 -160
rect 543554 -216 543622 -160
rect 543678 -216 543774 -160
rect 543154 -284 543774 -216
rect 543154 -340 543250 -284
rect 543306 -340 543374 -284
rect 543430 -340 543498 -284
rect 543554 -340 543622 -284
rect 543678 -340 543774 -284
rect 543154 -408 543774 -340
rect 543154 -464 543250 -408
rect 543306 -464 543374 -408
rect 543430 -464 543498 -408
rect 543554 -464 543622 -408
rect 543678 -464 543774 -408
rect 543154 -532 543774 -464
rect 543154 -588 543250 -532
rect 543306 -588 543374 -532
rect 543430 -588 543498 -532
rect 543554 -588 543622 -532
rect 543678 -588 543774 -532
rect 543154 -1644 543774 -588
rect 546874 28350 547494 41266
rect 546874 28294 546970 28350
rect 547026 28294 547094 28350
rect 547150 28294 547218 28350
rect 547274 28294 547342 28350
rect 547398 28294 547494 28350
rect 546874 28226 547494 28294
rect 546874 28170 546970 28226
rect 547026 28170 547094 28226
rect 547150 28170 547218 28226
rect 547274 28170 547342 28226
rect 547398 28170 547494 28226
rect 546874 28102 547494 28170
rect 546874 28046 546970 28102
rect 547026 28046 547094 28102
rect 547150 28046 547218 28102
rect 547274 28046 547342 28102
rect 547398 28046 547494 28102
rect 546874 27978 547494 28046
rect 546874 27922 546970 27978
rect 547026 27922 547094 27978
rect 547150 27922 547218 27978
rect 547274 27922 547342 27978
rect 547398 27922 547494 27978
rect 546874 10350 547494 27922
rect 548492 21364 548548 54602
rect 548716 54592 548772 54602
rect 548716 51598 548772 51608
rect 548604 49798 548660 49808
rect 548604 23156 548660 49742
rect 548604 23090 548660 23100
rect 548716 21476 548772 51542
rect 548828 38388 548884 55412
rect 548828 38322 548884 38332
rect 548940 42308 548996 42318
rect 548940 21700 548996 42252
rect 548940 21634 548996 21644
rect 548716 21410 548772 21420
rect 548492 21298 548548 21308
rect 546874 10294 546970 10350
rect 547026 10294 547094 10350
rect 547150 10294 547218 10350
rect 547274 10294 547342 10350
rect 547398 10294 547494 10350
rect 546874 10226 547494 10294
rect 546874 10170 546970 10226
rect 547026 10170 547094 10226
rect 547150 10170 547218 10226
rect 547274 10170 547342 10226
rect 547398 10170 547494 10226
rect 546874 10102 547494 10170
rect 546874 10046 546970 10102
rect 547026 10046 547094 10102
rect 547150 10046 547218 10102
rect 547274 10046 547342 10102
rect 547398 10046 547494 10102
rect 546874 9978 547494 10046
rect 546874 9922 546970 9978
rect 547026 9922 547094 9978
rect 547150 9922 547218 9978
rect 547274 9922 547342 9978
rect 547398 9922 547494 9978
rect 546874 -1120 547494 9922
rect 549052 9156 549108 377244
rect 549276 50428 549332 462700
rect 553532 460068 553588 460078
rect 550172 392868 550228 392878
rect 549388 217700 549444 217710
rect 549388 214340 549444 217644
rect 549388 214274 549444 214284
rect 549388 124964 549444 124974
rect 549388 54838 549444 124908
rect 549500 75684 549556 75694
rect 549500 67228 549556 75628
rect 549500 67172 549668 67228
rect 549388 54782 549556 54838
rect 549388 54658 549444 54668
rect 549388 54404 549444 54602
rect 549388 54338 549444 54348
rect 549388 51716 549444 51726
rect 549388 51598 549444 51660
rect 549388 51532 549444 51542
rect 549164 50372 549332 50428
rect 549164 38668 549220 50372
rect 549388 49812 549444 49822
rect 549388 49718 549444 49742
rect 549276 48692 549332 48702
rect 549276 42308 549332 48636
rect 549276 42242 549332 42252
rect 549164 38612 549332 38668
rect 549276 35218 549332 38612
rect 549500 36820 549556 54782
rect 549500 36754 549556 36764
rect 549612 36708 549668 67172
rect 550060 60004 550116 60014
rect 550060 59878 550116 59948
rect 550060 59812 550116 59822
rect 549612 36642 549668 36652
rect 549276 35152 549332 35162
rect 550172 34468 550228 392812
rect 550284 390180 550340 390190
rect 550284 41518 550340 390124
rect 550284 41452 550340 41462
rect 550956 377524 551012 377534
rect 550844 38098 550900 38108
rect 550844 37986 550900 37996
rect 550172 34402 550228 34412
rect 549052 8036 549108 9100
rect 549052 7970 549108 7980
rect 550956 5012 551012 377468
rect 552636 377412 552692 377422
rect 551852 226884 551908 226894
rect 551852 217028 551908 226828
rect 551628 189812 551684 189822
rect 551068 42778 551124 42788
rect 551068 42308 551124 42722
rect 551068 42242 551124 42252
rect 551628 31948 551684 189756
rect 551516 31892 551684 31948
rect 551516 27658 551572 31892
rect 551292 27478 551348 27488
rect 551292 26964 551348 27422
rect 551516 27076 551572 27602
rect 551516 27010 551572 27020
rect 551292 26898 551348 26908
rect 551852 15428 551908 216972
rect 552524 216580 552580 216590
rect 552076 199892 552132 199902
rect 552076 26964 552132 199836
rect 552300 193284 552356 193294
rect 552300 27748 552356 193228
rect 552300 27682 552356 27692
rect 552076 26898 552132 26908
rect 551852 15362 551908 15372
rect 552524 12740 552580 216524
rect 552524 12674 552580 12684
rect 551068 11638 551124 11648
rect 551068 7924 551124 11582
rect 552636 11638 552692 377356
rect 552748 229460 552804 229470
rect 552748 134820 552804 229404
rect 552860 224420 552916 224430
rect 552860 144676 552916 224364
rect 552860 144610 552916 144620
rect 552748 134754 552804 134764
rect 553308 115108 553364 115118
rect 552972 95396 553028 95406
rect 552748 55972 552804 55982
rect 552748 35028 552804 55916
rect 552972 36596 553028 95340
rect 552972 36530 553028 36540
rect 553084 85540 553140 85550
rect 553084 36372 553140 85484
rect 553084 36306 553140 36316
rect 553196 65828 553252 65838
rect 553196 35252 553252 65772
rect 553196 35186 553252 35196
rect 552748 34962 552804 34972
rect 553308 34692 553364 115052
rect 553420 105252 553476 105262
rect 553420 34804 553476 105196
rect 553532 39956 553588 460012
rect 560028 457380 560084 457390
rect 560028 456418 560084 457324
rect 559916 456362 560084 456418
rect 554540 454692 554596 454702
rect 554428 441252 554484 441262
rect 553980 44218 554036 44228
rect 553980 41300 554036 44162
rect 553980 41234 554036 41244
rect 554428 40516 554484 441196
rect 554540 41338 554596 454636
rect 554652 452004 554708 452014
rect 554652 67228 554708 451948
rect 559804 443940 559860 443950
rect 559692 438564 559748 438574
rect 555212 427812 555268 427822
rect 554652 67172 554820 67228
rect 554764 50428 554820 67172
rect 554652 50372 554820 50428
rect 554652 47068 554708 50372
rect 555212 47068 555268 427756
rect 554652 47012 554820 47068
rect 554540 41272 554596 41282
rect 554428 40450 554484 40460
rect 554652 40292 554708 40302
rect 554764 40292 554820 47012
rect 554708 40236 554820 40292
rect 554876 47012 555268 47068
rect 555324 419748 555380 419758
rect 554652 40226 554708 40236
rect 553532 39890 553588 39900
rect 554652 39284 554708 39294
rect 554876 39284 554932 47012
rect 555324 44218 555380 419692
rect 555324 44152 555380 44162
rect 556892 400932 556948 400942
rect 556892 42958 556948 400876
rect 559356 395556 559412 395566
rect 556892 42892 556948 42902
rect 557004 387492 557060 387502
rect 554708 39228 554932 39284
rect 554652 39218 554708 39228
rect 554540 37918 554596 37928
rect 554540 37604 554596 37862
rect 554316 36838 554372 36848
rect 554316 36260 554372 36782
rect 554316 36194 554372 36204
rect 553420 34738 553476 34748
rect 553308 34626 553364 34636
rect 554540 31948 554596 37548
rect 557004 37738 557060 387436
rect 557116 384804 557172 384814
rect 557116 43708 557172 384748
rect 557676 377188 557732 377198
rect 557340 47818 557396 47828
rect 557116 43652 557284 43708
rect 554540 31892 554708 31948
rect 554540 30100 554596 30110
rect 554540 29458 554596 30044
rect 554540 29392 554596 29402
rect 554428 26578 554484 26588
rect 554428 25844 554484 26522
rect 554540 26404 554596 26414
rect 554540 26038 554596 26348
rect 554540 25972 554596 25982
rect 554428 25778 554484 25788
rect 554540 25858 554596 25868
rect 554540 25508 554596 25802
rect 554540 25442 554596 25452
rect 552636 10738 552692 11582
rect 552636 10672 552692 10682
rect 554652 10164 554708 31892
rect 554652 10098 554708 10108
rect 556892 29458 556948 29468
rect 556892 9716 556948 29402
rect 557004 9940 557060 37682
rect 557228 38098 557284 43652
rect 557116 26578 557172 26588
rect 557116 10388 557172 26522
rect 557228 13078 557284 38042
rect 557228 13012 557284 13022
rect 557340 37738 557396 47762
rect 557676 37918 557732 377132
rect 559356 43138 559412 395500
rect 559356 43072 559412 43082
rect 557988 40412 559228 40446
rect 557988 40356 558022 40412
rect 558078 40356 558146 40412
rect 558202 40356 558270 40412
rect 558326 40356 558394 40412
rect 558450 40356 558518 40412
rect 558574 40356 558642 40412
rect 558698 40356 558766 40412
rect 558822 40356 558890 40412
rect 558946 40356 559014 40412
rect 559070 40356 559138 40412
rect 559194 40356 559228 40412
rect 557988 40288 559228 40356
rect 557988 40232 558022 40288
rect 558078 40232 558146 40288
rect 558202 40232 558270 40288
rect 558326 40232 558394 40288
rect 558450 40232 558518 40288
rect 558574 40232 558642 40288
rect 558698 40232 558766 40288
rect 558822 40232 558890 40288
rect 558946 40232 559014 40288
rect 559070 40232 559138 40288
rect 559194 40232 559228 40288
rect 557988 40164 559228 40232
rect 557988 40108 558022 40164
rect 558078 40108 558146 40164
rect 558202 40108 558270 40164
rect 558326 40108 558394 40164
rect 558450 40108 558518 40164
rect 558574 40108 558642 40164
rect 558698 40108 558766 40164
rect 558822 40108 558890 40164
rect 558946 40108 559014 40164
rect 559070 40108 559138 40164
rect 559194 40108 559228 40164
rect 557988 40040 559228 40108
rect 557988 39984 558022 40040
rect 558078 39984 558146 40040
rect 558202 39984 558270 40040
rect 558326 39984 558394 40040
rect 558450 39984 558518 40040
rect 558574 39984 558642 40040
rect 558698 39984 558766 40040
rect 558822 39984 558890 40040
rect 558946 39984 559014 40040
rect 559070 39984 559138 40040
rect 559194 39984 559228 40040
rect 557988 39916 559228 39984
rect 557988 39860 558022 39916
rect 558078 39860 558146 39916
rect 558202 39860 558270 39916
rect 558326 39860 558394 39916
rect 558450 39860 558518 39916
rect 558574 39860 558642 39916
rect 558698 39860 558766 39916
rect 558822 39860 558890 39916
rect 558946 39860 559014 39916
rect 559070 39860 559138 39916
rect 559194 39860 559228 39916
rect 557988 39826 559228 39860
rect 559692 39358 559748 438508
rect 559804 39538 559860 443884
rect 559916 41158 559972 456362
rect 560252 455308 560308 465388
rect 567988 460350 568308 460384
rect 567988 460294 568058 460350
rect 568114 460294 568182 460350
rect 568238 460294 568308 460350
rect 567988 460226 568308 460294
rect 567988 460170 568058 460226
rect 568114 460170 568182 460226
rect 568238 460170 568308 460226
rect 567988 460102 568308 460170
rect 567988 460046 568058 460102
rect 568114 460046 568182 460102
rect 568238 460046 568308 460102
rect 567988 459978 568308 460046
rect 567988 459922 568058 459978
rect 568114 459922 568182 459978
rect 568238 459922 568308 459978
rect 567988 459888 568308 459922
rect 574792 460350 575112 460384
rect 574792 460294 574862 460350
rect 574918 460294 574986 460350
rect 575042 460294 575112 460350
rect 574792 460226 575112 460294
rect 574792 460170 574862 460226
rect 574918 460170 574986 460226
rect 575042 460170 575112 460226
rect 574792 460102 575112 460170
rect 574792 460046 574862 460102
rect 574918 460046 574986 460102
rect 575042 460046 575112 460102
rect 574792 459978 575112 460046
rect 574792 459922 574862 459978
rect 574918 459922 574986 459978
rect 575042 459922 575112 459978
rect 574792 459888 575112 459922
rect 581596 460350 581916 460384
rect 581596 460294 581666 460350
rect 581722 460294 581790 460350
rect 581846 460294 581916 460350
rect 581596 460226 581916 460294
rect 581596 460170 581666 460226
rect 581722 460170 581790 460226
rect 581846 460170 581916 460226
rect 581596 460102 581916 460170
rect 581596 460046 581666 460102
rect 581722 460046 581790 460102
rect 581846 460046 581916 460102
rect 581596 459978 581916 460046
rect 581596 459922 581666 459978
rect 581722 459922 581790 459978
rect 581846 459922 581916 459978
rect 581596 459888 581916 459922
rect 588400 460350 588720 460384
rect 588400 460294 588470 460350
rect 588526 460294 588594 460350
rect 588650 460294 588720 460350
rect 588400 460226 588720 460294
rect 588400 460170 588470 460226
rect 588526 460170 588594 460226
rect 588650 460170 588720 460226
rect 588400 460102 588720 460170
rect 588400 460046 588470 460102
rect 588526 460046 588594 460102
rect 588650 460046 588720 460102
rect 588400 459978 588720 460046
rect 588400 459922 588470 459978
rect 588526 459922 588594 459978
rect 588650 459922 588720 459978
rect 588400 459888 588720 459922
rect 559916 41092 559972 41102
rect 560028 455252 560308 455308
rect 560028 39718 560084 455252
rect 564586 454350 564906 454384
rect 564586 454294 564656 454350
rect 564712 454294 564780 454350
rect 564836 454294 564906 454350
rect 564586 454226 564906 454294
rect 564586 454170 564656 454226
rect 564712 454170 564780 454226
rect 564836 454170 564906 454226
rect 564586 454102 564906 454170
rect 564586 454046 564656 454102
rect 564712 454046 564780 454102
rect 564836 454046 564906 454102
rect 564586 453978 564906 454046
rect 564586 453922 564656 453978
rect 564712 453922 564780 453978
rect 564836 453922 564906 453978
rect 564586 453888 564906 453922
rect 571390 454350 571710 454384
rect 571390 454294 571460 454350
rect 571516 454294 571584 454350
rect 571640 454294 571710 454350
rect 571390 454226 571710 454294
rect 571390 454170 571460 454226
rect 571516 454170 571584 454226
rect 571640 454170 571710 454226
rect 571390 454102 571710 454170
rect 571390 454046 571460 454102
rect 571516 454046 571584 454102
rect 571640 454046 571710 454102
rect 571390 453978 571710 454046
rect 571390 453922 571460 453978
rect 571516 453922 571584 453978
rect 571640 453922 571710 453978
rect 571390 453888 571710 453922
rect 578194 454350 578514 454384
rect 578194 454294 578264 454350
rect 578320 454294 578388 454350
rect 578444 454294 578514 454350
rect 578194 454226 578514 454294
rect 578194 454170 578264 454226
rect 578320 454170 578388 454226
rect 578444 454170 578514 454226
rect 578194 454102 578514 454170
rect 578194 454046 578264 454102
rect 578320 454046 578388 454102
rect 578444 454046 578514 454102
rect 578194 453978 578514 454046
rect 578194 453922 578264 453978
rect 578320 453922 578388 453978
rect 578444 453922 578514 453978
rect 578194 453888 578514 453922
rect 584998 454350 585318 454384
rect 584998 454294 585068 454350
rect 585124 454294 585192 454350
rect 585248 454294 585318 454350
rect 584998 454226 585318 454294
rect 584998 454170 585068 454226
rect 585124 454170 585192 454226
rect 585248 454170 585318 454226
rect 584998 454102 585318 454170
rect 584998 454046 585068 454102
rect 585124 454046 585192 454102
rect 585248 454046 585318 454102
rect 584998 453978 585318 454046
rect 584998 453922 585068 453978
rect 585124 453922 585192 453978
rect 585248 453922 585318 453978
rect 584998 453888 585318 453922
rect 596400 454350 597020 471922
rect 596400 454294 596496 454350
rect 596552 454294 596620 454350
rect 596676 454294 596744 454350
rect 596800 454294 596868 454350
rect 596924 454294 597020 454350
rect 596400 454226 597020 454294
rect 596400 454170 596496 454226
rect 596552 454170 596620 454226
rect 596676 454170 596744 454226
rect 596800 454170 596868 454226
rect 596924 454170 597020 454226
rect 596400 454102 597020 454170
rect 596400 454046 596496 454102
rect 596552 454046 596620 454102
rect 596676 454046 596744 454102
rect 596800 454046 596868 454102
rect 596924 454046 597020 454102
rect 596400 453978 597020 454046
rect 596400 453922 596496 453978
rect 596552 453922 596620 453978
rect 596676 453922 596744 453978
rect 596800 453922 596868 453978
rect 596924 453922 597020 453978
rect 567988 442350 568308 442384
rect 567988 442294 568058 442350
rect 568114 442294 568182 442350
rect 568238 442294 568308 442350
rect 567988 442226 568308 442294
rect 567988 442170 568058 442226
rect 568114 442170 568182 442226
rect 568238 442170 568308 442226
rect 567988 442102 568308 442170
rect 567988 442046 568058 442102
rect 568114 442046 568182 442102
rect 568238 442046 568308 442102
rect 567988 441978 568308 442046
rect 567988 441922 568058 441978
rect 568114 441922 568182 441978
rect 568238 441922 568308 441978
rect 567988 441888 568308 441922
rect 574792 442350 575112 442384
rect 574792 442294 574862 442350
rect 574918 442294 574986 442350
rect 575042 442294 575112 442350
rect 574792 442226 575112 442294
rect 574792 442170 574862 442226
rect 574918 442170 574986 442226
rect 575042 442170 575112 442226
rect 574792 442102 575112 442170
rect 574792 442046 574862 442102
rect 574918 442046 574986 442102
rect 575042 442046 575112 442102
rect 574792 441978 575112 442046
rect 574792 441922 574862 441978
rect 574918 441922 574986 441978
rect 575042 441922 575112 441978
rect 574792 441888 575112 441922
rect 581596 442350 581916 442384
rect 581596 442294 581666 442350
rect 581722 442294 581790 442350
rect 581846 442294 581916 442350
rect 581596 442226 581916 442294
rect 581596 442170 581666 442226
rect 581722 442170 581790 442226
rect 581846 442170 581916 442226
rect 581596 442102 581916 442170
rect 581596 442046 581666 442102
rect 581722 442046 581790 442102
rect 581846 442046 581916 442102
rect 581596 441978 581916 442046
rect 581596 441922 581666 441978
rect 581722 441922 581790 441978
rect 581846 441922 581916 441978
rect 581596 441888 581916 441922
rect 588400 442350 588720 442384
rect 588400 442294 588470 442350
rect 588526 442294 588594 442350
rect 588650 442294 588720 442350
rect 588400 442226 588720 442294
rect 588400 442170 588470 442226
rect 588526 442170 588594 442226
rect 588650 442170 588720 442226
rect 588400 442102 588720 442170
rect 588400 442046 588470 442102
rect 588526 442046 588594 442102
rect 588650 442046 588720 442102
rect 588400 441978 588720 442046
rect 588400 441922 588470 441978
rect 588526 441922 588594 441978
rect 588650 441922 588720 441978
rect 588400 441888 588720 441922
rect 564586 436350 564906 436384
rect 564586 436294 564656 436350
rect 564712 436294 564780 436350
rect 564836 436294 564906 436350
rect 564586 436226 564906 436294
rect 564586 436170 564656 436226
rect 564712 436170 564780 436226
rect 564836 436170 564906 436226
rect 564586 436102 564906 436170
rect 564586 436046 564656 436102
rect 564712 436046 564780 436102
rect 564836 436046 564906 436102
rect 564586 435978 564906 436046
rect 564586 435922 564656 435978
rect 564712 435922 564780 435978
rect 564836 435922 564906 435978
rect 564586 435888 564906 435922
rect 571390 436350 571710 436384
rect 571390 436294 571460 436350
rect 571516 436294 571584 436350
rect 571640 436294 571710 436350
rect 571390 436226 571710 436294
rect 571390 436170 571460 436226
rect 571516 436170 571584 436226
rect 571640 436170 571710 436226
rect 571390 436102 571710 436170
rect 571390 436046 571460 436102
rect 571516 436046 571584 436102
rect 571640 436046 571710 436102
rect 571390 435978 571710 436046
rect 571390 435922 571460 435978
rect 571516 435922 571584 435978
rect 571640 435922 571710 435978
rect 571390 435888 571710 435922
rect 578194 436350 578514 436384
rect 578194 436294 578264 436350
rect 578320 436294 578388 436350
rect 578444 436294 578514 436350
rect 578194 436226 578514 436294
rect 578194 436170 578264 436226
rect 578320 436170 578388 436226
rect 578444 436170 578514 436226
rect 578194 436102 578514 436170
rect 578194 436046 578264 436102
rect 578320 436046 578388 436102
rect 578444 436046 578514 436102
rect 578194 435978 578514 436046
rect 578194 435922 578264 435978
rect 578320 435922 578388 435978
rect 578444 435922 578514 435978
rect 578194 435888 578514 435922
rect 584998 436350 585318 436384
rect 584998 436294 585068 436350
rect 585124 436294 585192 436350
rect 585248 436294 585318 436350
rect 584998 436226 585318 436294
rect 584998 436170 585068 436226
rect 585124 436170 585192 436226
rect 585248 436170 585318 436226
rect 584998 436102 585318 436170
rect 584998 436046 585068 436102
rect 585124 436046 585192 436102
rect 585248 436046 585318 436102
rect 584998 435978 585318 436046
rect 584998 435922 585068 435978
rect 585124 435922 585192 435978
rect 585248 435922 585318 435978
rect 584998 435888 585318 435922
rect 596400 436350 597020 453922
rect 596400 436294 596496 436350
rect 596552 436294 596620 436350
rect 596676 436294 596744 436350
rect 596800 436294 596868 436350
rect 596924 436294 597020 436350
rect 596400 436226 597020 436294
rect 596400 436170 596496 436226
rect 596552 436170 596620 436226
rect 596676 436170 596744 436226
rect 596800 436170 596868 436226
rect 596924 436170 597020 436226
rect 596400 436102 597020 436170
rect 596400 436046 596496 436102
rect 596552 436046 596620 436102
rect 596676 436046 596744 436102
rect 596800 436046 596868 436102
rect 596924 436046 597020 436102
rect 596400 435978 597020 436046
rect 596400 435922 596496 435978
rect 596552 435922 596620 435978
rect 596676 435922 596744 435978
rect 596800 435922 596868 435978
rect 596924 435922 597020 435978
rect 567988 424350 568308 424384
rect 567988 424294 568058 424350
rect 568114 424294 568182 424350
rect 568238 424294 568308 424350
rect 567988 424226 568308 424294
rect 567988 424170 568058 424226
rect 568114 424170 568182 424226
rect 568238 424170 568308 424226
rect 567988 424102 568308 424170
rect 567988 424046 568058 424102
rect 568114 424046 568182 424102
rect 568238 424046 568308 424102
rect 567988 423978 568308 424046
rect 567988 423922 568058 423978
rect 568114 423922 568182 423978
rect 568238 423922 568308 423978
rect 567988 423888 568308 423922
rect 574792 424350 575112 424384
rect 574792 424294 574862 424350
rect 574918 424294 574986 424350
rect 575042 424294 575112 424350
rect 574792 424226 575112 424294
rect 574792 424170 574862 424226
rect 574918 424170 574986 424226
rect 575042 424170 575112 424226
rect 574792 424102 575112 424170
rect 574792 424046 574862 424102
rect 574918 424046 574986 424102
rect 575042 424046 575112 424102
rect 574792 423978 575112 424046
rect 574792 423922 574862 423978
rect 574918 423922 574986 423978
rect 575042 423922 575112 423978
rect 574792 423888 575112 423922
rect 581596 424350 581916 424384
rect 581596 424294 581666 424350
rect 581722 424294 581790 424350
rect 581846 424294 581916 424350
rect 581596 424226 581916 424294
rect 581596 424170 581666 424226
rect 581722 424170 581790 424226
rect 581846 424170 581916 424226
rect 581596 424102 581916 424170
rect 581596 424046 581666 424102
rect 581722 424046 581790 424102
rect 581846 424046 581916 424102
rect 581596 423978 581916 424046
rect 581596 423922 581666 423978
rect 581722 423922 581790 423978
rect 581846 423922 581916 423978
rect 581596 423888 581916 423922
rect 588400 424350 588720 424384
rect 588400 424294 588470 424350
rect 588526 424294 588594 424350
rect 588650 424294 588720 424350
rect 588400 424226 588720 424294
rect 588400 424170 588470 424226
rect 588526 424170 588594 424226
rect 588650 424170 588720 424226
rect 588400 424102 588720 424170
rect 588400 424046 588470 424102
rect 588526 424046 588594 424102
rect 588650 424046 588720 424102
rect 588400 423978 588720 424046
rect 588400 423922 588470 423978
rect 588526 423922 588594 423978
rect 588650 423922 588720 423978
rect 588400 423888 588720 423922
rect 564586 418350 564906 418384
rect 564586 418294 564656 418350
rect 564712 418294 564780 418350
rect 564836 418294 564906 418350
rect 564586 418226 564906 418294
rect 564586 418170 564656 418226
rect 564712 418170 564780 418226
rect 564836 418170 564906 418226
rect 564586 418102 564906 418170
rect 564586 418046 564656 418102
rect 564712 418046 564780 418102
rect 564836 418046 564906 418102
rect 564586 417978 564906 418046
rect 564586 417922 564656 417978
rect 564712 417922 564780 417978
rect 564836 417922 564906 417978
rect 564586 417888 564906 417922
rect 571390 418350 571710 418384
rect 571390 418294 571460 418350
rect 571516 418294 571584 418350
rect 571640 418294 571710 418350
rect 571390 418226 571710 418294
rect 571390 418170 571460 418226
rect 571516 418170 571584 418226
rect 571640 418170 571710 418226
rect 571390 418102 571710 418170
rect 571390 418046 571460 418102
rect 571516 418046 571584 418102
rect 571640 418046 571710 418102
rect 571390 417978 571710 418046
rect 571390 417922 571460 417978
rect 571516 417922 571584 417978
rect 571640 417922 571710 417978
rect 571390 417888 571710 417922
rect 578194 418350 578514 418384
rect 578194 418294 578264 418350
rect 578320 418294 578388 418350
rect 578444 418294 578514 418350
rect 578194 418226 578514 418294
rect 578194 418170 578264 418226
rect 578320 418170 578388 418226
rect 578444 418170 578514 418226
rect 578194 418102 578514 418170
rect 578194 418046 578264 418102
rect 578320 418046 578388 418102
rect 578444 418046 578514 418102
rect 578194 417978 578514 418046
rect 578194 417922 578264 417978
rect 578320 417922 578388 417978
rect 578444 417922 578514 417978
rect 578194 417888 578514 417922
rect 584998 418350 585318 418384
rect 584998 418294 585068 418350
rect 585124 418294 585192 418350
rect 585248 418294 585318 418350
rect 584998 418226 585318 418294
rect 584998 418170 585068 418226
rect 585124 418170 585192 418226
rect 585248 418170 585318 418226
rect 584998 418102 585318 418170
rect 584998 418046 585068 418102
rect 585124 418046 585192 418102
rect 585248 418046 585318 418102
rect 584998 417978 585318 418046
rect 584998 417922 585068 417978
rect 585124 417922 585192 417978
rect 585248 417922 585318 417978
rect 584998 417888 585318 417922
rect 596400 418350 597020 435922
rect 596400 418294 596496 418350
rect 596552 418294 596620 418350
rect 596676 418294 596744 418350
rect 596800 418294 596868 418350
rect 596924 418294 597020 418350
rect 596400 418226 597020 418294
rect 596400 418170 596496 418226
rect 596552 418170 596620 418226
rect 596676 418170 596744 418226
rect 596800 418170 596868 418226
rect 596924 418170 597020 418226
rect 596400 418102 597020 418170
rect 596400 418046 596496 418102
rect 596552 418046 596620 418102
rect 596676 418046 596744 418102
rect 596800 418046 596868 418102
rect 596924 418046 597020 418102
rect 596400 417978 597020 418046
rect 596400 417922 596496 417978
rect 596552 417922 596620 417978
rect 596676 417922 596744 417978
rect 596800 417922 596868 417978
rect 596924 417922 597020 417978
rect 567988 406350 568308 406384
rect 567988 406294 568058 406350
rect 568114 406294 568182 406350
rect 568238 406294 568308 406350
rect 567988 406226 568308 406294
rect 567988 406170 568058 406226
rect 568114 406170 568182 406226
rect 568238 406170 568308 406226
rect 567988 406102 568308 406170
rect 567988 406046 568058 406102
rect 568114 406046 568182 406102
rect 568238 406046 568308 406102
rect 567988 405978 568308 406046
rect 567988 405922 568058 405978
rect 568114 405922 568182 405978
rect 568238 405922 568308 405978
rect 567988 405888 568308 405922
rect 574792 406350 575112 406384
rect 574792 406294 574862 406350
rect 574918 406294 574986 406350
rect 575042 406294 575112 406350
rect 574792 406226 575112 406294
rect 574792 406170 574862 406226
rect 574918 406170 574986 406226
rect 575042 406170 575112 406226
rect 574792 406102 575112 406170
rect 574792 406046 574862 406102
rect 574918 406046 574986 406102
rect 575042 406046 575112 406102
rect 574792 405978 575112 406046
rect 574792 405922 574862 405978
rect 574918 405922 574986 405978
rect 575042 405922 575112 405978
rect 574792 405888 575112 405922
rect 581596 406350 581916 406384
rect 581596 406294 581666 406350
rect 581722 406294 581790 406350
rect 581846 406294 581916 406350
rect 581596 406226 581916 406294
rect 581596 406170 581666 406226
rect 581722 406170 581790 406226
rect 581846 406170 581916 406226
rect 581596 406102 581916 406170
rect 581596 406046 581666 406102
rect 581722 406046 581790 406102
rect 581846 406046 581916 406102
rect 581596 405978 581916 406046
rect 581596 405922 581666 405978
rect 581722 405922 581790 405978
rect 581846 405922 581916 405978
rect 581596 405888 581916 405922
rect 588400 406350 588720 406384
rect 588400 406294 588470 406350
rect 588526 406294 588594 406350
rect 588650 406294 588720 406350
rect 588400 406226 588720 406294
rect 588400 406170 588470 406226
rect 588526 406170 588594 406226
rect 588650 406170 588720 406226
rect 588400 406102 588720 406170
rect 588400 406046 588470 406102
rect 588526 406046 588594 406102
rect 588650 406046 588720 406102
rect 588400 405978 588720 406046
rect 588400 405922 588470 405978
rect 588526 405922 588594 405978
rect 588650 405922 588720 405978
rect 588400 405888 588720 405922
rect 564586 400350 564906 400384
rect 564586 400294 564656 400350
rect 564712 400294 564780 400350
rect 564836 400294 564906 400350
rect 564586 400226 564906 400294
rect 564586 400170 564656 400226
rect 564712 400170 564780 400226
rect 564836 400170 564906 400226
rect 564586 400102 564906 400170
rect 564586 400046 564656 400102
rect 564712 400046 564780 400102
rect 564836 400046 564906 400102
rect 564586 399978 564906 400046
rect 564586 399922 564656 399978
rect 564712 399922 564780 399978
rect 564836 399922 564906 399978
rect 564586 399888 564906 399922
rect 571390 400350 571710 400384
rect 571390 400294 571460 400350
rect 571516 400294 571584 400350
rect 571640 400294 571710 400350
rect 571390 400226 571710 400294
rect 571390 400170 571460 400226
rect 571516 400170 571584 400226
rect 571640 400170 571710 400226
rect 571390 400102 571710 400170
rect 571390 400046 571460 400102
rect 571516 400046 571584 400102
rect 571640 400046 571710 400102
rect 571390 399978 571710 400046
rect 571390 399922 571460 399978
rect 571516 399922 571584 399978
rect 571640 399922 571710 399978
rect 571390 399888 571710 399922
rect 578194 400350 578514 400384
rect 578194 400294 578264 400350
rect 578320 400294 578388 400350
rect 578444 400294 578514 400350
rect 578194 400226 578514 400294
rect 578194 400170 578264 400226
rect 578320 400170 578388 400226
rect 578444 400170 578514 400226
rect 578194 400102 578514 400170
rect 578194 400046 578264 400102
rect 578320 400046 578388 400102
rect 578444 400046 578514 400102
rect 578194 399978 578514 400046
rect 578194 399922 578264 399978
rect 578320 399922 578388 399978
rect 578444 399922 578514 399978
rect 578194 399888 578514 399922
rect 584998 400350 585318 400384
rect 584998 400294 585068 400350
rect 585124 400294 585192 400350
rect 585248 400294 585318 400350
rect 584998 400226 585318 400294
rect 584998 400170 585068 400226
rect 585124 400170 585192 400226
rect 585248 400170 585318 400226
rect 584998 400102 585318 400170
rect 584998 400046 585068 400102
rect 585124 400046 585192 400102
rect 585248 400046 585318 400102
rect 584998 399978 585318 400046
rect 584998 399922 585068 399978
rect 585124 399922 585192 399978
rect 585248 399922 585318 399978
rect 584998 399888 585318 399922
rect 596400 400350 597020 417922
rect 596400 400294 596496 400350
rect 596552 400294 596620 400350
rect 596676 400294 596744 400350
rect 596800 400294 596868 400350
rect 596924 400294 597020 400350
rect 596400 400226 597020 400294
rect 596400 400170 596496 400226
rect 596552 400170 596620 400226
rect 596676 400170 596744 400226
rect 596800 400170 596868 400226
rect 596924 400170 597020 400226
rect 596400 400102 597020 400170
rect 596400 400046 596496 400102
rect 596552 400046 596620 400102
rect 596676 400046 596744 400102
rect 596800 400046 596868 400102
rect 596924 400046 597020 400102
rect 596400 399978 597020 400046
rect 596400 399922 596496 399978
rect 596552 399922 596620 399978
rect 596676 399922 596744 399978
rect 596800 399922 596868 399978
rect 596924 399922 597020 399978
rect 567988 388350 568308 388384
rect 567988 388294 568058 388350
rect 568114 388294 568182 388350
rect 568238 388294 568308 388350
rect 567988 388226 568308 388294
rect 567988 388170 568058 388226
rect 568114 388170 568182 388226
rect 568238 388170 568308 388226
rect 567988 388102 568308 388170
rect 567988 388046 568058 388102
rect 568114 388046 568182 388102
rect 568238 388046 568308 388102
rect 567988 387978 568308 388046
rect 567988 387922 568058 387978
rect 568114 387922 568182 387978
rect 568238 387922 568308 387978
rect 567988 387888 568308 387922
rect 574792 388350 575112 388384
rect 574792 388294 574862 388350
rect 574918 388294 574986 388350
rect 575042 388294 575112 388350
rect 574792 388226 575112 388294
rect 574792 388170 574862 388226
rect 574918 388170 574986 388226
rect 575042 388170 575112 388226
rect 574792 388102 575112 388170
rect 574792 388046 574862 388102
rect 574918 388046 574986 388102
rect 575042 388046 575112 388102
rect 574792 387978 575112 388046
rect 574792 387922 574862 387978
rect 574918 387922 574986 387978
rect 575042 387922 575112 387978
rect 574792 387888 575112 387922
rect 581596 388350 581916 388384
rect 581596 388294 581666 388350
rect 581722 388294 581790 388350
rect 581846 388294 581916 388350
rect 581596 388226 581916 388294
rect 581596 388170 581666 388226
rect 581722 388170 581790 388226
rect 581846 388170 581916 388226
rect 581596 388102 581916 388170
rect 581596 388046 581666 388102
rect 581722 388046 581790 388102
rect 581846 388046 581916 388102
rect 581596 387978 581916 388046
rect 581596 387922 581666 387978
rect 581722 387922 581790 387978
rect 581846 387922 581916 387978
rect 581596 387888 581916 387922
rect 588400 388350 588720 388384
rect 588400 388294 588470 388350
rect 588526 388294 588594 388350
rect 588650 388294 588720 388350
rect 588400 388226 588720 388294
rect 588400 388170 588470 388226
rect 588526 388170 588594 388226
rect 588650 388170 588720 388226
rect 588400 388102 588720 388170
rect 588400 388046 588470 388102
rect 588526 388046 588594 388102
rect 588650 388046 588720 388102
rect 588400 387978 588720 388046
rect 588400 387922 588470 387978
rect 588526 387922 588594 387978
rect 588650 387922 588720 387978
rect 588400 387888 588720 387922
rect 564586 382350 564906 382384
rect 564586 382294 564656 382350
rect 564712 382294 564780 382350
rect 564836 382294 564906 382350
rect 564586 382226 564906 382294
rect 564586 382170 564656 382226
rect 564712 382170 564780 382226
rect 564836 382170 564906 382226
rect 564586 382102 564906 382170
rect 564586 382046 564656 382102
rect 564712 382046 564780 382102
rect 564836 382046 564906 382102
rect 564586 381978 564906 382046
rect 564586 381922 564656 381978
rect 564712 381922 564780 381978
rect 564836 381922 564906 381978
rect 564586 381888 564906 381922
rect 571390 382350 571710 382384
rect 571390 382294 571460 382350
rect 571516 382294 571584 382350
rect 571640 382294 571710 382350
rect 571390 382226 571710 382294
rect 571390 382170 571460 382226
rect 571516 382170 571584 382226
rect 571640 382170 571710 382226
rect 571390 382102 571710 382170
rect 571390 382046 571460 382102
rect 571516 382046 571584 382102
rect 571640 382046 571710 382102
rect 571390 381978 571710 382046
rect 571390 381922 571460 381978
rect 571516 381922 571584 381978
rect 571640 381922 571710 381978
rect 571390 381888 571710 381922
rect 578194 382350 578514 382384
rect 578194 382294 578264 382350
rect 578320 382294 578388 382350
rect 578444 382294 578514 382350
rect 578194 382226 578514 382294
rect 578194 382170 578264 382226
rect 578320 382170 578388 382226
rect 578444 382170 578514 382226
rect 578194 382102 578514 382170
rect 578194 382046 578264 382102
rect 578320 382046 578388 382102
rect 578444 382046 578514 382102
rect 578194 381978 578514 382046
rect 578194 381922 578264 381978
rect 578320 381922 578388 381978
rect 578444 381922 578514 381978
rect 578194 381888 578514 381922
rect 584998 382350 585318 382384
rect 584998 382294 585068 382350
rect 585124 382294 585192 382350
rect 585248 382294 585318 382350
rect 584998 382226 585318 382294
rect 584998 382170 585068 382226
rect 585124 382170 585192 382226
rect 585248 382170 585318 382226
rect 584998 382102 585318 382170
rect 584998 382046 585068 382102
rect 585124 382046 585192 382102
rect 585248 382046 585318 382102
rect 584998 381978 585318 382046
rect 584998 381922 585068 381978
rect 585124 381922 585192 381978
rect 585248 381922 585318 381978
rect 584998 381888 585318 381922
rect 596400 382350 597020 399922
rect 596400 382294 596496 382350
rect 596552 382294 596620 382350
rect 596676 382294 596744 382350
rect 596800 382294 596868 382350
rect 596924 382294 597020 382350
rect 596400 382226 597020 382294
rect 596400 382170 596496 382226
rect 596552 382170 596620 382226
rect 596676 382170 596744 382226
rect 596800 382170 596868 382226
rect 596924 382170 597020 382226
rect 596400 382102 597020 382170
rect 596400 382046 596496 382102
rect 596552 382046 596620 382102
rect 596676 382046 596744 382102
rect 596800 382046 596868 382102
rect 596924 382046 597020 382102
rect 596400 381978 597020 382046
rect 596400 381922 596496 381978
rect 596552 381922 596620 381978
rect 596676 381922 596744 381978
rect 596800 381922 596868 381978
rect 596924 381922 597020 381978
rect 561154 364350 561774 380034
rect 561154 364294 561250 364350
rect 561306 364294 561374 364350
rect 561430 364294 561498 364350
rect 561554 364294 561622 364350
rect 561678 364294 561774 364350
rect 561154 364226 561774 364294
rect 561154 364170 561250 364226
rect 561306 364170 561374 364226
rect 561430 364170 561498 364226
rect 561554 364170 561622 364226
rect 561678 364170 561774 364226
rect 561154 364102 561774 364170
rect 561154 364046 561250 364102
rect 561306 364046 561374 364102
rect 561430 364046 561498 364102
rect 561554 364046 561622 364102
rect 561678 364046 561774 364102
rect 561154 363978 561774 364046
rect 561154 363922 561250 363978
rect 561306 363922 561374 363978
rect 561430 363922 561498 363978
rect 561554 363922 561622 363978
rect 561678 363922 561774 363978
rect 561154 346350 561774 363922
rect 561154 346294 561250 346350
rect 561306 346294 561374 346350
rect 561430 346294 561498 346350
rect 561554 346294 561622 346350
rect 561678 346294 561774 346350
rect 561154 346226 561774 346294
rect 561154 346170 561250 346226
rect 561306 346170 561374 346226
rect 561430 346170 561498 346226
rect 561554 346170 561622 346226
rect 561678 346170 561774 346226
rect 561154 346102 561774 346170
rect 561154 346046 561250 346102
rect 561306 346046 561374 346102
rect 561430 346046 561498 346102
rect 561554 346046 561622 346102
rect 561678 346046 561774 346102
rect 561154 345978 561774 346046
rect 561154 345922 561250 345978
rect 561306 345922 561374 345978
rect 561430 345922 561498 345978
rect 561554 345922 561622 345978
rect 561678 345922 561774 345978
rect 561154 328350 561774 345922
rect 561154 328294 561250 328350
rect 561306 328294 561374 328350
rect 561430 328294 561498 328350
rect 561554 328294 561622 328350
rect 561678 328294 561774 328350
rect 561154 328226 561774 328294
rect 561154 328170 561250 328226
rect 561306 328170 561374 328226
rect 561430 328170 561498 328226
rect 561554 328170 561622 328226
rect 561678 328170 561774 328226
rect 561154 328102 561774 328170
rect 561154 328046 561250 328102
rect 561306 328046 561374 328102
rect 561430 328046 561498 328102
rect 561554 328046 561622 328102
rect 561678 328046 561774 328102
rect 561154 327978 561774 328046
rect 561154 327922 561250 327978
rect 561306 327922 561374 327978
rect 561430 327922 561498 327978
rect 561554 327922 561622 327978
rect 561678 327922 561774 327978
rect 561154 310350 561774 327922
rect 561154 310294 561250 310350
rect 561306 310294 561374 310350
rect 561430 310294 561498 310350
rect 561554 310294 561622 310350
rect 561678 310294 561774 310350
rect 561154 310226 561774 310294
rect 561154 310170 561250 310226
rect 561306 310170 561374 310226
rect 561430 310170 561498 310226
rect 561554 310170 561622 310226
rect 561678 310170 561774 310226
rect 561154 310102 561774 310170
rect 561154 310046 561250 310102
rect 561306 310046 561374 310102
rect 561430 310046 561498 310102
rect 561554 310046 561622 310102
rect 561678 310046 561774 310102
rect 561154 309978 561774 310046
rect 561154 309922 561250 309978
rect 561306 309922 561374 309978
rect 561430 309922 561498 309978
rect 561554 309922 561622 309978
rect 561678 309922 561774 309978
rect 561154 292350 561774 309922
rect 561154 292294 561250 292350
rect 561306 292294 561374 292350
rect 561430 292294 561498 292350
rect 561554 292294 561622 292350
rect 561678 292294 561774 292350
rect 561154 292226 561774 292294
rect 561154 292170 561250 292226
rect 561306 292170 561374 292226
rect 561430 292170 561498 292226
rect 561554 292170 561622 292226
rect 561678 292170 561774 292226
rect 561154 292102 561774 292170
rect 561154 292046 561250 292102
rect 561306 292046 561374 292102
rect 561430 292046 561498 292102
rect 561554 292046 561622 292102
rect 561678 292046 561774 292102
rect 561154 291978 561774 292046
rect 561154 291922 561250 291978
rect 561306 291922 561374 291978
rect 561430 291922 561498 291978
rect 561554 291922 561622 291978
rect 561678 291922 561774 291978
rect 561154 274350 561774 291922
rect 561154 274294 561250 274350
rect 561306 274294 561374 274350
rect 561430 274294 561498 274350
rect 561554 274294 561622 274350
rect 561678 274294 561774 274350
rect 561154 274226 561774 274294
rect 561154 274170 561250 274226
rect 561306 274170 561374 274226
rect 561430 274170 561498 274226
rect 561554 274170 561622 274226
rect 561678 274170 561774 274226
rect 561154 274102 561774 274170
rect 561154 274046 561250 274102
rect 561306 274046 561374 274102
rect 561430 274046 561498 274102
rect 561554 274046 561622 274102
rect 561678 274046 561774 274102
rect 561154 273978 561774 274046
rect 561154 273922 561250 273978
rect 561306 273922 561374 273978
rect 561430 273922 561498 273978
rect 561554 273922 561622 273978
rect 561678 273922 561774 273978
rect 561154 256350 561774 273922
rect 561154 256294 561250 256350
rect 561306 256294 561374 256350
rect 561430 256294 561498 256350
rect 561554 256294 561622 256350
rect 561678 256294 561774 256350
rect 561154 256226 561774 256294
rect 561154 256170 561250 256226
rect 561306 256170 561374 256226
rect 561430 256170 561498 256226
rect 561554 256170 561622 256226
rect 561678 256170 561774 256226
rect 561154 256102 561774 256170
rect 561154 256046 561250 256102
rect 561306 256046 561374 256102
rect 561430 256046 561498 256102
rect 561554 256046 561622 256102
rect 561678 256046 561774 256102
rect 561154 255978 561774 256046
rect 561154 255922 561250 255978
rect 561306 255922 561374 255978
rect 561430 255922 561498 255978
rect 561554 255922 561622 255978
rect 561678 255922 561774 255978
rect 561154 238350 561774 255922
rect 561154 238294 561250 238350
rect 561306 238294 561374 238350
rect 561430 238294 561498 238350
rect 561554 238294 561622 238350
rect 561678 238294 561774 238350
rect 561154 238226 561774 238294
rect 561154 238170 561250 238226
rect 561306 238170 561374 238226
rect 561430 238170 561498 238226
rect 561554 238170 561622 238226
rect 561678 238170 561774 238226
rect 561154 238102 561774 238170
rect 561154 238046 561250 238102
rect 561306 238046 561374 238102
rect 561430 238046 561498 238102
rect 561554 238046 561622 238102
rect 561678 238046 561774 238102
rect 561154 237978 561774 238046
rect 561154 237922 561250 237978
rect 561306 237922 561374 237978
rect 561430 237922 561498 237978
rect 561554 237922 561622 237978
rect 561678 237922 561774 237978
rect 561154 220350 561774 237922
rect 561154 220294 561250 220350
rect 561306 220294 561374 220350
rect 561430 220294 561498 220350
rect 561554 220294 561622 220350
rect 561678 220294 561774 220350
rect 561154 220226 561774 220294
rect 561154 220170 561250 220226
rect 561306 220170 561374 220226
rect 561430 220170 561498 220226
rect 561554 220170 561622 220226
rect 561678 220170 561774 220226
rect 561154 220102 561774 220170
rect 561154 220046 561250 220102
rect 561306 220046 561374 220102
rect 561430 220046 561498 220102
rect 561554 220046 561622 220102
rect 561678 220046 561774 220102
rect 561154 219978 561774 220046
rect 561154 219922 561250 219978
rect 561306 219922 561374 219978
rect 561430 219922 561498 219978
rect 561554 219922 561622 219978
rect 561678 219922 561774 219978
rect 561154 202350 561774 219922
rect 561154 202294 561250 202350
rect 561306 202294 561374 202350
rect 561430 202294 561498 202350
rect 561554 202294 561622 202350
rect 561678 202294 561774 202350
rect 561154 202226 561774 202294
rect 561154 202170 561250 202226
rect 561306 202170 561374 202226
rect 561430 202170 561498 202226
rect 561554 202170 561622 202226
rect 561678 202170 561774 202226
rect 561154 202102 561774 202170
rect 561154 202046 561250 202102
rect 561306 202046 561374 202102
rect 561430 202046 561498 202102
rect 561554 202046 561622 202102
rect 561678 202046 561774 202102
rect 561154 201978 561774 202046
rect 561154 201922 561250 201978
rect 561306 201922 561374 201978
rect 561430 201922 561498 201978
rect 561554 201922 561622 201978
rect 561678 201922 561774 201978
rect 561154 184350 561774 201922
rect 561154 184294 561250 184350
rect 561306 184294 561374 184350
rect 561430 184294 561498 184350
rect 561554 184294 561622 184350
rect 561678 184294 561774 184350
rect 561154 184226 561774 184294
rect 561154 184170 561250 184226
rect 561306 184170 561374 184226
rect 561430 184170 561498 184226
rect 561554 184170 561622 184226
rect 561678 184170 561774 184226
rect 561154 184102 561774 184170
rect 561154 184046 561250 184102
rect 561306 184046 561374 184102
rect 561430 184046 561498 184102
rect 561554 184046 561622 184102
rect 561678 184046 561774 184102
rect 561154 183978 561774 184046
rect 561154 183922 561250 183978
rect 561306 183922 561374 183978
rect 561430 183922 561498 183978
rect 561554 183922 561622 183978
rect 561678 183922 561774 183978
rect 561154 166350 561774 183922
rect 561154 166294 561250 166350
rect 561306 166294 561374 166350
rect 561430 166294 561498 166350
rect 561554 166294 561622 166350
rect 561678 166294 561774 166350
rect 561154 166226 561774 166294
rect 561154 166170 561250 166226
rect 561306 166170 561374 166226
rect 561430 166170 561498 166226
rect 561554 166170 561622 166226
rect 561678 166170 561774 166226
rect 561154 166102 561774 166170
rect 561154 166046 561250 166102
rect 561306 166046 561374 166102
rect 561430 166046 561498 166102
rect 561554 166046 561622 166102
rect 561678 166046 561774 166102
rect 561154 165978 561774 166046
rect 561154 165922 561250 165978
rect 561306 165922 561374 165978
rect 561430 165922 561498 165978
rect 561554 165922 561622 165978
rect 561678 165922 561774 165978
rect 561154 148350 561774 165922
rect 561154 148294 561250 148350
rect 561306 148294 561374 148350
rect 561430 148294 561498 148350
rect 561554 148294 561622 148350
rect 561678 148294 561774 148350
rect 561154 148226 561774 148294
rect 561154 148170 561250 148226
rect 561306 148170 561374 148226
rect 561430 148170 561498 148226
rect 561554 148170 561622 148226
rect 561678 148170 561774 148226
rect 561154 148102 561774 148170
rect 561154 148046 561250 148102
rect 561306 148046 561374 148102
rect 561430 148046 561498 148102
rect 561554 148046 561622 148102
rect 561678 148046 561774 148102
rect 561154 147978 561774 148046
rect 561154 147922 561250 147978
rect 561306 147922 561374 147978
rect 561430 147922 561498 147978
rect 561554 147922 561622 147978
rect 561678 147922 561774 147978
rect 561154 130350 561774 147922
rect 564396 376516 564452 376526
rect 561154 130294 561250 130350
rect 561306 130294 561374 130350
rect 561430 130294 561498 130350
rect 561554 130294 561622 130350
rect 561678 130294 561774 130350
rect 561154 130226 561774 130294
rect 561154 130170 561250 130226
rect 561306 130170 561374 130226
rect 561430 130170 561498 130226
rect 561554 130170 561622 130226
rect 561678 130170 561774 130226
rect 561154 130102 561774 130170
rect 561154 130046 561250 130102
rect 561306 130046 561374 130102
rect 561430 130046 561498 130102
rect 561554 130046 561622 130102
rect 561678 130046 561774 130102
rect 561154 129978 561774 130046
rect 561154 129922 561250 129978
rect 561306 129922 561374 129978
rect 561430 129922 561498 129978
rect 561554 129922 561622 129978
rect 561678 129922 561774 129978
rect 561154 112350 561774 129922
rect 561154 112294 561250 112350
rect 561306 112294 561374 112350
rect 561430 112294 561498 112350
rect 561554 112294 561622 112350
rect 561678 112294 561774 112350
rect 561154 112226 561774 112294
rect 561154 112170 561250 112226
rect 561306 112170 561374 112226
rect 561430 112170 561498 112226
rect 561554 112170 561622 112226
rect 561678 112170 561774 112226
rect 561154 112102 561774 112170
rect 561154 112046 561250 112102
rect 561306 112046 561374 112102
rect 561430 112046 561498 112102
rect 561554 112046 561622 112102
rect 561678 112046 561774 112102
rect 561154 111978 561774 112046
rect 561154 111922 561250 111978
rect 561306 111922 561374 111978
rect 561430 111922 561498 111978
rect 561554 111922 561622 111978
rect 561678 111922 561774 111978
rect 561154 94350 561774 111922
rect 561154 94294 561250 94350
rect 561306 94294 561374 94350
rect 561430 94294 561498 94350
rect 561554 94294 561622 94350
rect 561678 94294 561774 94350
rect 561154 94226 561774 94294
rect 561154 94170 561250 94226
rect 561306 94170 561374 94226
rect 561430 94170 561498 94226
rect 561554 94170 561622 94226
rect 561678 94170 561774 94226
rect 561154 94102 561774 94170
rect 561154 94046 561250 94102
rect 561306 94046 561374 94102
rect 561430 94046 561498 94102
rect 561554 94046 561622 94102
rect 561678 94046 561774 94102
rect 561154 93978 561774 94046
rect 561154 93922 561250 93978
rect 561306 93922 561374 93978
rect 561430 93922 561498 93978
rect 561554 93922 561622 93978
rect 561678 93922 561774 93978
rect 561154 76350 561774 93922
rect 561154 76294 561250 76350
rect 561306 76294 561374 76350
rect 561430 76294 561498 76350
rect 561554 76294 561622 76350
rect 561678 76294 561774 76350
rect 561154 76226 561774 76294
rect 561154 76170 561250 76226
rect 561306 76170 561374 76226
rect 561430 76170 561498 76226
rect 561554 76170 561622 76226
rect 561678 76170 561774 76226
rect 561154 76102 561774 76170
rect 561154 76046 561250 76102
rect 561306 76046 561374 76102
rect 561430 76046 561498 76102
rect 561554 76046 561622 76102
rect 561678 76046 561774 76102
rect 561154 75978 561774 76046
rect 561154 75922 561250 75978
rect 561306 75922 561374 75978
rect 561430 75922 561498 75978
rect 561554 75922 561622 75978
rect 561678 75922 561774 75978
rect 561154 58350 561774 75922
rect 561154 58294 561250 58350
rect 561306 58294 561374 58350
rect 561430 58294 561498 58350
rect 561554 58294 561622 58350
rect 561678 58294 561774 58350
rect 561154 58226 561774 58294
rect 561154 58170 561250 58226
rect 561306 58170 561374 58226
rect 561430 58170 561498 58226
rect 561554 58170 561622 58226
rect 561678 58170 561774 58226
rect 561154 58102 561774 58170
rect 561154 58046 561250 58102
rect 561306 58046 561374 58102
rect 561430 58046 561498 58102
rect 561554 58046 561622 58102
rect 561678 58046 561774 58102
rect 561154 57978 561774 58046
rect 561154 57922 561250 57978
rect 561306 57922 561374 57978
rect 561430 57922 561498 57978
rect 561554 57922 561622 57978
rect 561678 57922 561774 57978
rect 560252 44578 560308 44588
rect 560028 39652 560084 39662
rect 560140 41158 560196 41168
rect 559804 39472 559860 39482
rect 559692 39292 559748 39302
rect 560140 37918 560196 41102
rect 557676 37862 557844 37918
rect 557340 10612 557396 37682
rect 557788 29638 557844 37862
rect 560140 37852 560196 37862
rect 557788 28738 557844 29582
rect 557340 10546 557396 10556
rect 557452 28682 557844 28738
rect 557452 10500 557508 28682
rect 559356 26038 559412 26048
rect 557564 25858 557620 25868
rect 557564 10612 557620 25802
rect 557564 10546 557620 10556
rect 557676 24418 557732 24428
rect 557452 10434 557508 10444
rect 557116 10322 557172 10332
rect 557676 10276 557732 24362
rect 557988 22412 559228 22446
rect 557988 22356 558022 22412
rect 558078 22356 558146 22412
rect 558202 22356 558270 22412
rect 558326 22356 558394 22412
rect 558450 22356 558518 22412
rect 558574 22356 558642 22412
rect 558698 22356 558766 22412
rect 558822 22356 558890 22412
rect 558946 22356 559014 22412
rect 559070 22356 559138 22412
rect 559194 22356 559228 22412
rect 557988 22288 559228 22356
rect 557988 22232 558022 22288
rect 558078 22232 558146 22288
rect 558202 22232 558270 22288
rect 558326 22232 558394 22288
rect 558450 22232 558518 22288
rect 558574 22232 558642 22288
rect 558698 22232 558766 22288
rect 558822 22232 558890 22288
rect 558946 22232 559014 22288
rect 559070 22232 559138 22288
rect 559194 22232 559228 22288
rect 557988 22164 559228 22232
rect 557988 22108 558022 22164
rect 558078 22108 558146 22164
rect 558202 22108 558270 22164
rect 558326 22108 558394 22164
rect 558450 22108 558518 22164
rect 558574 22108 558642 22164
rect 558698 22108 558766 22164
rect 558822 22108 558890 22164
rect 558946 22108 559014 22164
rect 559070 22108 559138 22164
rect 559194 22108 559228 22164
rect 557988 22040 559228 22108
rect 557988 21984 558022 22040
rect 558078 21984 558146 22040
rect 558202 21984 558270 22040
rect 558326 21984 558394 22040
rect 558450 21984 558518 22040
rect 558574 21984 558642 22040
rect 558698 21984 558766 22040
rect 558822 21984 558890 22040
rect 558946 21984 559014 22040
rect 559070 21984 559138 22040
rect 559194 21984 559228 22040
rect 557988 21916 559228 21984
rect 557988 21860 558022 21916
rect 558078 21860 558146 21916
rect 558202 21860 558270 21916
rect 558326 21860 558394 21916
rect 558450 21860 558518 21916
rect 558574 21860 558642 21916
rect 558698 21860 558766 21916
rect 558822 21860 558890 21916
rect 558946 21860 559014 21916
rect 559070 21860 559138 21916
rect 559194 21860 559228 21916
rect 557988 21826 559228 21860
rect 559356 10500 559412 25982
rect 560252 25858 560308 44522
rect 560252 25792 560308 25802
rect 561154 40350 561774 57922
rect 563612 140308 563668 140318
rect 561154 40294 561250 40350
rect 561306 40294 561374 40350
rect 561430 40294 561498 40350
rect 561554 40294 561622 40350
rect 561678 40294 561774 40350
rect 561154 40226 561774 40294
rect 561154 40170 561250 40226
rect 561306 40170 561374 40226
rect 561430 40170 561498 40226
rect 561554 40170 561622 40226
rect 561678 40170 561774 40226
rect 561154 40102 561774 40170
rect 561154 40046 561250 40102
rect 561306 40046 561374 40102
rect 561430 40046 561498 40102
rect 561554 40046 561622 40102
rect 561678 40046 561774 40102
rect 561154 39978 561774 40046
rect 561154 39922 561250 39978
rect 561306 39922 561374 39978
rect 561430 39922 561498 39978
rect 561554 39922 561622 39978
rect 561678 39922 561774 39978
rect 561154 22350 561774 39922
rect 561932 42778 561988 42788
rect 561932 26578 561988 42722
rect 561932 26512 561988 26522
rect 563612 24778 563668 140252
rect 564396 31948 564452 376460
rect 563612 24712 563668 24722
rect 563724 31892 564452 31948
rect 564874 370350 565494 379396
rect 573244 377412 573300 377422
rect 571340 376852 571396 376862
rect 571228 376740 571284 376750
rect 569884 376628 569940 376638
rect 564874 370294 564970 370350
rect 565026 370294 565094 370350
rect 565150 370294 565218 370350
rect 565274 370294 565342 370350
rect 565398 370294 565494 370350
rect 564874 370226 565494 370294
rect 564874 370170 564970 370226
rect 565026 370170 565094 370226
rect 565150 370170 565218 370226
rect 565274 370170 565342 370226
rect 565398 370170 565494 370226
rect 564874 370102 565494 370170
rect 564874 370046 564970 370102
rect 565026 370046 565094 370102
rect 565150 370046 565218 370102
rect 565274 370046 565342 370102
rect 565398 370046 565494 370102
rect 564874 369978 565494 370046
rect 564874 369922 564970 369978
rect 565026 369922 565094 369978
rect 565150 369922 565218 369978
rect 565274 369922 565342 369978
rect 565398 369922 565494 369978
rect 564874 352350 565494 369922
rect 564874 352294 564970 352350
rect 565026 352294 565094 352350
rect 565150 352294 565218 352350
rect 565274 352294 565342 352350
rect 565398 352294 565494 352350
rect 564874 352226 565494 352294
rect 564874 352170 564970 352226
rect 565026 352170 565094 352226
rect 565150 352170 565218 352226
rect 565274 352170 565342 352226
rect 565398 352170 565494 352226
rect 564874 352102 565494 352170
rect 564874 352046 564970 352102
rect 565026 352046 565094 352102
rect 565150 352046 565218 352102
rect 565274 352046 565342 352102
rect 565398 352046 565494 352102
rect 564874 351978 565494 352046
rect 564874 351922 564970 351978
rect 565026 351922 565094 351978
rect 565150 351922 565218 351978
rect 565274 351922 565342 351978
rect 565398 351922 565494 351978
rect 564874 334350 565494 351922
rect 564874 334294 564970 334350
rect 565026 334294 565094 334350
rect 565150 334294 565218 334350
rect 565274 334294 565342 334350
rect 565398 334294 565494 334350
rect 564874 334226 565494 334294
rect 564874 334170 564970 334226
rect 565026 334170 565094 334226
rect 565150 334170 565218 334226
rect 565274 334170 565342 334226
rect 565398 334170 565494 334226
rect 564874 334102 565494 334170
rect 564874 334046 564970 334102
rect 565026 334046 565094 334102
rect 565150 334046 565218 334102
rect 565274 334046 565342 334102
rect 565398 334046 565494 334102
rect 564874 333978 565494 334046
rect 564874 333922 564970 333978
rect 565026 333922 565094 333978
rect 565150 333922 565218 333978
rect 565274 333922 565342 333978
rect 565398 333922 565494 333978
rect 564874 316350 565494 333922
rect 564874 316294 564970 316350
rect 565026 316294 565094 316350
rect 565150 316294 565218 316350
rect 565274 316294 565342 316350
rect 565398 316294 565494 316350
rect 564874 316226 565494 316294
rect 564874 316170 564970 316226
rect 565026 316170 565094 316226
rect 565150 316170 565218 316226
rect 565274 316170 565342 316226
rect 565398 316170 565494 316226
rect 564874 316102 565494 316170
rect 564874 316046 564970 316102
rect 565026 316046 565094 316102
rect 565150 316046 565218 316102
rect 565274 316046 565342 316102
rect 565398 316046 565494 316102
rect 564874 315978 565494 316046
rect 564874 315922 564970 315978
rect 565026 315922 565094 315978
rect 565150 315922 565218 315978
rect 565274 315922 565342 315978
rect 565398 315922 565494 315978
rect 564874 298350 565494 315922
rect 564874 298294 564970 298350
rect 565026 298294 565094 298350
rect 565150 298294 565218 298350
rect 565274 298294 565342 298350
rect 565398 298294 565494 298350
rect 564874 298226 565494 298294
rect 564874 298170 564970 298226
rect 565026 298170 565094 298226
rect 565150 298170 565218 298226
rect 565274 298170 565342 298226
rect 565398 298170 565494 298226
rect 564874 298102 565494 298170
rect 564874 298046 564970 298102
rect 565026 298046 565094 298102
rect 565150 298046 565218 298102
rect 565274 298046 565342 298102
rect 565398 298046 565494 298102
rect 564874 297978 565494 298046
rect 564874 297922 564970 297978
rect 565026 297922 565094 297978
rect 565150 297922 565218 297978
rect 565274 297922 565342 297978
rect 565398 297922 565494 297978
rect 564874 280350 565494 297922
rect 564874 280294 564970 280350
rect 565026 280294 565094 280350
rect 565150 280294 565218 280350
rect 565274 280294 565342 280350
rect 565398 280294 565494 280350
rect 564874 280226 565494 280294
rect 564874 280170 564970 280226
rect 565026 280170 565094 280226
rect 565150 280170 565218 280226
rect 565274 280170 565342 280226
rect 565398 280170 565494 280226
rect 564874 280102 565494 280170
rect 564874 280046 564970 280102
rect 565026 280046 565094 280102
rect 565150 280046 565218 280102
rect 565274 280046 565342 280102
rect 565398 280046 565494 280102
rect 564874 279978 565494 280046
rect 564874 279922 564970 279978
rect 565026 279922 565094 279978
rect 565150 279922 565218 279978
rect 565274 279922 565342 279978
rect 565398 279922 565494 279978
rect 564874 262350 565494 279922
rect 564874 262294 564970 262350
rect 565026 262294 565094 262350
rect 565150 262294 565218 262350
rect 565274 262294 565342 262350
rect 565398 262294 565494 262350
rect 564874 262226 565494 262294
rect 564874 262170 564970 262226
rect 565026 262170 565094 262226
rect 565150 262170 565218 262226
rect 565274 262170 565342 262226
rect 565398 262170 565494 262226
rect 564874 262102 565494 262170
rect 564874 262046 564970 262102
rect 565026 262046 565094 262102
rect 565150 262046 565218 262102
rect 565274 262046 565342 262102
rect 565398 262046 565494 262102
rect 564874 261978 565494 262046
rect 564874 261922 564970 261978
rect 565026 261922 565094 261978
rect 565150 261922 565218 261978
rect 565274 261922 565342 261978
rect 565398 261922 565494 261978
rect 564874 244350 565494 261922
rect 564874 244294 564970 244350
rect 565026 244294 565094 244350
rect 565150 244294 565218 244350
rect 565274 244294 565342 244350
rect 565398 244294 565494 244350
rect 564874 244226 565494 244294
rect 564874 244170 564970 244226
rect 565026 244170 565094 244226
rect 565150 244170 565218 244226
rect 565274 244170 565342 244226
rect 565398 244170 565494 244226
rect 564874 244102 565494 244170
rect 564874 244046 564970 244102
rect 565026 244046 565094 244102
rect 565150 244046 565218 244102
rect 565274 244046 565342 244102
rect 565398 244046 565494 244102
rect 564874 243978 565494 244046
rect 564874 243922 564970 243978
rect 565026 243922 565094 243978
rect 565150 243922 565218 243978
rect 565274 243922 565342 243978
rect 565398 243922 565494 243978
rect 564874 226350 565494 243922
rect 564874 226294 564970 226350
rect 565026 226294 565094 226350
rect 565150 226294 565218 226350
rect 565274 226294 565342 226350
rect 565398 226294 565494 226350
rect 564874 226226 565494 226294
rect 564874 226170 564970 226226
rect 565026 226170 565094 226226
rect 565150 226170 565218 226226
rect 565274 226170 565342 226226
rect 565398 226170 565494 226226
rect 564874 226102 565494 226170
rect 564874 226046 564970 226102
rect 565026 226046 565094 226102
rect 565150 226046 565218 226102
rect 565274 226046 565342 226102
rect 565398 226046 565494 226102
rect 564874 225978 565494 226046
rect 564874 225922 564970 225978
rect 565026 225922 565094 225978
rect 565150 225922 565218 225978
rect 565274 225922 565342 225978
rect 565398 225922 565494 225978
rect 564874 208350 565494 225922
rect 564874 208294 564970 208350
rect 565026 208294 565094 208350
rect 565150 208294 565218 208350
rect 565274 208294 565342 208350
rect 565398 208294 565494 208350
rect 564874 208226 565494 208294
rect 564874 208170 564970 208226
rect 565026 208170 565094 208226
rect 565150 208170 565218 208226
rect 565274 208170 565342 208226
rect 565398 208170 565494 208226
rect 564874 208102 565494 208170
rect 564874 208046 564970 208102
rect 565026 208046 565094 208102
rect 565150 208046 565218 208102
rect 565274 208046 565342 208102
rect 565398 208046 565494 208102
rect 564874 207978 565494 208046
rect 564874 207922 564970 207978
rect 565026 207922 565094 207978
rect 565150 207922 565218 207978
rect 565274 207922 565342 207978
rect 565398 207922 565494 207978
rect 564874 190350 565494 207922
rect 564874 190294 564970 190350
rect 565026 190294 565094 190350
rect 565150 190294 565218 190350
rect 565274 190294 565342 190350
rect 565398 190294 565494 190350
rect 564874 190226 565494 190294
rect 564874 190170 564970 190226
rect 565026 190170 565094 190226
rect 565150 190170 565218 190226
rect 565274 190170 565342 190226
rect 565398 190170 565494 190226
rect 564874 190102 565494 190170
rect 564874 190046 564970 190102
rect 565026 190046 565094 190102
rect 565150 190046 565218 190102
rect 565274 190046 565342 190102
rect 565398 190046 565494 190102
rect 564874 189978 565494 190046
rect 564874 189922 564970 189978
rect 565026 189922 565094 189978
rect 565150 189922 565218 189978
rect 565274 189922 565342 189978
rect 565398 189922 565494 189978
rect 564874 172350 565494 189922
rect 564874 172294 564970 172350
rect 565026 172294 565094 172350
rect 565150 172294 565218 172350
rect 565274 172294 565342 172350
rect 565398 172294 565494 172350
rect 564874 172226 565494 172294
rect 564874 172170 564970 172226
rect 565026 172170 565094 172226
rect 565150 172170 565218 172226
rect 565274 172170 565342 172226
rect 565398 172170 565494 172226
rect 564874 172102 565494 172170
rect 564874 172046 564970 172102
rect 565026 172046 565094 172102
rect 565150 172046 565218 172102
rect 565274 172046 565342 172102
rect 565398 172046 565494 172102
rect 564874 171978 565494 172046
rect 564874 171922 564970 171978
rect 565026 171922 565094 171978
rect 565150 171922 565218 171978
rect 565274 171922 565342 171978
rect 565398 171922 565494 171978
rect 564874 154350 565494 171922
rect 564874 154294 564970 154350
rect 565026 154294 565094 154350
rect 565150 154294 565218 154350
rect 565274 154294 565342 154350
rect 565398 154294 565494 154350
rect 564874 154226 565494 154294
rect 564874 154170 564970 154226
rect 565026 154170 565094 154226
rect 565150 154170 565218 154226
rect 565274 154170 565342 154226
rect 565398 154170 565494 154226
rect 564874 154102 565494 154170
rect 564874 154046 564970 154102
rect 565026 154046 565094 154102
rect 565150 154046 565218 154102
rect 565274 154046 565342 154102
rect 565398 154046 565494 154102
rect 564874 153978 565494 154046
rect 564874 153922 564970 153978
rect 565026 153922 565094 153978
rect 565150 153922 565218 153978
rect 565274 153922 565342 153978
rect 565398 153922 565494 153978
rect 564874 136350 565494 153922
rect 564874 136294 564970 136350
rect 565026 136294 565094 136350
rect 565150 136294 565218 136350
rect 565274 136294 565342 136350
rect 565398 136294 565494 136350
rect 564874 136226 565494 136294
rect 564874 136170 564970 136226
rect 565026 136170 565094 136226
rect 565150 136170 565218 136226
rect 565274 136170 565342 136226
rect 565398 136170 565494 136226
rect 564874 136102 565494 136170
rect 564874 136046 564970 136102
rect 565026 136046 565094 136102
rect 565150 136046 565218 136102
rect 565274 136046 565342 136102
rect 565398 136046 565494 136102
rect 564874 135978 565494 136046
rect 564874 135922 564970 135978
rect 565026 135922 565094 135978
rect 565150 135922 565218 135978
rect 565274 135922 565342 135978
rect 565398 135922 565494 135978
rect 564874 118350 565494 135922
rect 564874 118294 564970 118350
rect 565026 118294 565094 118350
rect 565150 118294 565218 118350
rect 565274 118294 565342 118350
rect 565398 118294 565494 118350
rect 564874 118226 565494 118294
rect 564874 118170 564970 118226
rect 565026 118170 565094 118226
rect 565150 118170 565218 118226
rect 565274 118170 565342 118226
rect 565398 118170 565494 118226
rect 564874 118102 565494 118170
rect 564874 118046 564970 118102
rect 565026 118046 565094 118102
rect 565150 118046 565218 118102
rect 565274 118046 565342 118102
rect 565398 118046 565494 118102
rect 564874 117978 565494 118046
rect 564874 117922 564970 117978
rect 565026 117922 565094 117978
rect 565150 117922 565218 117978
rect 565274 117922 565342 117978
rect 565398 117922 565494 117978
rect 564874 100350 565494 117922
rect 564874 100294 564970 100350
rect 565026 100294 565094 100350
rect 565150 100294 565218 100350
rect 565274 100294 565342 100350
rect 565398 100294 565494 100350
rect 564874 100226 565494 100294
rect 564874 100170 564970 100226
rect 565026 100170 565094 100226
rect 565150 100170 565218 100226
rect 565274 100170 565342 100226
rect 565398 100170 565494 100226
rect 564874 100102 565494 100170
rect 564874 100046 564970 100102
rect 565026 100046 565094 100102
rect 565150 100046 565218 100102
rect 565274 100046 565342 100102
rect 565398 100046 565494 100102
rect 564874 99978 565494 100046
rect 564874 99922 564970 99978
rect 565026 99922 565094 99978
rect 565150 99922 565218 99978
rect 565274 99922 565342 99978
rect 565398 99922 565494 99978
rect 564874 82350 565494 99922
rect 564874 82294 564970 82350
rect 565026 82294 565094 82350
rect 565150 82294 565218 82350
rect 565274 82294 565342 82350
rect 565398 82294 565494 82350
rect 564874 82226 565494 82294
rect 564874 82170 564970 82226
rect 565026 82170 565094 82226
rect 565150 82170 565218 82226
rect 565274 82170 565342 82226
rect 565398 82170 565494 82226
rect 564874 82102 565494 82170
rect 564874 82046 564970 82102
rect 565026 82046 565094 82102
rect 565150 82046 565218 82102
rect 565274 82046 565342 82102
rect 565398 82046 565494 82102
rect 564874 81978 565494 82046
rect 564874 81922 564970 81978
rect 565026 81922 565094 81978
rect 565150 81922 565218 81978
rect 565274 81922 565342 81978
rect 565398 81922 565494 81978
rect 564874 64350 565494 81922
rect 564874 64294 564970 64350
rect 565026 64294 565094 64350
rect 565150 64294 565218 64350
rect 565274 64294 565342 64350
rect 565398 64294 565494 64350
rect 564874 64226 565494 64294
rect 564874 64170 564970 64226
rect 565026 64170 565094 64226
rect 565150 64170 565218 64226
rect 565274 64170 565342 64226
rect 565398 64170 565494 64226
rect 564874 64102 565494 64170
rect 564874 64046 564970 64102
rect 565026 64046 565094 64102
rect 565150 64046 565218 64102
rect 565274 64046 565342 64102
rect 565398 64046 565494 64102
rect 564874 63978 565494 64046
rect 564874 63922 564970 63978
rect 565026 63922 565094 63978
rect 565150 63922 565218 63978
rect 565274 63922 565342 63978
rect 565398 63922 565494 63978
rect 564874 46350 565494 63922
rect 564874 46294 564970 46350
rect 565026 46294 565094 46350
rect 565150 46294 565218 46350
rect 565274 46294 565342 46350
rect 565398 46294 565494 46350
rect 564874 46226 565494 46294
rect 564874 46170 564970 46226
rect 565026 46170 565094 46226
rect 565150 46170 565218 46226
rect 565274 46170 565342 46226
rect 565398 46170 565494 46226
rect 564874 46102 565494 46170
rect 564874 46046 564970 46102
rect 565026 46046 565094 46102
rect 565150 46046 565218 46102
rect 565274 46046 565342 46102
rect 565398 46046 565494 46102
rect 564874 45978 565494 46046
rect 564874 45922 564970 45978
rect 565026 45922 565094 45978
rect 565150 45922 565218 45978
rect 565274 45922 565342 45978
rect 565398 45922 565494 45978
rect 563724 25318 563780 31892
rect 561154 22294 561250 22350
rect 561306 22294 561374 22350
rect 561430 22294 561498 22350
rect 561554 22294 561622 22350
rect 561678 22294 561774 22350
rect 561154 22226 561774 22294
rect 561154 22170 561250 22226
rect 561306 22170 561374 22226
rect 561430 22170 561498 22226
rect 561554 22170 561622 22226
rect 561678 22170 561774 22226
rect 561154 22102 561774 22170
rect 561154 22046 561250 22102
rect 561306 22046 561374 22102
rect 561430 22046 561498 22102
rect 561554 22046 561622 22102
rect 561678 22046 561774 22102
rect 561154 21978 561774 22046
rect 561154 21922 561250 21978
rect 561306 21922 561374 21978
rect 561430 21922 561498 21978
rect 561554 21922 561622 21978
rect 561678 21922 561774 21978
rect 561154 20830 561774 21922
rect 563724 20098 563780 25262
rect 564874 28350 565494 45922
rect 566972 375620 567028 375630
rect 565740 38638 565796 38648
rect 564874 28294 564970 28350
rect 565026 28294 565094 28350
rect 565150 28294 565218 28350
rect 565274 28294 565342 28350
rect 565398 28294 565494 28350
rect 564874 28226 565494 28294
rect 564874 28170 564970 28226
rect 565026 28170 565094 28226
rect 565150 28170 565218 28226
rect 565274 28170 565342 28226
rect 565398 28170 565494 28226
rect 564874 28102 565494 28170
rect 564874 28046 564970 28102
rect 565026 28046 565094 28102
rect 565150 28046 565218 28102
rect 565274 28046 565342 28102
rect 565398 28046 565494 28102
rect 564874 27978 565494 28046
rect 564874 27922 564970 27978
rect 565026 27922 565094 27978
rect 565150 27922 565218 27978
rect 565274 27922 565342 27978
rect 565398 27922 565494 27978
rect 564874 20830 565494 27922
rect 565628 37738 565684 37748
rect 565628 26038 565684 37682
rect 565740 29458 565796 38582
rect 566972 36838 567028 375564
rect 567988 46412 569228 46446
rect 567988 46356 568022 46412
rect 568078 46356 568146 46412
rect 568202 46356 568270 46412
rect 568326 46356 568394 46412
rect 568450 46356 568518 46412
rect 568574 46356 568642 46412
rect 568698 46356 568766 46412
rect 568822 46356 568890 46412
rect 568946 46356 569014 46412
rect 569070 46356 569138 46412
rect 569194 46356 569228 46412
rect 567988 46288 569228 46356
rect 567988 46232 568022 46288
rect 568078 46232 568146 46288
rect 568202 46232 568270 46288
rect 568326 46232 568394 46288
rect 568450 46232 568518 46288
rect 568574 46232 568642 46288
rect 568698 46232 568766 46288
rect 568822 46232 568890 46288
rect 568946 46232 569014 46288
rect 569070 46232 569138 46288
rect 569194 46232 569228 46288
rect 567988 46164 569228 46232
rect 567988 46108 568022 46164
rect 568078 46108 568146 46164
rect 568202 46108 568270 46164
rect 568326 46108 568394 46164
rect 568450 46108 568518 46164
rect 568574 46108 568642 46164
rect 568698 46108 568766 46164
rect 568822 46108 568890 46164
rect 568946 46108 569014 46164
rect 569070 46108 569138 46164
rect 569194 46108 569228 46164
rect 567988 46040 569228 46108
rect 567988 45984 568022 46040
rect 568078 45984 568146 46040
rect 568202 45984 568270 46040
rect 568326 45984 568394 46040
rect 568450 45984 568518 46040
rect 568574 45984 568642 46040
rect 568698 45984 568766 46040
rect 568822 45984 568890 46040
rect 568946 45984 569014 46040
rect 569070 45984 569138 46040
rect 569194 45984 569228 46040
rect 567988 45916 569228 45984
rect 567988 45860 568022 45916
rect 568078 45860 568146 45916
rect 568202 45860 568270 45916
rect 568326 45860 568394 45916
rect 568450 45860 568518 45916
rect 568574 45860 568642 45916
rect 568698 45860 568766 45916
rect 568822 45860 568890 45916
rect 568946 45860 569014 45916
rect 569070 45860 569138 45916
rect 569194 45860 569228 45916
rect 567988 45826 569228 45860
rect 566972 36772 567028 36782
rect 567756 42958 567812 42968
rect 565740 29392 565796 29402
rect 565628 25972 565684 25982
rect 567756 24958 567812 42902
rect 567988 28412 569228 28446
rect 567988 28356 568022 28412
rect 568078 28356 568146 28412
rect 568202 28356 568270 28412
rect 568326 28356 568394 28412
rect 568450 28356 568518 28412
rect 568574 28356 568642 28412
rect 568698 28356 568766 28412
rect 568822 28356 568890 28412
rect 568946 28356 569014 28412
rect 569070 28356 569138 28412
rect 569194 28356 569228 28412
rect 567988 28288 569228 28356
rect 567988 28232 568022 28288
rect 568078 28232 568146 28288
rect 568202 28232 568270 28288
rect 568326 28232 568394 28288
rect 568450 28232 568518 28288
rect 568574 28232 568642 28288
rect 568698 28232 568766 28288
rect 568822 28232 568890 28288
rect 568946 28232 569014 28288
rect 569070 28232 569138 28288
rect 569194 28232 569228 28288
rect 567988 28164 569228 28232
rect 567988 28108 568022 28164
rect 568078 28108 568146 28164
rect 568202 28108 568270 28164
rect 568326 28108 568394 28164
rect 568450 28108 568518 28164
rect 568574 28108 568642 28164
rect 568698 28108 568766 28164
rect 568822 28108 568890 28164
rect 568946 28108 569014 28164
rect 569070 28108 569138 28164
rect 569194 28108 569228 28164
rect 567988 28040 569228 28108
rect 567988 27984 568022 28040
rect 568078 27984 568146 28040
rect 568202 27984 568270 28040
rect 568326 27984 568394 28040
rect 568450 27984 568518 28040
rect 568574 27984 568642 28040
rect 568698 27984 568766 28040
rect 568822 27984 568890 28040
rect 568946 27984 569014 28040
rect 569070 27984 569138 28040
rect 569194 27984 569228 28040
rect 567988 27916 569228 27984
rect 567988 27860 568022 27916
rect 568078 27860 568146 27916
rect 568202 27860 568270 27916
rect 568326 27860 568394 27916
rect 568450 27860 568518 27916
rect 568574 27860 568642 27916
rect 568698 27860 568766 27916
rect 568822 27860 568890 27916
rect 568946 27860 569014 27916
rect 569070 27860 569138 27916
rect 569194 27860 569228 27916
rect 567988 27826 569228 27860
rect 567756 24892 567812 24902
rect 563724 20032 563780 20042
rect 559356 10434 559412 10444
rect 560028 13078 560084 13088
rect 557676 10210 557732 10220
rect 558012 10388 558068 10398
rect 558012 10164 558068 10332
rect 560028 10388 560084 13022
rect 560028 10322 560084 10332
rect 558012 10098 558068 10108
rect 557004 9874 557060 9884
rect 556892 9650 556948 9660
rect 551068 7858 551124 7868
rect 550956 4946 551012 4956
rect 546874 -1176 546970 -1120
rect 547026 -1176 547094 -1120
rect 547150 -1176 547218 -1120
rect 547274 -1176 547342 -1120
rect 547398 -1176 547494 -1120
rect 546874 -1244 547494 -1176
rect 546874 -1300 546970 -1244
rect 547026 -1300 547094 -1244
rect 547150 -1300 547218 -1244
rect 547274 -1300 547342 -1244
rect 547398 -1300 547494 -1244
rect 546874 -1368 547494 -1300
rect 546874 -1424 546970 -1368
rect 547026 -1424 547094 -1368
rect 547150 -1424 547218 -1368
rect 547274 -1424 547342 -1368
rect 547398 -1424 547494 -1368
rect 546874 -1492 547494 -1424
rect 546874 -1548 546970 -1492
rect 547026 -1548 547094 -1492
rect 547150 -1548 547218 -1492
rect 547274 -1548 547342 -1492
rect 547398 -1548 547494 -1492
rect 546874 -1644 547494 -1548
rect 561154 4350 561774 11154
rect 561154 4294 561250 4350
rect 561306 4294 561374 4350
rect 561430 4294 561498 4350
rect 561554 4294 561622 4350
rect 561678 4294 561774 4350
rect 561154 4226 561774 4294
rect 561154 4170 561250 4226
rect 561306 4170 561374 4226
rect 561430 4170 561498 4226
rect 561554 4170 561622 4226
rect 561678 4170 561774 4226
rect 561154 4102 561774 4170
rect 561154 4046 561250 4102
rect 561306 4046 561374 4102
rect 561430 4046 561498 4102
rect 561554 4046 561622 4102
rect 561678 4046 561774 4102
rect 561154 3978 561774 4046
rect 561154 3922 561250 3978
rect 561306 3922 561374 3978
rect 561430 3922 561498 3978
rect 561554 3922 561622 3978
rect 561678 3922 561774 3978
rect 561154 -160 561774 3922
rect 561154 -216 561250 -160
rect 561306 -216 561374 -160
rect 561430 -216 561498 -160
rect 561554 -216 561622 -160
rect 561678 -216 561774 -160
rect 561154 -284 561774 -216
rect 561154 -340 561250 -284
rect 561306 -340 561374 -284
rect 561430 -340 561498 -284
rect 561554 -340 561622 -284
rect 561678 -340 561774 -284
rect 561154 -408 561774 -340
rect 561154 -464 561250 -408
rect 561306 -464 561374 -408
rect 561430 -464 561498 -408
rect 561554 -464 561622 -408
rect 561678 -464 561774 -408
rect 561154 -532 561774 -464
rect 561154 -588 561250 -532
rect 561306 -588 561374 -532
rect 561430 -588 561498 -532
rect 561554 -588 561622 -532
rect 561678 -588 561774 -532
rect 561154 -1644 561774 -588
rect 564874 10350 565494 11154
rect 564874 10294 564970 10350
rect 565026 10294 565094 10350
rect 565150 10294 565218 10350
rect 565274 10294 565342 10350
rect 565398 10294 565494 10350
rect 564874 10226 565494 10294
rect 564874 10170 564970 10226
rect 565026 10170 565094 10226
rect 565150 10170 565218 10226
rect 565274 10170 565342 10226
rect 565398 10170 565494 10226
rect 564874 10102 565494 10170
rect 564874 10046 564970 10102
rect 565026 10046 565094 10102
rect 565150 10046 565218 10102
rect 565274 10046 565342 10102
rect 565398 10046 565494 10102
rect 564874 9978 565494 10046
rect 564874 9922 564970 9978
rect 565026 9922 565094 9978
rect 565150 9922 565218 9978
rect 565274 9922 565342 9978
rect 565398 9922 565494 9978
rect 564874 -1120 565494 9922
rect 569884 7700 569940 376572
rect 571116 376628 571172 376638
rect 569884 7634 569940 7644
rect 569996 376516 570052 376526
rect 569996 8036 570052 376460
rect 571004 376516 571060 376526
rect 570108 24958 570164 24968
rect 570108 9940 570164 24902
rect 570108 9874 570164 9884
rect 569996 7028 570052 7980
rect 569996 6962 570052 6972
rect 571004 7498 571060 376460
rect 571004 308 571060 7442
rect 571116 7924 571172 376572
rect 571116 6244 571172 7868
rect 571228 8148 571284 376684
rect 571228 6804 571284 8092
rect 571340 7700 571396 376796
rect 572684 376628 572740 376638
rect 571340 7252 571396 7644
rect 571340 7186 571396 7196
rect 572572 376516 572628 376526
rect 572572 7858 572628 376460
rect 571228 6738 571284 6748
rect 571116 6178 571172 6188
rect 571004 242 571060 252
rect 572572 84 572628 7802
rect 572684 7678 572740 376572
rect 572684 196 572740 7622
rect 572796 376516 572852 376526
rect 572796 8038 572852 376460
rect 572908 37018 572964 37028
rect 572908 8372 572964 36962
rect 572908 8306 572964 8316
rect 572796 6132 572852 7982
rect 573244 7140 573300 377356
rect 574812 377300 574868 377310
rect 574364 376628 574420 376638
rect 573692 376292 573748 376302
rect 573692 38638 573748 376236
rect 573692 38572 573748 38582
rect 573244 7074 573300 7084
rect 574364 10500 574420 376572
rect 574588 376628 574644 376638
rect 574476 376516 574532 376526
rect 574476 10612 574532 376460
rect 574476 10546 574532 10556
rect 572796 6066 572852 6076
rect 574364 6020 574420 10444
rect 574588 9604 574644 376572
rect 574588 9538 574644 9548
rect 574812 8428 574868 377244
rect 577052 376740 577108 376750
rect 576268 376516 576324 376526
rect 575372 376404 575428 376414
rect 575372 9940 575428 376348
rect 575372 9874 575428 9884
rect 576268 9380 576324 376460
rect 577052 42958 577108 376684
rect 577948 376516 578004 376526
rect 577948 56998 578004 376460
rect 579154 364350 579774 380034
rect 579964 376964 580020 376974
rect 579154 364294 579250 364350
rect 579306 364294 579374 364350
rect 579430 364294 579498 364350
rect 579554 364294 579622 364350
rect 579678 364294 579774 364350
rect 579154 364226 579774 364294
rect 579154 364170 579250 364226
rect 579306 364170 579374 364226
rect 579430 364170 579498 364226
rect 579554 364170 579622 364226
rect 579678 364170 579774 364226
rect 579154 364102 579774 364170
rect 579154 364046 579250 364102
rect 579306 364046 579374 364102
rect 579430 364046 579498 364102
rect 579554 364046 579622 364102
rect 579678 364046 579774 364102
rect 579154 363978 579774 364046
rect 579154 363922 579250 363978
rect 579306 363922 579374 363978
rect 579430 363922 579498 363978
rect 579554 363922 579622 363978
rect 579678 363922 579774 363978
rect 579154 346350 579774 363922
rect 579154 346294 579250 346350
rect 579306 346294 579374 346350
rect 579430 346294 579498 346350
rect 579554 346294 579622 346350
rect 579678 346294 579774 346350
rect 579154 346226 579774 346294
rect 579154 346170 579250 346226
rect 579306 346170 579374 346226
rect 579430 346170 579498 346226
rect 579554 346170 579622 346226
rect 579678 346170 579774 346226
rect 579154 346102 579774 346170
rect 579154 346046 579250 346102
rect 579306 346046 579374 346102
rect 579430 346046 579498 346102
rect 579554 346046 579622 346102
rect 579678 346046 579774 346102
rect 579154 345978 579774 346046
rect 579154 345922 579250 345978
rect 579306 345922 579374 345978
rect 579430 345922 579498 345978
rect 579554 345922 579622 345978
rect 579678 345922 579774 345978
rect 579154 328350 579774 345922
rect 579154 328294 579250 328350
rect 579306 328294 579374 328350
rect 579430 328294 579498 328350
rect 579554 328294 579622 328350
rect 579678 328294 579774 328350
rect 579154 328226 579774 328294
rect 579154 328170 579250 328226
rect 579306 328170 579374 328226
rect 579430 328170 579498 328226
rect 579554 328170 579622 328226
rect 579678 328170 579774 328226
rect 579154 328102 579774 328170
rect 579154 328046 579250 328102
rect 579306 328046 579374 328102
rect 579430 328046 579498 328102
rect 579554 328046 579622 328102
rect 579678 328046 579774 328102
rect 579154 327978 579774 328046
rect 579154 327922 579250 327978
rect 579306 327922 579374 327978
rect 579430 327922 579498 327978
rect 579554 327922 579622 327978
rect 579678 327922 579774 327978
rect 579154 310350 579774 327922
rect 579154 310294 579250 310350
rect 579306 310294 579374 310350
rect 579430 310294 579498 310350
rect 579554 310294 579622 310350
rect 579678 310294 579774 310350
rect 579154 310226 579774 310294
rect 579154 310170 579250 310226
rect 579306 310170 579374 310226
rect 579430 310170 579498 310226
rect 579554 310170 579622 310226
rect 579678 310170 579774 310226
rect 579154 310102 579774 310170
rect 579154 310046 579250 310102
rect 579306 310046 579374 310102
rect 579430 310046 579498 310102
rect 579554 310046 579622 310102
rect 579678 310046 579774 310102
rect 579154 309978 579774 310046
rect 579154 309922 579250 309978
rect 579306 309922 579374 309978
rect 579430 309922 579498 309978
rect 579554 309922 579622 309978
rect 579678 309922 579774 309978
rect 579154 292350 579774 309922
rect 579154 292294 579250 292350
rect 579306 292294 579374 292350
rect 579430 292294 579498 292350
rect 579554 292294 579622 292350
rect 579678 292294 579774 292350
rect 579154 292226 579774 292294
rect 579154 292170 579250 292226
rect 579306 292170 579374 292226
rect 579430 292170 579498 292226
rect 579554 292170 579622 292226
rect 579678 292170 579774 292226
rect 579154 292102 579774 292170
rect 579154 292046 579250 292102
rect 579306 292046 579374 292102
rect 579430 292046 579498 292102
rect 579554 292046 579622 292102
rect 579678 292046 579774 292102
rect 579154 291978 579774 292046
rect 579154 291922 579250 291978
rect 579306 291922 579374 291978
rect 579430 291922 579498 291978
rect 579554 291922 579622 291978
rect 579678 291922 579774 291978
rect 579154 274350 579774 291922
rect 579154 274294 579250 274350
rect 579306 274294 579374 274350
rect 579430 274294 579498 274350
rect 579554 274294 579622 274350
rect 579678 274294 579774 274350
rect 579154 274226 579774 274294
rect 579154 274170 579250 274226
rect 579306 274170 579374 274226
rect 579430 274170 579498 274226
rect 579554 274170 579622 274226
rect 579678 274170 579774 274226
rect 579154 274102 579774 274170
rect 579154 274046 579250 274102
rect 579306 274046 579374 274102
rect 579430 274046 579498 274102
rect 579554 274046 579622 274102
rect 579678 274046 579774 274102
rect 579154 273978 579774 274046
rect 579154 273922 579250 273978
rect 579306 273922 579374 273978
rect 579430 273922 579498 273978
rect 579554 273922 579622 273978
rect 579678 273922 579774 273978
rect 579154 256350 579774 273922
rect 579154 256294 579250 256350
rect 579306 256294 579374 256350
rect 579430 256294 579498 256350
rect 579554 256294 579622 256350
rect 579678 256294 579774 256350
rect 579154 256226 579774 256294
rect 579154 256170 579250 256226
rect 579306 256170 579374 256226
rect 579430 256170 579498 256226
rect 579554 256170 579622 256226
rect 579678 256170 579774 256226
rect 579154 256102 579774 256170
rect 579154 256046 579250 256102
rect 579306 256046 579374 256102
rect 579430 256046 579498 256102
rect 579554 256046 579622 256102
rect 579678 256046 579774 256102
rect 579154 255978 579774 256046
rect 579154 255922 579250 255978
rect 579306 255922 579374 255978
rect 579430 255922 579498 255978
rect 579554 255922 579622 255978
rect 579678 255922 579774 255978
rect 579154 238350 579774 255922
rect 579154 238294 579250 238350
rect 579306 238294 579374 238350
rect 579430 238294 579498 238350
rect 579554 238294 579622 238350
rect 579678 238294 579774 238350
rect 579154 238226 579774 238294
rect 579154 238170 579250 238226
rect 579306 238170 579374 238226
rect 579430 238170 579498 238226
rect 579554 238170 579622 238226
rect 579678 238170 579774 238226
rect 579154 238102 579774 238170
rect 579154 238046 579250 238102
rect 579306 238046 579374 238102
rect 579430 238046 579498 238102
rect 579554 238046 579622 238102
rect 579678 238046 579774 238102
rect 579154 237978 579774 238046
rect 579154 237922 579250 237978
rect 579306 237922 579374 237978
rect 579430 237922 579498 237978
rect 579554 237922 579622 237978
rect 579678 237922 579774 237978
rect 579154 220350 579774 237922
rect 579154 220294 579250 220350
rect 579306 220294 579374 220350
rect 579430 220294 579498 220350
rect 579554 220294 579622 220350
rect 579678 220294 579774 220350
rect 579154 220226 579774 220294
rect 579154 220170 579250 220226
rect 579306 220170 579374 220226
rect 579430 220170 579498 220226
rect 579554 220170 579622 220226
rect 579678 220170 579774 220226
rect 579154 220102 579774 220170
rect 579154 220046 579250 220102
rect 579306 220046 579374 220102
rect 579430 220046 579498 220102
rect 579554 220046 579622 220102
rect 579678 220046 579774 220102
rect 579154 219978 579774 220046
rect 579154 219922 579250 219978
rect 579306 219922 579374 219978
rect 579430 219922 579498 219978
rect 579554 219922 579622 219978
rect 579678 219922 579774 219978
rect 579154 202350 579774 219922
rect 579154 202294 579250 202350
rect 579306 202294 579374 202350
rect 579430 202294 579498 202350
rect 579554 202294 579622 202350
rect 579678 202294 579774 202350
rect 579154 202226 579774 202294
rect 579154 202170 579250 202226
rect 579306 202170 579374 202226
rect 579430 202170 579498 202226
rect 579554 202170 579622 202226
rect 579678 202170 579774 202226
rect 579154 202102 579774 202170
rect 579154 202046 579250 202102
rect 579306 202046 579374 202102
rect 579430 202046 579498 202102
rect 579554 202046 579622 202102
rect 579678 202046 579774 202102
rect 579154 201978 579774 202046
rect 579154 201922 579250 201978
rect 579306 201922 579374 201978
rect 579430 201922 579498 201978
rect 579554 201922 579622 201978
rect 579678 201922 579774 201978
rect 579154 184350 579774 201922
rect 579154 184294 579250 184350
rect 579306 184294 579374 184350
rect 579430 184294 579498 184350
rect 579554 184294 579622 184350
rect 579678 184294 579774 184350
rect 579154 184226 579774 184294
rect 579154 184170 579250 184226
rect 579306 184170 579374 184226
rect 579430 184170 579498 184226
rect 579554 184170 579622 184226
rect 579678 184170 579774 184226
rect 579154 184102 579774 184170
rect 579154 184046 579250 184102
rect 579306 184046 579374 184102
rect 579430 184046 579498 184102
rect 579554 184046 579622 184102
rect 579678 184046 579774 184102
rect 579154 183978 579774 184046
rect 579154 183922 579250 183978
rect 579306 183922 579374 183978
rect 579430 183922 579498 183978
rect 579554 183922 579622 183978
rect 579678 183922 579774 183978
rect 579154 166350 579774 183922
rect 579154 166294 579250 166350
rect 579306 166294 579374 166350
rect 579430 166294 579498 166350
rect 579554 166294 579622 166350
rect 579678 166294 579774 166350
rect 579154 166226 579774 166294
rect 579154 166170 579250 166226
rect 579306 166170 579374 166226
rect 579430 166170 579498 166226
rect 579554 166170 579622 166226
rect 579678 166170 579774 166226
rect 579154 166102 579774 166170
rect 579154 166046 579250 166102
rect 579306 166046 579374 166102
rect 579430 166046 579498 166102
rect 579554 166046 579622 166102
rect 579678 166046 579774 166102
rect 579154 165978 579774 166046
rect 579154 165922 579250 165978
rect 579306 165922 579374 165978
rect 579430 165922 579498 165978
rect 579554 165922 579622 165978
rect 579678 165922 579774 165978
rect 579154 148350 579774 165922
rect 579154 148294 579250 148350
rect 579306 148294 579374 148350
rect 579430 148294 579498 148350
rect 579554 148294 579622 148350
rect 579678 148294 579774 148350
rect 579154 148226 579774 148294
rect 579154 148170 579250 148226
rect 579306 148170 579374 148226
rect 579430 148170 579498 148226
rect 579554 148170 579622 148226
rect 579678 148170 579774 148226
rect 579154 148102 579774 148170
rect 579154 148046 579250 148102
rect 579306 148046 579374 148102
rect 579430 148046 579498 148102
rect 579554 148046 579622 148102
rect 579678 148046 579774 148102
rect 579154 147978 579774 148046
rect 579154 147922 579250 147978
rect 579306 147922 579374 147978
rect 579430 147922 579498 147978
rect 579554 147922 579622 147978
rect 579678 147922 579774 147978
rect 579154 130350 579774 147922
rect 579154 130294 579250 130350
rect 579306 130294 579374 130350
rect 579430 130294 579498 130350
rect 579554 130294 579622 130350
rect 579678 130294 579774 130350
rect 579154 130226 579774 130294
rect 579154 130170 579250 130226
rect 579306 130170 579374 130226
rect 579430 130170 579498 130226
rect 579554 130170 579622 130226
rect 579678 130170 579774 130226
rect 579154 130102 579774 130170
rect 579154 130046 579250 130102
rect 579306 130046 579374 130102
rect 579430 130046 579498 130102
rect 579554 130046 579622 130102
rect 579678 130046 579774 130102
rect 579154 129978 579774 130046
rect 579154 129922 579250 129978
rect 579306 129922 579374 129978
rect 579430 129922 579498 129978
rect 579554 129922 579622 129978
rect 579678 129922 579774 129978
rect 579154 112350 579774 129922
rect 579154 112294 579250 112350
rect 579306 112294 579374 112350
rect 579430 112294 579498 112350
rect 579554 112294 579622 112350
rect 579678 112294 579774 112350
rect 579154 112226 579774 112294
rect 579154 112170 579250 112226
rect 579306 112170 579374 112226
rect 579430 112170 579498 112226
rect 579554 112170 579622 112226
rect 579678 112170 579774 112226
rect 579154 112102 579774 112170
rect 579154 112046 579250 112102
rect 579306 112046 579374 112102
rect 579430 112046 579498 112102
rect 579554 112046 579622 112102
rect 579678 112046 579774 112102
rect 579154 111978 579774 112046
rect 579154 111922 579250 111978
rect 579306 111922 579374 111978
rect 579430 111922 579498 111978
rect 579554 111922 579622 111978
rect 579678 111922 579774 111978
rect 579154 94350 579774 111922
rect 579154 94294 579250 94350
rect 579306 94294 579374 94350
rect 579430 94294 579498 94350
rect 579554 94294 579622 94350
rect 579678 94294 579774 94350
rect 579154 94226 579774 94294
rect 579154 94170 579250 94226
rect 579306 94170 579374 94226
rect 579430 94170 579498 94226
rect 579554 94170 579622 94226
rect 579678 94170 579774 94226
rect 579154 94102 579774 94170
rect 579154 94046 579250 94102
rect 579306 94046 579374 94102
rect 579430 94046 579498 94102
rect 579554 94046 579622 94102
rect 579678 94046 579774 94102
rect 579154 93978 579774 94046
rect 579154 93922 579250 93978
rect 579306 93922 579374 93978
rect 579430 93922 579498 93978
rect 579554 93922 579622 93978
rect 579678 93922 579774 93978
rect 579154 76350 579774 93922
rect 579154 76294 579250 76350
rect 579306 76294 579374 76350
rect 579430 76294 579498 76350
rect 579554 76294 579622 76350
rect 579678 76294 579774 76350
rect 579154 76226 579774 76294
rect 579154 76170 579250 76226
rect 579306 76170 579374 76226
rect 579430 76170 579498 76226
rect 579554 76170 579622 76226
rect 579678 76170 579774 76226
rect 579154 76102 579774 76170
rect 579154 76046 579250 76102
rect 579306 76046 579374 76102
rect 579430 76046 579498 76102
rect 579554 76046 579622 76102
rect 579678 76046 579774 76102
rect 579154 75978 579774 76046
rect 579154 75922 579250 75978
rect 579306 75922 579374 75978
rect 579430 75922 579498 75978
rect 579554 75922 579622 75978
rect 579678 75922 579774 75978
rect 579154 58428 579774 75922
rect 579852 376628 579908 376638
rect 577052 42892 577108 42902
rect 577164 56942 578004 56998
rect 577164 37018 577220 56942
rect 577988 40412 579228 40446
rect 577988 40356 578022 40412
rect 578078 40356 578146 40412
rect 578202 40356 578270 40412
rect 578326 40356 578394 40412
rect 578450 40356 578518 40412
rect 578574 40356 578642 40412
rect 578698 40356 578766 40412
rect 578822 40356 578890 40412
rect 578946 40356 579014 40412
rect 579070 40356 579138 40412
rect 579194 40356 579228 40412
rect 577988 40288 579228 40356
rect 577988 40232 578022 40288
rect 578078 40232 578146 40288
rect 578202 40232 578270 40288
rect 578326 40232 578394 40288
rect 578450 40232 578518 40288
rect 578574 40232 578642 40288
rect 578698 40232 578766 40288
rect 578822 40232 578890 40288
rect 578946 40232 579014 40288
rect 579070 40232 579138 40288
rect 579194 40232 579228 40288
rect 577988 40164 579228 40232
rect 577988 40108 578022 40164
rect 578078 40108 578146 40164
rect 578202 40108 578270 40164
rect 578326 40108 578394 40164
rect 578450 40108 578518 40164
rect 578574 40108 578642 40164
rect 578698 40108 578766 40164
rect 578822 40108 578890 40164
rect 578946 40108 579014 40164
rect 579070 40108 579138 40164
rect 579194 40108 579228 40164
rect 577988 40040 579228 40108
rect 577988 39984 578022 40040
rect 578078 39984 578146 40040
rect 578202 39984 578270 40040
rect 578326 39984 578394 40040
rect 578450 39984 578518 40040
rect 578574 39984 578642 40040
rect 578698 39984 578766 40040
rect 578822 39984 578890 40040
rect 578946 39984 579014 40040
rect 579070 39984 579138 40040
rect 579194 39984 579228 40040
rect 577988 39916 579228 39984
rect 577988 39860 578022 39916
rect 578078 39860 578146 39916
rect 578202 39860 578270 39916
rect 578326 39860 578394 39916
rect 578450 39860 578518 39916
rect 578574 39860 578642 39916
rect 578698 39860 578766 39916
rect 578822 39860 578890 39916
rect 578946 39860 579014 39916
rect 579070 39860 579138 39916
rect 579194 39860 579228 39916
rect 577988 39826 579228 39860
rect 577164 36952 577220 36962
rect 577052 25318 577108 25328
rect 577052 20188 577108 25262
rect 577988 22412 579228 22446
rect 577988 22356 578022 22412
rect 578078 22356 578146 22412
rect 578202 22356 578270 22412
rect 578326 22356 578394 22412
rect 578450 22356 578518 22412
rect 578574 22356 578642 22412
rect 578698 22356 578766 22412
rect 578822 22356 578890 22412
rect 578946 22356 579014 22412
rect 579070 22356 579138 22412
rect 579194 22356 579228 22412
rect 577988 22288 579228 22356
rect 577988 22232 578022 22288
rect 578078 22232 578146 22288
rect 578202 22232 578270 22288
rect 578326 22232 578394 22288
rect 578450 22232 578518 22288
rect 578574 22232 578642 22288
rect 578698 22232 578766 22288
rect 578822 22232 578890 22288
rect 578946 22232 579014 22288
rect 579070 22232 579138 22288
rect 579194 22232 579228 22288
rect 577988 22164 579228 22232
rect 577988 22108 578022 22164
rect 578078 22108 578146 22164
rect 578202 22108 578270 22164
rect 578326 22108 578394 22164
rect 578450 22108 578518 22164
rect 578574 22108 578642 22164
rect 578698 22108 578766 22164
rect 578822 22108 578890 22164
rect 578946 22108 579014 22164
rect 579070 22108 579138 22164
rect 579194 22108 579228 22164
rect 577988 22040 579228 22108
rect 577988 21984 578022 22040
rect 578078 21984 578146 22040
rect 578202 21984 578270 22040
rect 578326 21984 578394 22040
rect 578450 21984 578518 22040
rect 578574 21984 578642 22040
rect 578698 21984 578766 22040
rect 578822 21984 578890 22040
rect 578946 21984 579014 22040
rect 579070 21984 579138 22040
rect 579194 21984 579228 22040
rect 577988 21916 579228 21984
rect 577988 21860 578022 21916
rect 578078 21860 578146 21916
rect 578202 21860 578270 21916
rect 578326 21860 578394 21916
rect 578450 21860 578518 21916
rect 578574 21860 578642 21916
rect 578698 21860 578766 21916
rect 578822 21860 578890 21916
rect 578946 21860 579014 21916
rect 579070 21860 579138 21916
rect 579194 21860 579228 21916
rect 577988 21826 579228 21860
rect 577052 20132 577220 20188
rect 576268 9314 576324 9324
rect 574812 8372 575092 8428
rect 575036 8306 575092 8316
rect 577052 8260 577108 8270
rect 577052 8038 577108 8204
rect 577052 7972 577108 7982
rect 574364 5954 574420 5964
rect 574476 6916 574532 6926
rect 574476 5908 574532 6860
rect 577164 6804 577220 20132
rect 577948 8148 578004 8158
rect 577948 7858 578004 8092
rect 577948 7792 578004 7802
rect 578844 8148 578900 8158
rect 578844 7678 578900 8092
rect 578844 7612 578900 7622
rect 577164 6738 577220 6748
rect 574476 5842 574532 5852
rect 572684 130 572740 140
rect 579154 4350 579774 10964
rect 579852 9268 579908 376572
rect 579964 10388 580020 376908
rect 579964 10322 580020 10332
rect 581308 376852 581364 376862
rect 581308 9604 581364 376796
rect 581532 376516 581588 376526
rect 581532 361228 581588 376460
rect 581420 361172 581588 361228
rect 582092 376516 582148 376526
rect 581420 37738 581476 361172
rect 582092 44578 582148 376460
rect 582092 44512 582148 44522
rect 582874 370350 583494 380034
rect 582874 370294 582970 370350
rect 583026 370294 583094 370350
rect 583150 370294 583218 370350
rect 583274 370294 583342 370350
rect 583398 370294 583494 370350
rect 582874 370226 583494 370294
rect 582874 370170 582970 370226
rect 583026 370170 583094 370226
rect 583150 370170 583218 370226
rect 583274 370170 583342 370226
rect 583398 370170 583494 370226
rect 582874 370102 583494 370170
rect 582874 370046 582970 370102
rect 583026 370046 583094 370102
rect 583150 370046 583218 370102
rect 583274 370046 583342 370102
rect 583398 370046 583494 370102
rect 582874 369978 583494 370046
rect 582874 369922 582970 369978
rect 583026 369922 583094 369978
rect 583150 369922 583218 369978
rect 583274 369922 583342 369978
rect 583398 369922 583494 369978
rect 582874 352350 583494 369922
rect 582874 352294 582970 352350
rect 583026 352294 583094 352350
rect 583150 352294 583218 352350
rect 583274 352294 583342 352350
rect 583398 352294 583494 352350
rect 582874 352226 583494 352294
rect 582874 352170 582970 352226
rect 583026 352170 583094 352226
rect 583150 352170 583218 352226
rect 583274 352170 583342 352226
rect 583398 352170 583494 352226
rect 582874 352102 583494 352170
rect 582874 352046 582970 352102
rect 583026 352046 583094 352102
rect 583150 352046 583218 352102
rect 583274 352046 583342 352102
rect 583398 352046 583494 352102
rect 582874 351978 583494 352046
rect 582874 351922 582970 351978
rect 583026 351922 583094 351978
rect 583150 351922 583218 351978
rect 583274 351922 583342 351978
rect 583398 351922 583494 351978
rect 582874 334350 583494 351922
rect 582874 334294 582970 334350
rect 583026 334294 583094 334350
rect 583150 334294 583218 334350
rect 583274 334294 583342 334350
rect 583398 334294 583494 334350
rect 582874 334226 583494 334294
rect 582874 334170 582970 334226
rect 583026 334170 583094 334226
rect 583150 334170 583218 334226
rect 583274 334170 583342 334226
rect 583398 334170 583494 334226
rect 582874 334102 583494 334170
rect 582874 334046 582970 334102
rect 583026 334046 583094 334102
rect 583150 334046 583218 334102
rect 583274 334046 583342 334102
rect 583398 334046 583494 334102
rect 582874 333978 583494 334046
rect 582874 333922 582970 333978
rect 583026 333922 583094 333978
rect 583150 333922 583218 333978
rect 583274 333922 583342 333978
rect 583398 333922 583494 333978
rect 582874 316350 583494 333922
rect 582874 316294 582970 316350
rect 583026 316294 583094 316350
rect 583150 316294 583218 316350
rect 583274 316294 583342 316350
rect 583398 316294 583494 316350
rect 582874 316226 583494 316294
rect 582874 316170 582970 316226
rect 583026 316170 583094 316226
rect 583150 316170 583218 316226
rect 583274 316170 583342 316226
rect 583398 316170 583494 316226
rect 582874 316102 583494 316170
rect 582874 316046 582970 316102
rect 583026 316046 583094 316102
rect 583150 316046 583218 316102
rect 583274 316046 583342 316102
rect 583398 316046 583494 316102
rect 582874 315978 583494 316046
rect 582874 315922 582970 315978
rect 583026 315922 583094 315978
rect 583150 315922 583218 315978
rect 583274 315922 583342 315978
rect 583398 315922 583494 315978
rect 582874 298350 583494 315922
rect 582874 298294 582970 298350
rect 583026 298294 583094 298350
rect 583150 298294 583218 298350
rect 583274 298294 583342 298350
rect 583398 298294 583494 298350
rect 582874 298226 583494 298294
rect 582874 298170 582970 298226
rect 583026 298170 583094 298226
rect 583150 298170 583218 298226
rect 583274 298170 583342 298226
rect 583398 298170 583494 298226
rect 582874 298102 583494 298170
rect 582874 298046 582970 298102
rect 583026 298046 583094 298102
rect 583150 298046 583218 298102
rect 583274 298046 583342 298102
rect 583398 298046 583494 298102
rect 582874 297978 583494 298046
rect 582874 297922 582970 297978
rect 583026 297922 583094 297978
rect 583150 297922 583218 297978
rect 583274 297922 583342 297978
rect 583398 297922 583494 297978
rect 582874 280350 583494 297922
rect 582874 280294 582970 280350
rect 583026 280294 583094 280350
rect 583150 280294 583218 280350
rect 583274 280294 583342 280350
rect 583398 280294 583494 280350
rect 582874 280226 583494 280294
rect 582874 280170 582970 280226
rect 583026 280170 583094 280226
rect 583150 280170 583218 280226
rect 583274 280170 583342 280226
rect 583398 280170 583494 280226
rect 582874 280102 583494 280170
rect 582874 280046 582970 280102
rect 583026 280046 583094 280102
rect 583150 280046 583218 280102
rect 583274 280046 583342 280102
rect 583398 280046 583494 280102
rect 582874 279978 583494 280046
rect 582874 279922 582970 279978
rect 583026 279922 583094 279978
rect 583150 279922 583218 279978
rect 583274 279922 583342 279978
rect 583398 279922 583494 279978
rect 582874 262350 583494 279922
rect 582874 262294 582970 262350
rect 583026 262294 583094 262350
rect 583150 262294 583218 262350
rect 583274 262294 583342 262350
rect 583398 262294 583494 262350
rect 582874 262226 583494 262294
rect 582874 262170 582970 262226
rect 583026 262170 583094 262226
rect 583150 262170 583218 262226
rect 583274 262170 583342 262226
rect 583398 262170 583494 262226
rect 582874 262102 583494 262170
rect 582874 262046 582970 262102
rect 583026 262046 583094 262102
rect 583150 262046 583218 262102
rect 583274 262046 583342 262102
rect 583398 262046 583494 262102
rect 582874 261978 583494 262046
rect 582874 261922 582970 261978
rect 583026 261922 583094 261978
rect 583150 261922 583218 261978
rect 583274 261922 583342 261978
rect 583398 261922 583494 261978
rect 582874 244350 583494 261922
rect 582874 244294 582970 244350
rect 583026 244294 583094 244350
rect 583150 244294 583218 244350
rect 583274 244294 583342 244350
rect 583398 244294 583494 244350
rect 582874 244226 583494 244294
rect 582874 244170 582970 244226
rect 583026 244170 583094 244226
rect 583150 244170 583218 244226
rect 583274 244170 583342 244226
rect 583398 244170 583494 244226
rect 582874 244102 583494 244170
rect 582874 244046 582970 244102
rect 583026 244046 583094 244102
rect 583150 244046 583218 244102
rect 583274 244046 583342 244102
rect 583398 244046 583494 244102
rect 582874 243978 583494 244046
rect 582874 243922 582970 243978
rect 583026 243922 583094 243978
rect 583150 243922 583218 243978
rect 583274 243922 583342 243978
rect 583398 243922 583494 243978
rect 582874 226350 583494 243922
rect 582874 226294 582970 226350
rect 583026 226294 583094 226350
rect 583150 226294 583218 226350
rect 583274 226294 583342 226350
rect 583398 226294 583494 226350
rect 582874 226226 583494 226294
rect 582874 226170 582970 226226
rect 583026 226170 583094 226226
rect 583150 226170 583218 226226
rect 583274 226170 583342 226226
rect 583398 226170 583494 226226
rect 582874 226102 583494 226170
rect 582874 226046 582970 226102
rect 583026 226046 583094 226102
rect 583150 226046 583218 226102
rect 583274 226046 583342 226102
rect 583398 226046 583494 226102
rect 582874 225978 583494 226046
rect 582874 225922 582970 225978
rect 583026 225922 583094 225978
rect 583150 225922 583218 225978
rect 583274 225922 583342 225978
rect 583398 225922 583494 225978
rect 582874 208350 583494 225922
rect 582874 208294 582970 208350
rect 583026 208294 583094 208350
rect 583150 208294 583218 208350
rect 583274 208294 583342 208350
rect 583398 208294 583494 208350
rect 582874 208226 583494 208294
rect 582874 208170 582970 208226
rect 583026 208170 583094 208226
rect 583150 208170 583218 208226
rect 583274 208170 583342 208226
rect 583398 208170 583494 208226
rect 582874 208102 583494 208170
rect 582874 208046 582970 208102
rect 583026 208046 583094 208102
rect 583150 208046 583218 208102
rect 583274 208046 583342 208102
rect 583398 208046 583494 208102
rect 582874 207978 583494 208046
rect 582874 207922 582970 207978
rect 583026 207922 583094 207978
rect 583150 207922 583218 207978
rect 583274 207922 583342 207978
rect 583398 207922 583494 207978
rect 582874 190350 583494 207922
rect 582874 190294 582970 190350
rect 583026 190294 583094 190350
rect 583150 190294 583218 190350
rect 583274 190294 583342 190350
rect 583398 190294 583494 190350
rect 582874 190226 583494 190294
rect 582874 190170 582970 190226
rect 583026 190170 583094 190226
rect 583150 190170 583218 190226
rect 583274 190170 583342 190226
rect 583398 190170 583494 190226
rect 582874 190102 583494 190170
rect 582874 190046 582970 190102
rect 583026 190046 583094 190102
rect 583150 190046 583218 190102
rect 583274 190046 583342 190102
rect 583398 190046 583494 190102
rect 582874 189978 583494 190046
rect 582874 189922 582970 189978
rect 583026 189922 583094 189978
rect 583150 189922 583218 189978
rect 583274 189922 583342 189978
rect 583398 189922 583494 189978
rect 582874 172350 583494 189922
rect 582874 172294 582970 172350
rect 583026 172294 583094 172350
rect 583150 172294 583218 172350
rect 583274 172294 583342 172350
rect 583398 172294 583494 172350
rect 582874 172226 583494 172294
rect 582874 172170 582970 172226
rect 583026 172170 583094 172226
rect 583150 172170 583218 172226
rect 583274 172170 583342 172226
rect 583398 172170 583494 172226
rect 582874 172102 583494 172170
rect 582874 172046 582970 172102
rect 583026 172046 583094 172102
rect 583150 172046 583218 172102
rect 583274 172046 583342 172102
rect 583398 172046 583494 172102
rect 582874 171978 583494 172046
rect 582874 171922 582970 171978
rect 583026 171922 583094 171978
rect 583150 171922 583218 171978
rect 583274 171922 583342 171978
rect 583398 171922 583494 171978
rect 582874 154350 583494 171922
rect 582874 154294 582970 154350
rect 583026 154294 583094 154350
rect 583150 154294 583218 154350
rect 583274 154294 583342 154350
rect 583398 154294 583494 154350
rect 582874 154226 583494 154294
rect 582874 154170 582970 154226
rect 583026 154170 583094 154226
rect 583150 154170 583218 154226
rect 583274 154170 583342 154226
rect 583398 154170 583494 154226
rect 582874 154102 583494 154170
rect 582874 154046 582970 154102
rect 583026 154046 583094 154102
rect 583150 154046 583218 154102
rect 583274 154046 583342 154102
rect 583398 154046 583494 154102
rect 582874 153978 583494 154046
rect 582874 153922 582970 153978
rect 583026 153922 583094 153978
rect 583150 153922 583218 153978
rect 583274 153922 583342 153978
rect 583398 153922 583494 153978
rect 582874 136350 583494 153922
rect 582874 136294 582970 136350
rect 583026 136294 583094 136350
rect 583150 136294 583218 136350
rect 583274 136294 583342 136350
rect 583398 136294 583494 136350
rect 582874 136226 583494 136294
rect 582874 136170 582970 136226
rect 583026 136170 583094 136226
rect 583150 136170 583218 136226
rect 583274 136170 583342 136226
rect 583398 136170 583494 136226
rect 582874 136102 583494 136170
rect 582874 136046 582970 136102
rect 583026 136046 583094 136102
rect 583150 136046 583218 136102
rect 583274 136046 583342 136102
rect 583398 136046 583494 136102
rect 582874 135978 583494 136046
rect 582874 135922 582970 135978
rect 583026 135922 583094 135978
rect 583150 135922 583218 135978
rect 583274 135922 583342 135978
rect 583398 135922 583494 135978
rect 582874 118350 583494 135922
rect 582874 118294 582970 118350
rect 583026 118294 583094 118350
rect 583150 118294 583218 118350
rect 583274 118294 583342 118350
rect 583398 118294 583494 118350
rect 582874 118226 583494 118294
rect 582874 118170 582970 118226
rect 583026 118170 583094 118226
rect 583150 118170 583218 118226
rect 583274 118170 583342 118226
rect 583398 118170 583494 118226
rect 582874 118102 583494 118170
rect 582874 118046 582970 118102
rect 583026 118046 583094 118102
rect 583150 118046 583218 118102
rect 583274 118046 583342 118102
rect 583398 118046 583494 118102
rect 582874 117978 583494 118046
rect 582874 117922 582970 117978
rect 583026 117922 583094 117978
rect 583150 117922 583218 117978
rect 583274 117922 583342 117978
rect 583398 117922 583494 117978
rect 582874 100350 583494 117922
rect 582874 100294 582970 100350
rect 583026 100294 583094 100350
rect 583150 100294 583218 100350
rect 583274 100294 583342 100350
rect 583398 100294 583494 100350
rect 582874 100226 583494 100294
rect 582874 100170 582970 100226
rect 583026 100170 583094 100226
rect 583150 100170 583218 100226
rect 583274 100170 583342 100226
rect 583398 100170 583494 100226
rect 582874 100102 583494 100170
rect 582874 100046 582970 100102
rect 583026 100046 583094 100102
rect 583150 100046 583218 100102
rect 583274 100046 583342 100102
rect 583398 100046 583494 100102
rect 582874 99978 583494 100046
rect 582874 99922 582970 99978
rect 583026 99922 583094 99978
rect 583150 99922 583218 99978
rect 583274 99922 583342 99978
rect 583398 99922 583494 99978
rect 582874 82350 583494 99922
rect 582874 82294 582970 82350
rect 583026 82294 583094 82350
rect 583150 82294 583218 82350
rect 583274 82294 583342 82350
rect 583398 82294 583494 82350
rect 582874 82226 583494 82294
rect 582874 82170 582970 82226
rect 583026 82170 583094 82226
rect 583150 82170 583218 82226
rect 583274 82170 583342 82226
rect 583398 82170 583494 82226
rect 582874 82102 583494 82170
rect 582874 82046 582970 82102
rect 583026 82046 583094 82102
rect 583150 82046 583218 82102
rect 583274 82046 583342 82102
rect 583398 82046 583494 82102
rect 582874 81978 583494 82046
rect 582874 81922 582970 81978
rect 583026 81922 583094 81978
rect 583150 81922 583218 81978
rect 583274 81922 583342 81978
rect 583398 81922 583494 81978
rect 582874 64350 583494 81922
rect 582874 64294 582970 64350
rect 583026 64294 583094 64350
rect 583150 64294 583218 64350
rect 583274 64294 583342 64350
rect 583398 64294 583494 64350
rect 582874 64226 583494 64294
rect 582874 64170 582970 64226
rect 583026 64170 583094 64226
rect 583150 64170 583218 64226
rect 583274 64170 583342 64226
rect 583398 64170 583494 64226
rect 582874 64102 583494 64170
rect 582874 64046 582970 64102
rect 583026 64046 583094 64102
rect 583150 64046 583218 64102
rect 583274 64046 583342 64102
rect 583398 64046 583494 64102
rect 582874 63978 583494 64046
rect 582874 63922 582970 63978
rect 583026 63922 583094 63978
rect 583150 63922 583218 63978
rect 583274 63922 583342 63978
rect 583398 63922 583494 63978
rect 582874 46350 583494 63922
rect 582874 46294 582970 46350
rect 583026 46294 583094 46350
rect 583150 46294 583218 46350
rect 583274 46294 583342 46350
rect 583398 46294 583494 46350
rect 582874 46226 583494 46294
rect 582874 46170 582970 46226
rect 583026 46170 583094 46226
rect 583150 46170 583218 46226
rect 583274 46170 583342 46226
rect 583398 46170 583494 46226
rect 582874 46102 583494 46170
rect 582874 46046 582970 46102
rect 583026 46046 583094 46102
rect 583150 46046 583218 46102
rect 583274 46046 583342 46102
rect 583398 46046 583494 46102
rect 582874 45978 583494 46046
rect 582874 45922 582970 45978
rect 583026 45922 583094 45978
rect 583150 45922 583218 45978
rect 583274 45922 583342 45978
rect 583398 45922 583494 45978
rect 581420 37672 581476 37682
rect 581308 9538 581364 9548
rect 582874 28350 583494 45922
rect 582874 28294 582970 28350
rect 583026 28294 583094 28350
rect 583150 28294 583218 28350
rect 583274 28294 583342 28350
rect 583398 28294 583494 28350
rect 582874 28226 583494 28294
rect 582874 28170 582970 28226
rect 583026 28170 583094 28226
rect 583150 28170 583218 28226
rect 583274 28170 583342 28226
rect 583398 28170 583494 28226
rect 582874 28102 583494 28170
rect 582874 28046 582970 28102
rect 583026 28046 583094 28102
rect 583150 28046 583218 28102
rect 583274 28046 583342 28102
rect 583398 28046 583494 28102
rect 582874 27978 583494 28046
rect 582874 27922 582970 27978
rect 583026 27922 583094 27978
rect 583150 27922 583218 27978
rect 583274 27922 583342 27978
rect 583398 27922 583494 27978
rect 582874 10350 583494 27922
rect 582874 10294 582970 10350
rect 583026 10294 583094 10350
rect 583150 10294 583218 10350
rect 583274 10294 583342 10350
rect 583398 10294 583494 10350
rect 582874 10226 583494 10294
rect 582874 10170 582970 10226
rect 583026 10170 583094 10226
rect 583150 10170 583218 10226
rect 583274 10170 583342 10226
rect 583398 10170 583494 10226
rect 582874 10102 583494 10170
rect 582874 10046 582970 10102
rect 583026 10046 583094 10102
rect 583150 10046 583218 10102
rect 583274 10046 583342 10102
rect 583398 10046 583494 10102
rect 582874 9978 583494 10046
rect 582874 9922 582970 9978
rect 583026 9922 583094 9978
rect 583150 9922 583218 9978
rect 583274 9922 583342 9978
rect 583398 9922 583494 9978
rect 579852 9202 579908 9212
rect 579852 8148 579908 8158
rect 579852 7498 579908 8092
rect 579852 7432 579908 7442
rect 579154 4294 579250 4350
rect 579306 4294 579374 4350
rect 579430 4294 579498 4350
rect 579554 4294 579622 4350
rect 579678 4294 579774 4350
rect 579154 4226 579774 4294
rect 579154 4170 579250 4226
rect 579306 4170 579374 4226
rect 579430 4170 579498 4226
rect 579554 4170 579622 4226
rect 579678 4170 579774 4226
rect 579154 4102 579774 4170
rect 579154 4046 579250 4102
rect 579306 4046 579374 4102
rect 579430 4046 579498 4102
rect 579554 4046 579622 4102
rect 579678 4046 579774 4102
rect 579154 3978 579774 4046
rect 579154 3922 579250 3978
rect 579306 3922 579374 3978
rect 579430 3922 579498 3978
rect 579554 3922 579622 3978
rect 579678 3922 579774 3978
rect 572572 18 572628 28
rect 564874 -1176 564970 -1120
rect 565026 -1176 565094 -1120
rect 565150 -1176 565218 -1120
rect 565274 -1176 565342 -1120
rect 565398 -1176 565494 -1120
rect 564874 -1244 565494 -1176
rect 564874 -1300 564970 -1244
rect 565026 -1300 565094 -1244
rect 565150 -1300 565218 -1244
rect 565274 -1300 565342 -1244
rect 565398 -1300 565494 -1244
rect 564874 -1368 565494 -1300
rect 564874 -1424 564970 -1368
rect 565026 -1424 565094 -1368
rect 565150 -1424 565218 -1368
rect 565274 -1424 565342 -1368
rect 565398 -1424 565494 -1368
rect 564874 -1492 565494 -1424
rect 564874 -1548 564970 -1492
rect 565026 -1548 565094 -1492
rect 565150 -1548 565218 -1492
rect 565274 -1548 565342 -1492
rect 565398 -1548 565494 -1492
rect 564874 -1644 565494 -1548
rect 579154 -160 579774 3922
rect 579154 -216 579250 -160
rect 579306 -216 579374 -160
rect 579430 -216 579498 -160
rect 579554 -216 579622 -160
rect 579678 -216 579774 -160
rect 579154 -284 579774 -216
rect 579154 -340 579250 -284
rect 579306 -340 579374 -284
rect 579430 -340 579498 -284
rect 579554 -340 579622 -284
rect 579678 -340 579774 -284
rect 579154 -408 579774 -340
rect 579154 -464 579250 -408
rect 579306 -464 579374 -408
rect 579430 -464 579498 -408
rect 579554 -464 579622 -408
rect 579678 -464 579774 -408
rect 579154 -532 579774 -464
rect 579154 -588 579250 -532
rect 579306 -588 579374 -532
rect 579430 -588 579498 -532
rect 579554 -588 579622 -532
rect 579678 -588 579774 -532
rect 579154 -1644 579774 -588
rect 582874 -1120 583494 9922
rect 584668 377860 584724 377870
rect 584668 9716 584724 377804
rect 586460 377636 586516 377646
rect 584892 376628 584948 376638
rect 584780 376516 584836 376526
rect 584780 41158 584836 376460
rect 584892 47818 584948 376572
rect 584892 47752 584948 47762
rect 586348 376516 586404 376526
rect 584780 41092 584836 41102
rect 586012 10738 586068 10748
rect 586012 10612 586068 10682
rect 586012 10546 586068 10556
rect 586348 9828 586404 376460
rect 586460 42778 586516 377580
rect 596400 364350 597020 381922
rect 596400 364294 596496 364350
rect 596552 364294 596620 364350
rect 596676 364294 596744 364350
rect 596800 364294 596868 364350
rect 596924 364294 597020 364350
rect 596400 364226 597020 364294
rect 596400 364170 596496 364226
rect 596552 364170 596620 364226
rect 596676 364170 596744 364226
rect 596800 364170 596868 364226
rect 596924 364170 597020 364226
rect 596400 364102 597020 364170
rect 596400 364046 596496 364102
rect 596552 364046 596620 364102
rect 596676 364046 596744 364102
rect 596800 364046 596868 364102
rect 596924 364046 597020 364102
rect 596400 363978 597020 364046
rect 596400 363922 596496 363978
rect 596552 363922 596620 363978
rect 596676 363922 596744 363978
rect 596800 363922 596868 363978
rect 596924 363922 597020 363978
rect 596400 346350 597020 363922
rect 596400 346294 596496 346350
rect 596552 346294 596620 346350
rect 596676 346294 596744 346350
rect 596800 346294 596868 346350
rect 596924 346294 597020 346350
rect 596400 346226 597020 346294
rect 596400 346170 596496 346226
rect 596552 346170 596620 346226
rect 596676 346170 596744 346226
rect 596800 346170 596868 346226
rect 596924 346170 597020 346226
rect 596400 346102 597020 346170
rect 596400 346046 596496 346102
rect 596552 346046 596620 346102
rect 596676 346046 596744 346102
rect 596800 346046 596868 346102
rect 596924 346046 597020 346102
rect 596400 345978 597020 346046
rect 596400 345922 596496 345978
rect 596552 345922 596620 345978
rect 596676 345922 596744 345978
rect 596800 345922 596868 345978
rect 596924 345922 597020 345978
rect 596400 328350 597020 345922
rect 596400 328294 596496 328350
rect 596552 328294 596620 328350
rect 596676 328294 596744 328350
rect 596800 328294 596868 328350
rect 596924 328294 597020 328350
rect 596400 328226 597020 328294
rect 596400 328170 596496 328226
rect 596552 328170 596620 328226
rect 596676 328170 596744 328226
rect 596800 328170 596868 328226
rect 596924 328170 597020 328226
rect 596400 328102 597020 328170
rect 596400 328046 596496 328102
rect 596552 328046 596620 328102
rect 596676 328046 596744 328102
rect 596800 328046 596868 328102
rect 596924 328046 597020 328102
rect 596400 327978 597020 328046
rect 596400 327922 596496 327978
rect 596552 327922 596620 327978
rect 596676 327922 596744 327978
rect 596800 327922 596868 327978
rect 596924 327922 597020 327978
rect 596400 310350 597020 327922
rect 596400 310294 596496 310350
rect 596552 310294 596620 310350
rect 596676 310294 596744 310350
rect 596800 310294 596868 310350
rect 596924 310294 597020 310350
rect 596400 310226 597020 310294
rect 596400 310170 596496 310226
rect 596552 310170 596620 310226
rect 596676 310170 596744 310226
rect 596800 310170 596868 310226
rect 596924 310170 597020 310226
rect 596400 310102 597020 310170
rect 596400 310046 596496 310102
rect 596552 310046 596620 310102
rect 596676 310046 596744 310102
rect 596800 310046 596868 310102
rect 596924 310046 597020 310102
rect 596400 309978 597020 310046
rect 596400 309922 596496 309978
rect 596552 309922 596620 309978
rect 596676 309922 596744 309978
rect 596800 309922 596868 309978
rect 596924 309922 597020 309978
rect 596400 292350 597020 309922
rect 596400 292294 596496 292350
rect 596552 292294 596620 292350
rect 596676 292294 596744 292350
rect 596800 292294 596868 292350
rect 596924 292294 597020 292350
rect 596400 292226 597020 292294
rect 596400 292170 596496 292226
rect 596552 292170 596620 292226
rect 596676 292170 596744 292226
rect 596800 292170 596868 292226
rect 596924 292170 597020 292226
rect 596400 292102 597020 292170
rect 596400 292046 596496 292102
rect 596552 292046 596620 292102
rect 596676 292046 596744 292102
rect 596800 292046 596868 292102
rect 596924 292046 597020 292102
rect 596400 291978 597020 292046
rect 596400 291922 596496 291978
rect 596552 291922 596620 291978
rect 596676 291922 596744 291978
rect 596800 291922 596868 291978
rect 596924 291922 597020 291978
rect 596400 274350 597020 291922
rect 596400 274294 596496 274350
rect 596552 274294 596620 274350
rect 596676 274294 596744 274350
rect 596800 274294 596868 274350
rect 596924 274294 597020 274350
rect 596400 274226 597020 274294
rect 596400 274170 596496 274226
rect 596552 274170 596620 274226
rect 596676 274170 596744 274226
rect 596800 274170 596868 274226
rect 596924 274170 597020 274226
rect 596400 274102 597020 274170
rect 596400 274046 596496 274102
rect 596552 274046 596620 274102
rect 596676 274046 596744 274102
rect 596800 274046 596868 274102
rect 596924 274046 597020 274102
rect 596400 273978 597020 274046
rect 596400 273922 596496 273978
rect 596552 273922 596620 273978
rect 596676 273922 596744 273978
rect 596800 273922 596868 273978
rect 596924 273922 597020 273978
rect 591276 271460 591332 271470
rect 591164 245028 591220 245038
rect 591052 205380 591108 205390
rect 591052 60452 591108 205324
rect 591052 60386 591108 60396
rect 591164 60340 591220 244972
rect 591164 60274 591220 60284
rect 587988 46412 589228 46446
rect 587988 46356 588022 46412
rect 588078 46356 588146 46412
rect 588202 46356 588270 46412
rect 588326 46356 588394 46412
rect 588450 46356 588518 46412
rect 588574 46356 588642 46412
rect 588698 46356 588766 46412
rect 588822 46356 588890 46412
rect 588946 46356 589014 46412
rect 589070 46356 589138 46412
rect 589194 46356 589228 46412
rect 587988 46288 589228 46356
rect 587988 46232 588022 46288
rect 588078 46232 588146 46288
rect 588202 46232 588270 46288
rect 588326 46232 588394 46288
rect 588450 46232 588518 46288
rect 588574 46232 588642 46288
rect 588698 46232 588766 46288
rect 588822 46232 588890 46288
rect 588946 46232 589014 46288
rect 589070 46232 589138 46288
rect 589194 46232 589228 46288
rect 587988 46164 589228 46232
rect 587988 46108 588022 46164
rect 588078 46108 588146 46164
rect 588202 46108 588270 46164
rect 588326 46108 588394 46164
rect 588450 46108 588518 46164
rect 588574 46108 588642 46164
rect 588698 46108 588766 46164
rect 588822 46108 588890 46164
rect 588946 46108 589014 46164
rect 589070 46108 589138 46164
rect 589194 46108 589228 46164
rect 587988 46040 589228 46108
rect 587988 45984 588022 46040
rect 588078 45984 588146 46040
rect 588202 45984 588270 46040
rect 588326 45984 588394 46040
rect 588450 45984 588518 46040
rect 588574 45984 588642 46040
rect 588698 45984 588766 46040
rect 588822 45984 588890 46040
rect 588946 45984 589014 46040
rect 589070 45984 589138 46040
rect 589194 45984 589228 46040
rect 587988 45916 589228 45984
rect 587988 45860 588022 45916
rect 588078 45860 588146 45916
rect 588202 45860 588270 45916
rect 588326 45860 588394 45916
rect 588450 45860 588518 45916
rect 588574 45860 588642 45916
rect 588698 45860 588766 45916
rect 588822 45860 588890 45916
rect 588946 45860 589014 45916
rect 589070 45860 589138 45916
rect 589194 45860 589228 45916
rect 587988 45826 589228 45860
rect 586460 42712 586516 42722
rect 591276 30178 591332 271404
rect 596400 256350 597020 273922
rect 596400 256294 596496 256350
rect 596552 256294 596620 256350
rect 596676 256294 596744 256350
rect 596800 256294 596868 256350
rect 596924 256294 597020 256350
rect 596400 256226 597020 256294
rect 596400 256170 596496 256226
rect 596552 256170 596620 256226
rect 596676 256170 596744 256226
rect 596800 256170 596868 256226
rect 596924 256170 597020 256226
rect 596400 256102 597020 256170
rect 596400 256046 596496 256102
rect 596552 256046 596620 256102
rect 596676 256046 596744 256102
rect 596800 256046 596868 256102
rect 596924 256046 597020 256102
rect 596400 255978 597020 256046
rect 596400 255922 596496 255978
rect 596552 255922 596620 255978
rect 596676 255922 596744 255978
rect 596800 255922 596868 255978
rect 596924 255922 597020 255978
rect 596400 238350 597020 255922
rect 596400 238294 596496 238350
rect 596552 238294 596620 238350
rect 596676 238294 596744 238350
rect 596800 238294 596868 238350
rect 596924 238294 597020 238350
rect 596400 238226 597020 238294
rect 596400 238170 596496 238226
rect 596552 238170 596620 238226
rect 596676 238170 596744 238226
rect 596800 238170 596868 238226
rect 596924 238170 597020 238226
rect 596400 238102 597020 238170
rect 596400 238046 596496 238102
rect 596552 238046 596620 238102
rect 596676 238046 596744 238102
rect 596800 238046 596868 238102
rect 596924 238046 597020 238102
rect 596400 237978 597020 238046
rect 596400 237922 596496 237978
rect 596552 237922 596620 237978
rect 596676 237922 596744 237978
rect 596800 237922 596868 237978
rect 596924 237922 597020 237978
rect 592956 231924 593012 231934
rect 592956 60418 593012 231868
rect 596400 220350 597020 237922
rect 596400 220294 596496 220350
rect 596552 220294 596620 220350
rect 596676 220294 596744 220350
rect 596800 220294 596868 220350
rect 596924 220294 597020 220350
rect 596400 220226 597020 220294
rect 596400 220170 596496 220226
rect 596552 220170 596620 220226
rect 596676 220170 596744 220226
rect 596800 220170 596868 220226
rect 596924 220170 597020 220226
rect 596400 220102 597020 220170
rect 596400 220046 596496 220102
rect 596552 220046 596620 220102
rect 596676 220046 596744 220102
rect 596800 220046 596868 220102
rect 596924 220046 597020 220102
rect 596400 219978 597020 220046
rect 596400 219922 596496 219978
rect 596552 219922 596620 219978
rect 596676 219922 596744 219978
rect 596800 219922 596868 219978
rect 596924 219922 597020 219978
rect 596400 202350 597020 219922
rect 596400 202294 596496 202350
rect 596552 202294 596620 202350
rect 596676 202294 596744 202350
rect 596800 202294 596868 202350
rect 596924 202294 597020 202350
rect 596400 202226 597020 202294
rect 596400 202170 596496 202226
rect 596552 202170 596620 202226
rect 596676 202170 596744 202226
rect 596800 202170 596868 202226
rect 596924 202170 597020 202226
rect 596400 202102 597020 202170
rect 596400 202046 596496 202102
rect 596552 202046 596620 202102
rect 596676 202046 596744 202102
rect 596800 202046 596868 202102
rect 596924 202046 597020 202102
rect 596400 201978 597020 202046
rect 596400 201922 596496 201978
rect 596552 201922 596620 201978
rect 596676 201922 596744 201978
rect 596800 201922 596868 201978
rect 596924 201922 597020 201978
rect 596400 184350 597020 201922
rect 596400 184294 596496 184350
rect 596552 184294 596620 184350
rect 596676 184294 596744 184350
rect 596800 184294 596868 184350
rect 596924 184294 597020 184350
rect 596400 184226 597020 184294
rect 596400 184170 596496 184226
rect 596552 184170 596620 184226
rect 596676 184170 596744 184226
rect 596800 184170 596868 184226
rect 596924 184170 597020 184226
rect 596400 184102 597020 184170
rect 596400 184046 596496 184102
rect 596552 184046 596620 184102
rect 596676 184046 596744 184102
rect 596800 184046 596868 184102
rect 596924 184046 597020 184102
rect 596400 183978 597020 184046
rect 596400 183922 596496 183978
rect 596552 183922 596620 183978
rect 596676 183922 596744 183978
rect 596800 183922 596868 183978
rect 596924 183922 597020 183978
rect 596400 166350 597020 183922
rect 596400 166294 596496 166350
rect 596552 166294 596620 166350
rect 596676 166294 596744 166350
rect 596800 166294 596868 166350
rect 596924 166294 597020 166350
rect 596400 166226 597020 166294
rect 596400 166170 596496 166226
rect 596552 166170 596620 166226
rect 596676 166170 596744 166226
rect 596800 166170 596868 166226
rect 596924 166170 597020 166226
rect 596400 166102 597020 166170
rect 596400 166046 596496 166102
rect 596552 166046 596620 166102
rect 596676 166046 596744 166102
rect 596800 166046 596868 166102
rect 596924 166046 597020 166102
rect 596400 165978 597020 166046
rect 596400 165922 596496 165978
rect 596552 165922 596620 165978
rect 596676 165922 596744 165978
rect 596800 165922 596868 165978
rect 596924 165922 597020 165978
rect 596400 148350 597020 165922
rect 596400 148294 596496 148350
rect 596552 148294 596620 148350
rect 596676 148294 596744 148350
rect 596800 148294 596868 148350
rect 596924 148294 597020 148350
rect 596400 148226 597020 148294
rect 596400 148170 596496 148226
rect 596552 148170 596620 148226
rect 596676 148170 596744 148226
rect 596800 148170 596868 148226
rect 596924 148170 597020 148226
rect 596400 148102 597020 148170
rect 596400 148046 596496 148102
rect 596552 148046 596620 148102
rect 596676 148046 596744 148102
rect 596800 148046 596868 148102
rect 596924 148046 597020 148102
rect 596400 147978 597020 148046
rect 596400 147922 596496 147978
rect 596552 147922 596620 147978
rect 596676 147922 596744 147978
rect 596800 147922 596868 147978
rect 596924 147922 597020 147978
rect 596400 130350 597020 147922
rect 596400 130294 596496 130350
rect 596552 130294 596620 130350
rect 596676 130294 596744 130350
rect 596800 130294 596868 130350
rect 596924 130294 597020 130350
rect 596400 130226 597020 130294
rect 596400 130170 596496 130226
rect 596552 130170 596620 130226
rect 596676 130170 596744 130226
rect 596800 130170 596868 130226
rect 596924 130170 597020 130226
rect 596400 130102 597020 130170
rect 596400 130046 596496 130102
rect 596552 130046 596620 130102
rect 596676 130046 596744 130102
rect 596800 130046 596868 130102
rect 596924 130046 597020 130102
rect 596400 129978 597020 130046
rect 596400 129922 596496 129978
rect 596552 129922 596620 129978
rect 596676 129922 596744 129978
rect 596800 129922 596868 129978
rect 596924 129922 597020 129978
rect 596400 112350 597020 129922
rect 596400 112294 596496 112350
rect 596552 112294 596620 112350
rect 596676 112294 596744 112350
rect 596800 112294 596868 112350
rect 596924 112294 597020 112350
rect 596400 112226 597020 112294
rect 596400 112170 596496 112226
rect 596552 112170 596620 112226
rect 596676 112170 596744 112226
rect 596800 112170 596868 112226
rect 596924 112170 597020 112226
rect 596400 112102 597020 112170
rect 596400 112046 596496 112102
rect 596552 112046 596620 112102
rect 596676 112046 596744 112102
rect 596800 112046 596868 112102
rect 596924 112046 597020 112102
rect 596400 111978 597020 112046
rect 596400 111922 596496 111978
rect 596552 111922 596620 111978
rect 596676 111922 596744 111978
rect 596800 111922 596868 111978
rect 596924 111922 597020 111978
rect 596400 94350 597020 111922
rect 596400 94294 596496 94350
rect 596552 94294 596620 94350
rect 596676 94294 596744 94350
rect 596800 94294 596868 94350
rect 596924 94294 597020 94350
rect 596400 94226 597020 94294
rect 596400 94170 596496 94226
rect 596552 94170 596620 94226
rect 596676 94170 596744 94226
rect 596800 94170 596868 94226
rect 596924 94170 597020 94226
rect 596400 94102 597020 94170
rect 596400 94046 596496 94102
rect 596552 94046 596620 94102
rect 596676 94046 596744 94102
rect 596800 94046 596868 94102
rect 596924 94046 597020 94102
rect 596400 93978 597020 94046
rect 596400 93922 596496 93978
rect 596552 93922 596620 93978
rect 596676 93922 596744 93978
rect 596800 93922 596868 93978
rect 596924 93922 597020 93978
rect 596400 76350 597020 93922
rect 596400 76294 596496 76350
rect 596552 76294 596620 76350
rect 596676 76294 596744 76350
rect 596800 76294 596868 76350
rect 596924 76294 597020 76350
rect 596400 76226 597020 76294
rect 596400 76170 596496 76226
rect 596552 76170 596620 76226
rect 596676 76170 596744 76226
rect 596800 76170 596868 76226
rect 596924 76170 597020 76226
rect 596400 76102 597020 76170
rect 596400 76046 596496 76102
rect 596552 76046 596620 76102
rect 596676 76046 596744 76102
rect 596800 76046 596868 76102
rect 596924 76046 597020 76102
rect 596400 75978 597020 76046
rect 596400 75922 596496 75978
rect 596552 75922 596620 75978
rect 596676 75922 596744 75978
rect 596800 75922 596868 75978
rect 596924 75922 597020 75978
rect 593404 60452 593460 60462
rect 592956 60362 593124 60418
rect 591276 30112 591332 30122
rect 591388 60228 591444 60238
rect 587988 28412 589228 28446
rect 587988 28356 588022 28412
rect 588078 28356 588146 28412
rect 588202 28356 588270 28412
rect 588326 28356 588394 28412
rect 588450 28356 588518 28412
rect 588574 28356 588642 28412
rect 588698 28356 588766 28412
rect 588822 28356 588890 28412
rect 588946 28356 589014 28412
rect 589070 28356 589138 28412
rect 589194 28356 589228 28412
rect 587988 28288 589228 28356
rect 587988 28232 588022 28288
rect 588078 28232 588146 28288
rect 588202 28232 588270 28288
rect 588326 28232 588394 28288
rect 588450 28232 588518 28288
rect 588574 28232 588642 28288
rect 588698 28232 588766 28288
rect 588822 28232 588890 28288
rect 588946 28232 589014 28288
rect 589070 28232 589138 28288
rect 589194 28232 589228 28288
rect 587988 28164 589228 28232
rect 587988 28108 588022 28164
rect 588078 28108 588146 28164
rect 588202 28108 588270 28164
rect 588326 28108 588394 28164
rect 588450 28108 588518 28164
rect 588574 28108 588642 28164
rect 588698 28108 588766 28164
rect 588822 28108 588890 28164
rect 588946 28108 589014 28164
rect 589070 28108 589138 28164
rect 589194 28108 589228 28164
rect 587988 28040 589228 28108
rect 587988 27984 588022 28040
rect 588078 27984 588146 28040
rect 588202 27984 588270 28040
rect 588326 27984 588394 28040
rect 588450 27984 588518 28040
rect 588574 27984 588642 28040
rect 588698 27984 588766 28040
rect 588822 27984 588890 28040
rect 588946 27984 589014 28040
rect 589070 27984 589138 28040
rect 589194 27984 589228 28040
rect 587988 27916 589228 27984
rect 587988 27860 588022 27916
rect 588078 27860 588146 27916
rect 588202 27860 588270 27916
rect 588326 27860 588394 27916
rect 588450 27860 588518 27916
rect 588574 27860 588642 27916
rect 588698 27860 588766 27916
rect 588822 27860 588890 27916
rect 588946 27860 589014 27916
rect 589070 27860 589138 27916
rect 589194 27860 589228 27916
rect 587988 27826 589228 27860
rect 591388 25138 591444 60172
rect 593068 55468 593124 60362
rect 593068 55412 593348 55468
rect 593292 53284 593348 55412
rect 593292 53218 593348 53228
rect 593292 30178 593348 30188
rect 593292 28644 593348 30122
rect 593292 28578 593348 28588
rect 591388 10612 591444 25082
rect 593404 16324 593460 60396
rect 593516 60340 593572 60350
rect 593516 40964 593572 60284
rect 593516 40898 593572 40908
rect 596400 58350 597020 75922
rect 596400 58294 596496 58350
rect 596552 58294 596620 58350
rect 596676 58294 596744 58350
rect 596800 58294 596868 58350
rect 596924 58294 597020 58350
rect 596400 58226 597020 58294
rect 596400 58170 596496 58226
rect 596552 58170 596620 58226
rect 596676 58170 596744 58226
rect 596800 58170 596868 58226
rect 596924 58170 597020 58226
rect 596400 58102 597020 58170
rect 596400 58046 596496 58102
rect 596552 58046 596620 58102
rect 596676 58046 596744 58102
rect 596800 58046 596868 58102
rect 596924 58046 597020 58102
rect 596400 57978 597020 58046
rect 596400 57922 596496 57978
rect 596552 57922 596620 57978
rect 596676 57922 596744 57978
rect 596800 57922 596868 57978
rect 596924 57922 597020 57978
rect 593404 16258 593460 16268
rect 596400 40350 597020 57922
rect 596400 40294 596496 40350
rect 596552 40294 596620 40350
rect 596676 40294 596744 40350
rect 596800 40294 596868 40350
rect 596924 40294 597020 40350
rect 596400 40226 597020 40294
rect 596400 40170 596496 40226
rect 596552 40170 596620 40226
rect 596676 40170 596744 40226
rect 596800 40170 596868 40226
rect 596924 40170 597020 40226
rect 596400 40102 597020 40170
rect 596400 40046 596496 40102
rect 596552 40046 596620 40102
rect 596676 40046 596744 40102
rect 596800 40046 596868 40102
rect 596924 40046 597020 40102
rect 596400 39978 597020 40046
rect 596400 39922 596496 39978
rect 596552 39922 596620 39978
rect 596676 39922 596744 39978
rect 596800 39922 596868 39978
rect 596924 39922 597020 39978
rect 596400 22350 597020 39922
rect 596400 22294 596496 22350
rect 596552 22294 596620 22350
rect 596676 22294 596744 22350
rect 596800 22294 596868 22350
rect 596924 22294 597020 22350
rect 596400 22226 597020 22294
rect 596400 22170 596496 22226
rect 596552 22170 596620 22226
rect 596676 22170 596744 22226
rect 596800 22170 596868 22226
rect 596924 22170 597020 22226
rect 596400 22102 597020 22170
rect 596400 22046 596496 22102
rect 596552 22046 596620 22102
rect 596676 22046 596744 22102
rect 596800 22046 596868 22102
rect 596924 22046 597020 22102
rect 596400 21978 597020 22046
rect 596400 21922 596496 21978
rect 596552 21922 596620 21978
rect 596676 21922 596744 21978
rect 596800 21922 596868 21978
rect 596924 21922 597020 21978
rect 591388 10546 591444 10556
rect 586348 9762 586404 9772
rect 584668 9650 584724 9660
rect 596400 4350 597020 21922
rect 596400 4294 596496 4350
rect 596552 4294 596620 4350
rect 596676 4294 596744 4350
rect 596800 4294 596868 4350
rect 596924 4294 597020 4350
rect 596400 4226 597020 4294
rect 596400 4170 596496 4226
rect 596552 4170 596620 4226
rect 596676 4170 596744 4226
rect 596800 4170 596868 4226
rect 596924 4170 597020 4226
rect 596400 4102 597020 4170
rect 596400 4046 596496 4102
rect 596552 4046 596620 4102
rect 596676 4046 596744 4102
rect 596800 4046 596868 4102
rect 596924 4046 597020 4102
rect 596400 3978 597020 4046
rect 596400 3922 596496 3978
rect 596552 3922 596620 3978
rect 596676 3922 596744 3978
rect 596800 3922 596868 3978
rect 596924 3922 597020 3978
rect 596400 -160 597020 3922
rect 596400 -216 596496 -160
rect 596552 -216 596620 -160
rect 596676 -216 596744 -160
rect 596800 -216 596868 -160
rect 596924 -216 597020 -160
rect 596400 -284 597020 -216
rect 596400 -340 596496 -284
rect 596552 -340 596620 -284
rect 596676 -340 596744 -284
rect 596800 -340 596868 -284
rect 596924 -340 597020 -284
rect 596400 -408 597020 -340
rect 596400 -464 596496 -408
rect 596552 -464 596620 -408
rect 596676 -464 596744 -408
rect 596800 -464 596868 -408
rect 596924 -464 597020 -408
rect 596400 -532 597020 -464
rect 596400 -588 596496 -532
rect 596552 -588 596620 -532
rect 596676 -588 596744 -532
rect 596800 -588 596868 -532
rect 596924 -588 597020 -532
rect 596400 -684 597020 -588
rect 597360 586350 597980 597744
rect 597360 586294 597456 586350
rect 597512 586294 597580 586350
rect 597636 586294 597704 586350
rect 597760 586294 597828 586350
rect 597884 586294 597980 586350
rect 597360 586226 597980 586294
rect 597360 586170 597456 586226
rect 597512 586170 597580 586226
rect 597636 586170 597704 586226
rect 597760 586170 597828 586226
rect 597884 586170 597980 586226
rect 597360 586102 597980 586170
rect 597360 586046 597456 586102
rect 597512 586046 597580 586102
rect 597636 586046 597704 586102
rect 597760 586046 597828 586102
rect 597884 586046 597980 586102
rect 597360 585978 597980 586046
rect 597360 585922 597456 585978
rect 597512 585922 597580 585978
rect 597636 585922 597704 585978
rect 597760 585922 597828 585978
rect 597884 585922 597980 585978
rect 597360 568350 597980 585922
rect 597360 568294 597456 568350
rect 597512 568294 597580 568350
rect 597636 568294 597704 568350
rect 597760 568294 597828 568350
rect 597884 568294 597980 568350
rect 597360 568226 597980 568294
rect 597360 568170 597456 568226
rect 597512 568170 597580 568226
rect 597636 568170 597704 568226
rect 597760 568170 597828 568226
rect 597884 568170 597980 568226
rect 597360 568102 597980 568170
rect 597360 568046 597456 568102
rect 597512 568046 597580 568102
rect 597636 568046 597704 568102
rect 597760 568046 597828 568102
rect 597884 568046 597980 568102
rect 597360 567978 597980 568046
rect 597360 567922 597456 567978
rect 597512 567922 597580 567978
rect 597636 567922 597704 567978
rect 597760 567922 597828 567978
rect 597884 567922 597980 567978
rect 597360 550350 597980 567922
rect 597360 550294 597456 550350
rect 597512 550294 597580 550350
rect 597636 550294 597704 550350
rect 597760 550294 597828 550350
rect 597884 550294 597980 550350
rect 597360 550226 597980 550294
rect 597360 550170 597456 550226
rect 597512 550170 597580 550226
rect 597636 550170 597704 550226
rect 597760 550170 597828 550226
rect 597884 550170 597980 550226
rect 597360 550102 597980 550170
rect 597360 550046 597456 550102
rect 597512 550046 597580 550102
rect 597636 550046 597704 550102
rect 597760 550046 597828 550102
rect 597884 550046 597980 550102
rect 597360 549978 597980 550046
rect 597360 549922 597456 549978
rect 597512 549922 597580 549978
rect 597636 549922 597704 549978
rect 597760 549922 597828 549978
rect 597884 549922 597980 549978
rect 597360 532350 597980 549922
rect 597360 532294 597456 532350
rect 597512 532294 597580 532350
rect 597636 532294 597704 532350
rect 597760 532294 597828 532350
rect 597884 532294 597980 532350
rect 597360 532226 597980 532294
rect 597360 532170 597456 532226
rect 597512 532170 597580 532226
rect 597636 532170 597704 532226
rect 597760 532170 597828 532226
rect 597884 532170 597980 532226
rect 597360 532102 597980 532170
rect 597360 532046 597456 532102
rect 597512 532046 597580 532102
rect 597636 532046 597704 532102
rect 597760 532046 597828 532102
rect 597884 532046 597980 532102
rect 597360 531978 597980 532046
rect 597360 531922 597456 531978
rect 597512 531922 597580 531978
rect 597636 531922 597704 531978
rect 597760 531922 597828 531978
rect 597884 531922 597980 531978
rect 597360 514350 597980 531922
rect 597360 514294 597456 514350
rect 597512 514294 597580 514350
rect 597636 514294 597704 514350
rect 597760 514294 597828 514350
rect 597884 514294 597980 514350
rect 597360 514226 597980 514294
rect 597360 514170 597456 514226
rect 597512 514170 597580 514226
rect 597636 514170 597704 514226
rect 597760 514170 597828 514226
rect 597884 514170 597980 514226
rect 597360 514102 597980 514170
rect 597360 514046 597456 514102
rect 597512 514046 597580 514102
rect 597636 514046 597704 514102
rect 597760 514046 597828 514102
rect 597884 514046 597980 514102
rect 597360 513978 597980 514046
rect 597360 513922 597456 513978
rect 597512 513922 597580 513978
rect 597636 513922 597704 513978
rect 597760 513922 597828 513978
rect 597884 513922 597980 513978
rect 597360 496350 597980 513922
rect 597360 496294 597456 496350
rect 597512 496294 597580 496350
rect 597636 496294 597704 496350
rect 597760 496294 597828 496350
rect 597884 496294 597980 496350
rect 597360 496226 597980 496294
rect 597360 496170 597456 496226
rect 597512 496170 597580 496226
rect 597636 496170 597704 496226
rect 597760 496170 597828 496226
rect 597884 496170 597980 496226
rect 597360 496102 597980 496170
rect 597360 496046 597456 496102
rect 597512 496046 597580 496102
rect 597636 496046 597704 496102
rect 597760 496046 597828 496102
rect 597884 496046 597980 496102
rect 597360 495978 597980 496046
rect 597360 495922 597456 495978
rect 597512 495922 597580 495978
rect 597636 495922 597704 495978
rect 597760 495922 597828 495978
rect 597884 495922 597980 495978
rect 597360 478350 597980 495922
rect 597360 478294 597456 478350
rect 597512 478294 597580 478350
rect 597636 478294 597704 478350
rect 597760 478294 597828 478350
rect 597884 478294 597980 478350
rect 597360 478226 597980 478294
rect 597360 478170 597456 478226
rect 597512 478170 597580 478226
rect 597636 478170 597704 478226
rect 597760 478170 597828 478226
rect 597884 478170 597980 478226
rect 597360 478102 597980 478170
rect 597360 478046 597456 478102
rect 597512 478046 597580 478102
rect 597636 478046 597704 478102
rect 597760 478046 597828 478102
rect 597884 478046 597980 478102
rect 597360 477978 597980 478046
rect 597360 477922 597456 477978
rect 597512 477922 597580 477978
rect 597636 477922 597704 477978
rect 597760 477922 597828 477978
rect 597884 477922 597980 477978
rect 597360 460350 597980 477922
rect 597360 460294 597456 460350
rect 597512 460294 597580 460350
rect 597636 460294 597704 460350
rect 597760 460294 597828 460350
rect 597884 460294 597980 460350
rect 597360 460226 597980 460294
rect 597360 460170 597456 460226
rect 597512 460170 597580 460226
rect 597636 460170 597704 460226
rect 597760 460170 597828 460226
rect 597884 460170 597980 460226
rect 597360 460102 597980 460170
rect 597360 460046 597456 460102
rect 597512 460046 597580 460102
rect 597636 460046 597704 460102
rect 597760 460046 597828 460102
rect 597884 460046 597980 460102
rect 597360 459978 597980 460046
rect 597360 459922 597456 459978
rect 597512 459922 597580 459978
rect 597636 459922 597704 459978
rect 597760 459922 597828 459978
rect 597884 459922 597980 459978
rect 597360 442350 597980 459922
rect 597360 442294 597456 442350
rect 597512 442294 597580 442350
rect 597636 442294 597704 442350
rect 597760 442294 597828 442350
rect 597884 442294 597980 442350
rect 597360 442226 597980 442294
rect 597360 442170 597456 442226
rect 597512 442170 597580 442226
rect 597636 442170 597704 442226
rect 597760 442170 597828 442226
rect 597884 442170 597980 442226
rect 597360 442102 597980 442170
rect 597360 442046 597456 442102
rect 597512 442046 597580 442102
rect 597636 442046 597704 442102
rect 597760 442046 597828 442102
rect 597884 442046 597980 442102
rect 597360 441978 597980 442046
rect 597360 441922 597456 441978
rect 597512 441922 597580 441978
rect 597636 441922 597704 441978
rect 597760 441922 597828 441978
rect 597884 441922 597980 441978
rect 597360 424350 597980 441922
rect 597360 424294 597456 424350
rect 597512 424294 597580 424350
rect 597636 424294 597704 424350
rect 597760 424294 597828 424350
rect 597884 424294 597980 424350
rect 597360 424226 597980 424294
rect 597360 424170 597456 424226
rect 597512 424170 597580 424226
rect 597636 424170 597704 424226
rect 597760 424170 597828 424226
rect 597884 424170 597980 424226
rect 597360 424102 597980 424170
rect 597360 424046 597456 424102
rect 597512 424046 597580 424102
rect 597636 424046 597704 424102
rect 597760 424046 597828 424102
rect 597884 424046 597980 424102
rect 597360 423978 597980 424046
rect 597360 423922 597456 423978
rect 597512 423922 597580 423978
rect 597636 423922 597704 423978
rect 597760 423922 597828 423978
rect 597884 423922 597980 423978
rect 597360 406350 597980 423922
rect 597360 406294 597456 406350
rect 597512 406294 597580 406350
rect 597636 406294 597704 406350
rect 597760 406294 597828 406350
rect 597884 406294 597980 406350
rect 597360 406226 597980 406294
rect 597360 406170 597456 406226
rect 597512 406170 597580 406226
rect 597636 406170 597704 406226
rect 597760 406170 597828 406226
rect 597884 406170 597980 406226
rect 597360 406102 597980 406170
rect 597360 406046 597456 406102
rect 597512 406046 597580 406102
rect 597636 406046 597704 406102
rect 597760 406046 597828 406102
rect 597884 406046 597980 406102
rect 597360 405978 597980 406046
rect 597360 405922 597456 405978
rect 597512 405922 597580 405978
rect 597636 405922 597704 405978
rect 597760 405922 597828 405978
rect 597884 405922 597980 405978
rect 597360 388350 597980 405922
rect 597360 388294 597456 388350
rect 597512 388294 597580 388350
rect 597636 388294 597704 388350
rect 597760 388294 597828 388350
rect 597884 388294 597980 388350
rect 597360 388226 597980 388294
rect 597360 388170 597456 388226
rect 597512 388170 597580 388226
rect 597636 388170 597704 388226
rect 597760 388170 597828 388226
rect 597884 388170 597980 388226
rect 597360 388102 597980 388170
rect 597360 388046 597456 388102
rect 597512 388046 597580 388102
rect 597636 388046 597704 388102
rect 597760 388046 597828 388102
rect 597884 388046 597980 388102
rect 597360 387978 597980 388046
rect 597360 387922 597456 387978
rect 597512 387922 597580 387978
rect 597636 387922 597704 387978
rect 597760 387922 597828 387978
rect 597884 387922 597980 387978
rect 597360 370350 597980 387922
rect 597360 370294 597456 370350
rect 597512 370294 597580 370350
rect 597636 370294 597704 370350
rect 597760 370294 597828 370350
rect 597884 370294 597980 370350
rect 597360 370226 597980 370294
rect 597360 370170 597456 370226
rect 597512 370170 597580 370226
rect 597636 370170 597704 370226
rect 597760 370170 597828 370226
rect 597884 370170 597980 370226
rect 597360 370102 597980 370170
rect 597360 370046 597456 370102
rect 597512 370046 597580 370102
rect 597636 370046 597704 370102
rect 597760 370046 597828 370102
rect 597884 370046 597980 370102
rect 597360 369978 597980 370046
rect 597360 369922 597456 369978
rect 597512 369922 597580 369978
rect 597636 369922 597704 369978
rect 597760 369922 597828 369978
rect 597884 369922 597980 369978
rect 597360 352350 597980 369922
rect 597360 352294 597456 352350
rect 597512 352294 597580 352350
rect 597636 352294 597704 352350
rect 597760 352294 597828 352350
rect 597884 352294 597980 352350
rect 597360 352226 597980 352294
rect 597360 352170 597456 352226
rect 597512 352170 597580 352226
rect 597636 352170 597704 352226
rect 597760 352170 597828 352226
rect 597884 352170 597980 352226
rect 597360 352102 597980 352170
rect 597360 352046 597456 352102
rect 597512 352046 597580 352102
rect 597636 352046 597704 352102
rect 597760 352046 597828 352102
rect 597884 352046 597980 352102
rect 597360 351978 597980 352046
rect 597360 351922 597456 351978
rect 597512 351922 597580 351978
rect 597636 351922 597704 351978
rect 597760 351922 597828 351978
rect 597884 351922 597980 351978
rect 597360 334350 597980 351922
rect 597360 334294 597456 334350
rect 597512 334294 597580 334350
rect 597636 334294 597704 334350
rect 597760 334294 597828 334350
rect 597884 334294 597980 334350
rect 597360 334226 597980 334294
rect 597360 334170 597456 334226
rect 597512 334170 597580 334226
rect 597636 334170 597704 334226
rect 597760 334170 597828 334226
rect 597884 334170 597980 334226
rect 597360 334102 597980 334170
rect 597360 334046 597456 334102
rect 597512 334046 597580 334102
rect 597636 334046 597704 334102
rect 597760 334046 597828 334102
rect 597884 334046 597980 334102
rect 597360 333978 597980 334046
rect 597360 333922 597456 333978
rect 597512 333922 597580 333978
rect 597636 333922 597704 333978
rect 597760 333922 597828 333978
rect 597884 333922 597980 333978
rect 597360 316350 597980 333922
rect 597360 316294 597456 316350
rect 597512 316294 597580 316350
rect 597636 316294 597704 316350
rect 597760 316294 597828 316350
rect 597884 316294 597980 316350
rect 597360 316226 597980 316294
rect 597360 316170 597456 316226
rect 597512 316170 597580 316226
rect 597636 316170 597704 316226
rect 597760 316170 597828 316226
rect 597884 316170 597980 316226
rect 597360 316102 597980 316170
rect 597360 316046 597456 316102
rect 597512 316046 597580 316102
rect 597636 316046 597704 316102
rect 597760 316046 597828 316102
rect 597884 316046 597980 316102
rect 597360 315978 597980 316046
rect 597360 315922 597456 315978
rect 597512 315922 597580 315978
rect 597636 315922 597704 315978
rect 597760 315922 597828 315978
rect 597884 315922 597980 315978
rect 597360 298350 597980 315922
rect 597360 298294 597456 298350
rect 597512 298294 597580 298350
rect 597636 298294 597704 298350
rect 597760 298294 597828 298350
rect 597884 298294 597980 298350
rect 597360 298226 597980 298294
rect 597360 298170 597456 298226
rect 597512 298170 597580 298226
rect 597636 298170 597704 298226
rect 597760 298170 597828 298226
rect 597884 298170 597980 298226
rect 597360 298102 597980 298170
rect 597360 298046 597456 298102
rect 597512 298046 597580 298102
rect 597636 298046 597704 298102
rect 597760 298046 597828 298102
rect 597884 298046 597980 298102
rect 597360 297978 597980 298046
rect 597360 297922 597456 297978
rect 597512 297922 597580 297978
rect 597636 297922 597704 297978
rect 597760 297922 597828 297978
rect 597884 297922 597980 297978
rect 597360 280350 597980 297922
rect 597360 280294 597456 280350
rect 597512 280294 597580 280350
rect 597636 280294 597704 280350
rect 597760 280294 597828 280350
rect 597884 280294 597980 280350
rect 597360 280226 597980 280294
rect 597360 280170 597456 280226
rect 597512 280170 597580 280226
rect 597636 280170 597704 280226
rect 597760 280170 597828 280226
rect 597884 280170 597980 280226
rect 597360 280102 597980 280170
rect 597360 280046 597456 280102
rect 597512 280046 597580 280102
rect 597636 280046 597704 280102
rect 597760 280046 597828 280102
rect 597884 280046 597980 280102
rect 597360 279978 597980 280046
rect 597360 279922 597456 279978
rect 597512 279922 597580 279978
rect 597636 279922 597704 279978
rect 597760 279922 597828 279978
rect 597884 279922 597980 279978
rect 597360 262350 597980 279922
rect 597360 262294 597456 262350
rect 597512 262294 597580 262350
rect 597636 262294 597704 262350
rect 597760 262294 597828 262350
rect 597884 262294 597980 262350
rect 597360 262226 597980 262294
rect 597360 262170 597456 262226
rect 597512 262170 597580 262226
rect 597636 262170 597704 262226
rect 597760 262170 597828 262226
rect 597884 262170 597980 262226
rect 597360 262102 597980 262170
rect 597360 262046 597456 262102
rect 597512 262046 597580 262102
rect 597636 262046 597704 262102
rect 597760 262046 597828 262102
rect 597884 262046 597980 262102
rect 597360 261978 597980 262046
rect 597360 261922 597456 261978
rect 597512 261922 597580 261978
rect 597636 261922 597704 261978
rect 597760 261922 597828 261978
rect 597884 261922 597980 261978
rect 597360 244350 597980 261922
rect 597360 244294 597456 244350
rect 597512 244294 597580 244350
rect 597636 244294 597704 244350
rect 597760 244294 597828 244350
rect 597884 244294 597980 244350
rect 597360 244226 597980 244294
rect 597360 244170 597456 244226
rect 597512 244170 597580 244226
rect 597636 244170 597704 244226
rect 597760 244170 597828 244226
rect 597884 244170 597980 244226
rect 597360 244102 597980 244170
rect 597360 244046 597456 244102
rect 597512 244046 597580 244102
rect 597636 244046 597704 244102
rect 597760 244046 597828 244102
rect 597884 244046 597980 244102
rect 597360 243978 597980 244046
rect 597360 243922 597456 243978
rect 597512 243922 597580 243978
rect 597636 243922 597704 243978
rect 597760 243922 597828 243978
rect 597884 243922 597980 243978
rect 597360 226350 597980 243922
rect 597360 226294 597456 226350
rect 597512 226294 597580 226350
rect 597636 226294 597704 226350
rect 597760 226294 597828 226350
rect 597884 226294 597980 226350
rect 597360 226226 597980 226294
rect 597360 226170 597456 226226
rect 597512 226170 597580 226226
rect 597636 226170 597704 226226
rect 597760 226170 597828 226226
rect 597884 226170 597980 226226
rect 597360 226102 597980 226170
rect 597360 226046 597456 226102
rect 597512 226046 597580 226102
rect 597636 226046 597704 226102
rect 597760 226046 597828 226102
rect 597884 226046 597980 226102
rect 597360 225978 597980 226046
rect 597360 225922 597456 225978
rect 597512 225922 597580 225978
rect 597636 225922 597704 225978
rect 597760 225922 597828 225978
rect 597884 225922 597980 225978
rect 597360 208350 597980 225922
rect 597360 208294 597456 208350
rect 597512 208294 597580 208350
rect 597636 208294 597704 208350
rect 597760 208294 597828 208350
rect 597884 208294 597980 208350
rect 597360 208226 597980 208294
rect 597360 208170 597456 208226
rect 597512 208170 597580 208226
rect 597636 208170 597704 208226
rect 597760 208170 597828 208226
rect 597884 208170 597980 208226
rect 597360 208102 597980 208170
rect 597360 208046 597456 208102
rect 597512 208046 597580 208102
rect 597636 208046 597704 208102
rect 597760 208046 597828 208102
rect 597884 208046 597980 208102
rect 597360 207978 597980 208046
rect 597360 207922 597456 207978
rect 597512 207922 597580 207978
rect 597636 207922 597704 207978
rect 597760 207922 597828 207978
rect 597884 207922 597980 207978
rect 597360 190350 597980 207922
rect 597360 190294 597456 190350
rect 597512 190294 597580 190350
rect 597636 190294 597704 190350
rect 597760 190294 597828 190350
rect 597884 190294 597980 190350
rect 597360 190226 597980 190294
rect 597360 190170 597456 190226
rect 597512 190170 597580 190226
rect 597636 190170 597704 190226
rect 597760 190170 597828 190226
rect 597884 190170 597980 190226
rect 597360 190102 597980 190170
rect 597360 190046 597456 190102
rect 597512 190046 597580 190102
rect 597636 190046 597704 190102
rect 597760 190046 597828 190102
rect 597884 190046 597980 190102
rect 597360 189978 597980 190046
rect 597360 189922 597456 189978
rect 597512 189922 597580 189978
rect 597636 189922 597704 189978
rect 597760 189922 597828 189978
rect 597884 189922 597980 189978
rect 597360 172350 597980 189922
rect 597360 172294 597456 172350
rect 597512 172294 597580 172350
rect 597636 172294 597704 172350
rect 597760 172294 597828 172350
rect 597884 172294 597980 172350
rect 597360 172226 597980 172294
rect 597360 172170 597456 172226
rect 597512 172170 597580 172226
rect 597636 172170 597704 172226
rect 597760 172170 597828 172226
rect 597884 172170 597980 172226
rect 597360 172102 597980 172170
rect 597360 172046 597456 172102
rect 597512 172046 597580 172102
rect 597636 172046 597704 172102
rect 597760 172046 597828 172102
rect 597884 172046 597980 172102
rect 597360 171978 597980 172046
rect 597360 171922 597456 171978
rect 597512 171922 597580 171978
rect 597636 171922 597704 171978
rect 597760 171922 597828 171978
rect 597884 171922 597980 171978
rect 597360 154350 597980 171922
rect 597360 154294 597456 154350
rect 597512 154294 597580 154350
rect 597636 154294 597704 154350
rect 597760 154294 597828 154350
rect 597884 154294 597980 154350
rect 597360 154226 597980 154294
rect 597360 154170 597456 154226
rect 597512 154170 597580 154226
rect 597636 154170 597704 154226
rect 597760 154170 597828 154226
rect 597884 154170 597980 154226
rect 597360 154102 597980 154170
rect 597360 154046 597456 154102
rect 597512 154046 597580 154102
rect 597636 154046 597704 154102
rect 597760 154046 597828 154102
rect 597884 154046 597980 154102
rect 597360 153978 597980 154046
rect 597360 153922 597456 153978
rect 597512 153922 597580 153978
rect 597636 153922 597704 153978
rect 597760 153922 597828 153978
rect 597884 153922 597980 153978
rect 597360 136350 597980 153922
rect 597360 136294 597456 136350
rect 597512 136294 597580 136350
rect 597636 136294 597704 136350
rect 597760 136294 597828 136350
rect 597884 136294 597980 136350
rect 597360 136226 597980 136294
rect 597360 136170 597456 136226
rect 597512 136170 597580 136226
rect 597636 136170 597704 136226
rect 597760 136170 597828 136226
rect 597884 136170 597980 136226
rect 597360 136102 597980 136170
rect 597360 136046 597456 136102
rect 597512 136046 597580 136102
rect 597636 136046 597704 136102
rect 597760 136046 597828 136102
rect 597884 136046 597980 136102
rect 597360 135978 597980 136046
rect 597360 135922 597456 135978
rect 597512 135922 597580 135978
rect 597636 135922 597704 135978
rect 597760 135922 597828 135978
rect 597884 135922 597980 135978
rect 597360 118350 597980 135922
rect 597360 118294 597456 118350
rect 597512 118294 597580 118350
rect 597636 118294 597704 118350
rect 597760 118294 597828 118350
rect 597884 118294 597980 118350
rect 597360 118226 597980 118294
rect 597360 118170 597456 118226
rect 597512 118170 597580 118226
rect 597636 118170 597704 118226
rect 597760 118170 597828 118226
rect 597884 118170 597980 118226
rect 597360 118102 597980 118170
rect 597360 118046 597456 118102
rect 597512 118046 597580 118102
rect 597636 118046 597704 118102
rect 597760 118046 597828 118102
rect 597884 118046 597980 118102
rect 597360 117978 597980 118046
rect 597360 117922 597456 117978
rect 597512 117922 597580 117978
rect 597636 117922 597704 117978
rect 597760 117922 597828 117978
rect 597884 117922 597980 117978
rect 597360 100350 597980 117922
rect 597360 100294 597456 100350
rect 597512 100294 597580 100350
rect 597636 100294 597704 100350
rect 597760 100294 597828 100350
rect 597884 100294 597980 100350
rect 597360 100226 597980 100294
rect 597360 100170 597456 100226
rect 597512 100170 597580 100226
rect 597636 100170 597704 100226
rect 597760 100170 597828 100226
rect 597884 100170 597980 100226
rect 597360 100102 597980 100170
rect 597360 100046 597456 100102
rect 597512 100046 597580 100102
rect 597636 100046 597704 100102
rect 597760 100046 597828 100102
rect 597884 100046 597980 100102
rect 597360 99978 597980 100046
rect 597360 99922 597456 99978
rect 597512 99922 597580 99978
rect 597636 99922 597704 99978
rect 597760 99922 597828 99978
rect 597884 99922 597980 99978
rect 597360 82350 597980 99922
rect 597360 82294 597456 82350
rect 597512 82294 597580 82350
rect 597636 82294 597704 82350
rect 597760 82294 597828 82350
rect 597884 82294 597980 82350
rect 597360 82226 597980 82294
rect 597360 82170 597456 82226
rect 597512 82170 597580 82226
rect 597636 82170 597704 82226
rect 597760 82170 597828 82226
rect 597884 82170 597980 82226
rect 597360 82102 597980 82170
rect 597360 82046 597456 82102
rect 597512 82046 597580 82102
rect 597636 82046 597704 82102
rect 597760 82046 597828 82102
rect 597884 82046 597980 82102
rect 597360 81978 597980 82046
rect 597360 81922 597456 81978
rect 597512 81922 597580 81978
rect 597636 81922 597704 81978
rect 597760 81922 597828 81978
rect 597884 81922 597980 81978
rect 597360 64350 597980 81922
rect 597360 64294 597456 64350
rect 597512 64294 597580 64350
rect 597636 64294 597704 64350
rect 597760 64294 597828 64350
rect 597884 64294 597980 64350
rect 597360 64226 597980 64294
rect 597360 64170 597456 64226
rect 597512 64170 597580 64226
rect 597636 64170 597704 64226
rect 597760 64170 597828 64226
rect 597884 64170 597980 64226
rect 597360 64102 597980 64170
rect 597360 64046 597456 64102
rect 597512 64046 597580 64102
rect 597636 64046 597704 64102
rect 597760 64046 597828 64102
rect 597884 64046 597980 64102
rect 597360 63978 597980 64046
rect 597360 63922 597456 63978
rect 597512 63922 597580 63978
rect 597636 63922 597704 63978
rect 597760 63922 597828 63978
rect 597884 63922 597980 63978
rect 597360 46350 597980 63922
rect 597360 46294 597456 46350
rect 597512 46294 597580 46350
rect 597636 46294 597704 46350
rect 597760 46294 597828 46350
rect 597884 46294 597980 46350
rect 597360 46226 597980 46294
rect 597360 46170 597456 46226
rect 597512 46170 597580 46226
rect 597636 46170 597704 46226
rect 597760 46170 597828 46226
rect 597884 46170 597980 46226
rect 597360 46102 597980 46170
rect 597360 46046 597456 46102
rect 597512 46046 597580 46102
rect 597636 46046 597704 46102
rect 597760 46046 597828 46102
rect 597884 46046 597980 46102
rect 597360 45978 597980 46046
rect 597360 45922 597456 45978
rect 597512 45922 597580 45978
rect 597636 45922 597704 45978
rect 597760 45922 597828 45978
rect 597884 45922 597980 45978
rect 597360 28350 597980 45922
rect 597360 28294 597456 28350
rect 597512 28294 597580 28350
rect 597636 28294 597704 28350
rect 597760 28294 597828 28350
rect 597884 28294 597980 28350
rect 597360 28226 597980 28294
rect 597360 28170 597456 28226
rect 597512 28170 597580 28226
rect 597636 28170 597704 28226
rect 597760 28170 597828 28226
rect 597884 28170 597980 28226
rect 597360 28102 597980 28170
rect 597360 28046 597456 28102
rect 597512 28046 597580 28102
rect 597636 28046 597704 28102
rect 597760 28046 597828 28102
rect 597884 28046 597980 28102
rect 597360 27978 597980 28046
rect 597360 27922 597456 27978
rect 597512 27922 597580 27978
rect 597636 27922 597704 27978
rect 597760 27922 597828 27978
rect 597884 27922 597980 27978
rect 597360 10350 597980 27922
rect 597360 10294 597456 10350
rect 597512 10294 597580 10350
rect 597636 10294 597704 10350
rect 597760 10294 597828 10350
rect 597884 10294 597980 10350
rect 597360 10226 597980 10294
rect 597360 10170 597456 10226
rect 597512 10170 597580 10226
rect 597636 10170 597704 10226
rect 597760 10170 597828 10226
rect 597884 10170 597980 10226
rect 597360 10102 597980 10170
rect 597360 10046 597456 10102
rect 597512 10046 597580 10102
rect 597636 10046 597704 10102
rect 597760 10046 597828 10102
rect 597884 10046 597980 10102
rect 597360 9978 597980 10046
rect 597360 9922 597456 9978
rect 597512 9922 597580 9978
rect 597636 9922 597704 9978
rect 597760 9922 597828 9978
rect 597884 9922 597980 9978
rect 582874 -1176 582970 -1120
rect 583026 -1176 583094 -1120
rect 583150 -1176 583218 -1120
rect 583274 -1176 583342 -1120
rect 583398 -1176 583494 -1120
rect 582874 -1244 583494 -1176
rect 582874 -1300 582970 -1244
rect 583026 -1300 583094 -1244
rect 583150 -1300 583218 -1244
rect 583274 -1300 583342 -1244
rect 583398 -1300 583494 -1244
rect 582874 -1368 583494 -1300
rect 582874 -1424 582970 -1368
rect 583026 -1424 583094 -1368
rect 583150 -1424 583218 -1368
rect 583274 -1424 583342 -1368
rect 583398 -1424 583494 -1368
rect 582874 -1492 583494 -1424
rect 582874 -1548 582970 -1492
rect 583026 -1548 583094 -1492
rect 583150 -1548 583218 -1492
rect 583274 -1548 583342 -1492
rect 583398 -1548 583494 -1492
rect 582874 -1644 583494 -1548
rect 597360 -1120 597980 9922
rect 597360 -1176 597456 -1120
rect 597512 -1176 597580 -1120
rect 597636 -1176 597704 -1120
rect 597760 -1176 597828 -1120
rect 597884 -1176 597980 -1120
rect 597360 -1244 597980 -1176
rect 597360 -1300 597456 -1244
rect 597512 -1300 597580 -1244
rect 597636 -1300 597704 -1244
rect 597760 -1300 597828 -1244
rect 597884 -1300 597980 -1244
rect 597360 -1368 597980 -1300
rect 597360 -1424 597456 -1368
rect 597512 -1424 597580 -1368
rect 597636 -1424 597704 -1368
rect 597760 -1424 597828 -1368
rect 597884 -1424 597980 -1368
rect 597360 -1492 597980 -1424
rect 597360 -1548 597456 -1492
rect 597512 -1548 597580 -1492
rect 597636 -1548 597704 -1492
rect 597760 -1548 597828 -1492
rect 597884 -1548 597980 -1492
rect 597360 -1644 597980 -1548
<< via4 >>
rect -1820 598116 -1764 598172
rect -1696 598116 -1640 598172
rect -1572 598116 -1516 598172
rect -1448 598116 -1392 598172
rect -1820 597992 -1764 598048
rect -1696 597992 -1640 598048
rect -1572 597992 -1516 598048
rect -1448 597992 -1392 598048
rect -1820 597868 -1764 597924
rect -1696 597868 -1640 597924
rect -1572 597868 -1516 597924
rect -1448 597868 -1392 597924
rect -1820 597744 -1764 597800
rect -1696 597744 -1640 597800
rect -1572 597744 -1516 597800
rect -1448 597744 -1392 597800
rect -1820 586294 -1764 586350
rect -1696 586294 -1640 586350
rect -1572 586294 -1516 586350
rect -1448 586294 -1392 586350
rect -1820 586170 -1764 586226
rect -1696 586170 -1640 586226
rect -1572 586170 -1516 586226
rect -1448 586170 -1392 586226
rect -1820 586046 -1764 586102
rect -1696 586046 -1640 586102
rect -1572 586046 -1516 586102
rect -1448 586046 -1392 586102
rect -1820 585922 -1764 585978
rect -1696 585922 -1640 585978
rect -1572 585922 -1516 585978
rect -1448 585922 -1392 585978
rect -1820 568294 -1764 568350
rect -1696 568294 -1640 568350
rect -1572 568294 -1516 568350
rect -1448 568294 -1392 568350
rect -1820 568170 -1764 568226
rect -1696 568170 -1640 568226
rect -1572 568170 -1516 568226
rect -1448 568170 -1392 568226
rect -1820 568046 -1764 568102
rect -1696 568046 -1640 568102
rect -1572 568046 -1516 568102
rect -1448 568046 -1392 568102
rect -1820 567922 -1764 567978
rect -1696 567922 -1640 567978
rect -1572 567922 -1516 567978
rect -1448 567922 -1392 567978
rect -1820 550294 -1764 550350
rect -1696 550294 -1640 550350
rect -1572 550294 -1516 550350
rect -1448 550294 -1392 550350
rect -1820 550170 -1764 550226
rect -1696 550170 -1640 550226
rect -1572 550170 -1516 550226
rect -1448 550170 -1392 550226
rect -1820 550046 -1764 550102
rect -1696 550046 -1640 550102
rect -1572 550046 -1516 550102
rect -1448 550046 -1392 550102
rect -1820 549922 -1764 549978
rect -1696 549922 -1640 549978
rect -1572 549922 -1516 549978
rect -1448 549922 -1392 549978
rect -1820 532294 -1764 532350
rect -1696 532294 -1640 532350
rect -1572 532294 -1516 532350
rect -1448 532294 -1392 532350
rect -1820 532170 -1764 532226
rect -1696 532170 -1640 532226
rect -1572 532170 -1516 532226
rect -1448 532170 -1392 532226
rect -1820 532046 -1764 532102
rect -1696 532046 -1640 532102
rect -1572 532046 -1516 532102
rect -1448 532046 -1392 532102
rect -1820 531922 -1764 531978
rect -1696 531922 -1640 531978
rect -1572 531922 -1516 531978
rect -1448 531922 -1392 531978
rect -1820 514294 -1764 514350
rect -1696 514294 -1640 514350
rect -1572 514294 -1516 514350
rect -1448 514294 -1392 514350
rect -1820 514170 -1764 514226
rect -1696 514170 -1640 514226
rect -1572 514170 -1516 514226
rect -1448 514170 -1392 514226
rect -1820 514046 -1764 514102
rect -1696 514046 -1640 514102
rect -1572 514046 -1516 514102
rect -1448 514046 -1392 514102
rect -1820 513922 -1764 513978
rect -1696 513922 -1640 513978
rect -1572 513922 -1516 513978
rect -1448 513922 -1392 513978
rect -1820 496294 -1764 496350
rect -1696 496294 -1640 496350
rect -1572 496294 -1516 496350
rect -1448 496294 -1392 496350
rect -1820 496170 -1764 496226
rect -1696 496170 -1640 496226
rect -1572 496170 -1516 496226
rect -1448 496170 -1392 496226
rect -1820 496046 -1764 496102
rect -1696 496046 -1640 496102
rect -1572 496046 -1516 496102
rect -1448 496046 -1392 496102
rect -1820 495922 -1764 495978
rect -1696 495922 -1640 495978
rect -1572 495922 -1516 495978
rect -1448 495922 -1392 495978
rect -1820 478294 -1764 478350
rect -1696 478294 -1640 478350
rect -1572 478294 -1516 478350
rect -1448 478294 -1392 478350
rect -1820 478170 -1764 478226
rect -1696 478170 -1640 478226
rect -1572 478170 -1516 478226
rect -1448 478170 -1392 478226
rect -1820 478046 -1764 478102
rect -1696 478046 -1640 478102
rect -1572 478046 -1516 478102
rect -1448 478046 -1392 478102
rect -1820 477922 -1764 477978
rect -1696 477922 -1640 477978
rect -1572 477922 -1516 477978
rect -1448 477922 -1392 477978
rect -1820 460294 -1764 460350
rect -1696 460294 -1640 460350
rect -1572 460294 -1516 460350
rect -1448 460294 -1392 460350
rect -1820 460170 -1764 460226
rect -1696 460170 -1640 460226
rect -1572 460170 -1516 460226
rect -1448 460170 -1392 460226
rect -1820 460046 -1764 460102
rect -1696 460046 -1640 460102
rect -1572 460046 -1516 460102
rect -1448 460046 -1392 460102
rect -1820 459922 -1764 459978
rect -1696 459922 -1640 459978
rect -1572 459922 -1516 459978
rect -1448 459922 -1392 459978
rect -1820 442294 -1764 442350
rect -1696 442294 -1640 442350
rect -1572 442294 -1516 442350
rect -1448 442294 -1392 442350
rect -1820 442170 -1764 442226
rect -1696 442170 -1640 442226
rect -1572 442170 -1516 442226
rect -1448 442170 -1392 442226
rect -1820 442046 -1764 442102
rect -1696 442046 -1640 442102
rect -1572 442046 -1516 442102
rect -1448 442046 -1392 442102
rect -1820 441922 -1764 441978
rect -1696 441922 -1640 441978
rect -1572 441922 -1516 441978
rect -1448 441922 -1392 441978
rect -1820 424294 -1764 424350
rect -1696 424294 -1640 424350
rect -1572 424294 -1516 424350
rect -1448 424294 -1392 424350
rect -1820 424170 -1764 424226
rect -1696 424170 -1640 424226
rect -1572 424170 -1516 424226
rect -1448 424170 -1392 424226
rect -1820 424046 -1764 424102
rect -1696 424046 -1640 424102
rect -1572 424046 -1516 424102
rect -1448 424046 -1392 424102
rect -1820 423922 -1764 423978
rect -1696 423922 -1640 423978
rect -1572 423922 -1516 423978
rect -1448 423922 -1392 423978
rect -1820 406294 -1764 406350
rect -1696 406294 -1640 406350
rect -1572 406294 -1516 406350
rect -1448 406294 -1392 406350
rect -1820 406170 -1764 406226
rect -1696 406170 -1640 406226
rect -1572 406170 -1516 406226
rect -1448 406170 -1392 406226
rect -1820 406046 -1764 406102
rect -1696 406046 -1640 406102
rect -1572 406046 -1516 406102
rect -1448 406046 -1392 406102
rect -1820 405922 -1764 405978
rect -1696 405922 -1640 405978
rect -1572 405922 -1516 405978
rect -1448 405922 -1392 405978
rect -1820 388294 -1764 388350
rect -1696 388294 -1640 388350
rect -1572 388294 -1516 388350
rect -1448 388294 -1392 388350
rect -1820 388170 -1764 388226
rect -1696 388170 -1640 388226
rect -1572 388170 -1516 388226
rect -1448 388170 -1392 388226
rect -1820 388046 -1764 388102
rect -1696 388046 -1640 388102
rect -1572 388046 -1516 388102
rect -1448 388046 -1392 388102
rect -1820 387922 -1764 387978
rect -1696 387922 -1640 387978
rect -1572 387922 -1516 387978
rect -1448 387922 -1392 387978
rect -1820 370294 -1764 370350
rect -1696 370294 -1640 370350
rect -1572 370294 -1516 370350
rect -1448 370294 -1392 370350
rect -1820 370170 -1764 370226
rect -1696 370170 -1640 370226
rect -1572 370170 -1516 370226
rect -1448 370170 -1392 370226
rect -1820 370046 -1764 370102
rect -1696 370046 -1640 370102
rect -1572 370046 -1516 370102
rect -1448 370046 -1392 370102
rect -1820 369922 -1764 369978
rect -1696 369922 -1640 369978
rect -1572 369922 -1516 369978
rect -1448 369922 -1392 369978
rect -1820 352294 -1764 352350
rect -1696 352294 -1640 352350
rect -1572 352294 -1516 352350
rect -1448 352294 -1392 352350
rect -1820 352170 -1764 352226
rect -1696 352170 -1640 352226
rect -1572 352170 -1516 352226
rect -1448 352170 -1392 352226
rect -1820 352046 -1764 352102
rect -1696 352046 -1640 352102
rect -1572 352046 -1516 352102
rect -1448 352046 -1392 352102
rect -1820 351922 -1764 351978
rect -1696 351922 -1640 351978
rect -1572 351922 -1516 351978
rect -1448 351922 -1392 351978
rect -1820 334294 -1764 334350
rect -1696 334294 -1640 334350
rect -1572 334294 -1516 334350
rect -1448 334294 -1392 334350
rect -1820 334170 -1764 334226
rect -1696 334170 -1640 334226
rect -1572 334170 -1516 334226
rect -1448 334170 -1392 334226
rect -1820 334046 -1764 334102
rect -1696 334046 -1640 334102
rect -1572 334046 -1516 334102
rect -1448 334046 -1392 334102
rect -1820 333922 -1764 333978
rect -1696 333922 -1640 333978
rect -1572 333922 -1516 333978
rect -1448 333922 -1392 333978
rect -1820 316294 -1764 316350
rect -1696 316294 -1640 316350
rect -1572 316294 -1516 316350
rect -1448 316294 -1392 316350
rect -1820 316170 -1764 316226
rect -1696 316170 -1640 316226
rect -1572 316170 -1516 316226
rect -1448 316170 -1392 316226
rect -1820 316046 -1764 316102
rect -1696 316046 -1640 316102
rect -1572 316046 -1516 316102
rect -1448 316046 -1392 316102
rect -1820 315922 -1764 315978
rect -1696 315922 -1640 315978
rect -1572 315922 -1516 315978
rect -1448 315922 -1392 315978
rect -1820 298294 -1764 298350
rect -1696 298294 -1640 298350
rect -1572 298294 -1516 298350
rect -1448 298294 -1392 298350
rect -1820 298170 -1764 298226
rect -1696 298170 -1640 298226
rect -1572 298170 -1516 298226
rect -1448 298170 -1392 298226
rect -1820 298046 -1764 298102
rect -1696 298046 -1640 298102
rect -1572 298046 -1516 298102
rect -1448 298046 -1392 298102
rect -1820 297922 -1764 297978
rect -1696 297922 -1640 297978
rect -1572 297922 -1516 297978
rect -1448 297922 -1392 297978
rect -1820 280294 -1764 280350
rect -1696 280294 -1640 280350
rect -1572 280294 -1516 280350
rect -1448 280294 -1392 280350
rect -1820 280170 -1764 280226
rect -1696 280170 -1640 280226
rect -1572 280170 -1516 280226
rect -1448 280170 -1392 280226
rect -1820 280046 -1764 280102
rect -1696 280046 -1640 280102
rect -1572 280046 -1516 280102
rect -1448 280046 -1392 280102
rect -1820 279922 -1764 279978
rect -1696 279922 -1640 279978
rect -1572 279922 -1516 279978
rect -1448 279922 -1392 279978
rect -1820 262294 -1764 262350
rect -1696 262294 -1640 262350
rect -1572 262294 -1516 262350
rect -1448 262294 -1392 262350
rect -1820 262170 -1764 262226
rect -1696 262170 -1640 262226
rect -1572 262170 -1516 262226
rect -1448 262170 -1392 262226
rect -1820 262046 -1764 262102
rect -1696 262046 -1640 262102
rect -1572 262046 -1516 262102
rect -1448 262046 -1392 262102
rect -1820 261922 -1764 261978
rect -1696 261922 -1640 261978
rect -1572 261922 -1516 261978
rect -1448 261922 -1392 261978
rect -1820 244294 -1764 244350
rect -1696 244294 -1640 244350
rect -1572 244294 -1516 244350
rect -1448 244294 -1392 244350
rect -1820 244170 -1764 244226
rect -1696 244170 -1640 244226
rect -1572 244170 -1516 244226
rect -1448 244170 -1392 244226
rect -1820 244046 -1764 244102
rect -1696 244046 -1640 244102
rect -1572 244046 -1516 244102
rect -1448 244046 -1392 244102
rect -1820 243922 -1764 243978
rect -1696 243922 -1640 243978
rect -1572 243922 -1516 243978
rect -1448 243922 -1392 243978
rect -1820 226294 -1764 226350
rect -1696 226294 -1640 226350
rect -1572 226294 -1516 226350
rect -1448 226294 -1392 226350
rect -1820 226170 -1764 226226
rect -1696 226170 -1640 226226
rect -1572 226170 -1516 226226
rect -1448 226170 -1392 226226
rect -1820 226046 -1764 226102
rect -1696 226046 -1640 226102
rect -1572 226046 -1516 226102
rect -1448 226046 -1392 226102
rect -1820 225922 -1764 225978
rect -1696 225922 -1640 225978
rect -1572 225922 -1516 225978
rect -1448 225922 -1392 225978
rect -1820 208294 -1764 208350
rect -1696 208294 -1640 208350
rect -1572 208294 -1516 208350
rect -1448 208294 -1392 208350
rect -1820 208170 -1764 208226
rect -1696 208170 -1640 208226
rect -1572 208170 -1516 208226
rect -1448 208170 -1392 208226
rect -1820 208046 -1764 208102
rect -1696 208046 -1640 208102
rect -1572 208046 -1516 208102
rect -1448 208046 -1392 208102
rect -1820 207922 -1764 207978
rect -1696 207922 -1640 207978
rect -1572 207922 -1516 207978
rect -1448 207922 -1392 207978
rect -1820 190294 -1764 190350
rect -1696 190294 -1640 190350
rect -1572 190294 -1516 190350
rect -1448 190294 -1392 190350
rect -1820 190170 -1764 190226
rect -1696 190170 -1640 190226
rect -1572 190170 -1516 190226
rect -1448 190170 -1392 190226
rect -1820 190046 -1764 190102
rect -1696 190046 -1640 190102
rect -1572 190046 -1516 190102
rect -1448 190046 -1392 190102
rect -1820 189922 -1764 189978
rect -1696 189922 -1640 189978
rect -1572 189922 -1516 189978
rect -1448 189922 -1392 189978
rect -1820 172294 -1764 172350
rect -1696 172294 -1640 172350
rect -1572 172294 -1516 172350
rect -1448 172294 -1392 172350
rect -1820 172170 -1764 172226
rect -1696 172170 -1640 172226
rect -1572 172170 -1516 172226
rect -1448 172170 -1392 172226
rect -1820 172046 -1764 172102
rect -1696 172046 -1640 172102
rect -1572 172046 -1516 172102
rect -1448 172046 -1392 172102
rect -1820 171922 -1764 171978
rect -1696 171922 -1640 171978
rect -1572 171922 -1516 171978
rect -1448 171922 -1392 171978
rect -1820 154294 -1764 154350
rect -1696 154294 -1640 154350
rect -1572 154294 -1516 154350
rect -1448 154294 -1392 154350
rect -1820 154170 -1764 154226
rect -1696 154170 -1640 154226
rect -1572 154170 -1516 154226
rect -1448 154170 -1392 154226
rect -1820 154046 -1764 154102
rect -1696 154046 -1640 154102
rect -1572 154046 -1516 154102
rect -1448 154046 -1392 154102
rect -1820 153922 -1764 153978
rect -1696 153922 -1640 153978
rect -1572 153922 -1516 153978
rect -1448 153922 -1392 153978
rect -1820 136294 -1764 136350
rect -1696 136294 -1640 136350
rect -1572 136294 -1516 136350
rect -1448 136294 -1392 136350
rect -1820 136170 -1764 136226
rect -1696 136170 -1640 136226
rect -1572 136170 -1516 136226
rect -1448 136170 -1392 136226
rect -1820 136046 -1764 136102
rect -1696 136046 -1640 136102
rect -1572 136046 -1516 136102
rect -1448 136046 -1392 136102
rect -1820 135922 -1764 135978
rect -1696 135922 -1640 135978
rect -1572 135922 -1516 135978
rect -1448 135922 -1392 135978
rect -1820 118294 -1764 118350
rect -1696 118294 -1640 118350
rect -1572 118294 -1516 118350
rect -1448 118294 -1392 118350
rect -1820 118170 -1764 118226
rect -1696 118170 -1640 118226
rect -1572 118170 -1516 118226
rect -1448 118170 -1392 118226
rect -1820 118046 -1764 118102
rect -1696 118046 -1640 118102
rect -1572 118046 -1516 118102
rect -1448 118046 -1392 118102
rect -1820 117922 -1764 117978
rect -1696 117922 -1640 117978
rect -1572 117922 -1516 117978
rect -1448 117922 -1392 117978
rect -1820 100294 -1764 100350
rect -1696 100294 -1640 100350
rect -1572 100294 -1516 100350
rect -1448 100294 -1392 100350
rect -1820 100170 -1764 100226
rect -1696 100170 -1640 100226
rect -1572 100170 -1516 100226
rect -1448 100170 -1392 100226
rect -1820 100046 -1764 100102
rect -1696 100046 -1640 100102
rect -1572 100046 -1516 100102
rect -1448 100046 -1392 100102
rect -1820 99922 -1764 99978
rect -1696 99922 -1640 99978
rect -1572 99922 -1516 99978
rect -1448 99922 -1392 99978
rect -1820 82294 -1764 82350
rect -1696 82294 -1640 82350
rect -1572 82294 -1516 82350
rect -1448 82294 -1392 82350
rect -1820 82170 -1764 82226
rect -1696 82170 -1640 82226
rect -1572 82170 -1516 82226
rect -1448 82170 -1392 82226
rect -1820 82046 -1764 82102
rect -1696 82046 -1640 82102
rect -1572 82046 -1516 82102
rect -1448 82046 -1392 82102
rect -1820 81922 -1764 81978
rect -1696 81922 -1640 81978
rect -1572 81922 -1516 81978
rect -1448 81922 -1392 81978
rect -1820 64294 -1764 64350
rect -1696 64294 -1640 64350
rect -1572 64294 -1516 64350
rect -1448 64294 -1392 64350
rect -1820 64170 -1764 64226
rect -1696 64170 -1640 64226
rect -1572 64170 -1516 64226
rect -1448 64170 -1392 64226
rect -1820 64046 -1764 64102
rect -1696 64046 -1640 64102
rect -1572 64046 -1516 64102
rect -1448 64046 -1392 64102
rect -1820 63922 -1764 63978
rect -1696 63922 -1640 63978
rect -1572 63922 -1516 63978
rect -1448 63922 -1392 63978
rect -1820 46294 -1764 46350
rect -1696 46294 -1640 46350
rect -1572 46294 -1516 46350
rect -1448 46294 -1392 46350
rect -1820 46170 -1764 46226
rect -1696 46170 -1640 46226
rect -1572 46170 -1516 46226
rect -1448 46170 -1392 46226
rect -1820 46046 -1764 46102
rect -1696 46046 -1640 46102
rect -1572 46046 -1516 46102
rect -1448 46046 -1392 46102
rect -1820 45922 -1764 45978
rect -1696 45922 -1640 45978
rect -1572 45922 -1516 45978
rect -1448 45922 -1392 45978
rect -1820 28294 -1764 28350
rect -1696 28294 -1640 28350
rect -1572 28294 -1516 28350
rect -1448 28294 -1392 28350
rect -1820 28170 -1764 28226
rect -1696 28170 -1640 28226
rect -1572 28170 -1516 28226
rect -1448 28170 -1392 28226
rect -1820 28046 -1764 28102
rect -1696 28046 -1640 28102
rect -1572 28046 -1516 28102
rect -1448 28046 -1392 28102
rect -1820 27922 -1764 27978
rect -1696 27922 -1640 27978
rect -1572 27922 -1516 27978
rect -1448 27922 -1392 27978
rect -1820 10294 -1764 10350
rect -1696 10294 -1640 10350
rect -1572 10294 -1516 10350
rect -1448 10294 -1392 10350
rect -1820 10170 -1764 10226
rect -1696 10170 -1640 10226
rect -1572 10170 -1516 10226
rect -1448 10170 -1392 10226
rect -1820 10046 -1764 10102
rect -1696 10046 -1640 10102
rect -1572 10046 -1516 10102
rect -1448 10046 -1392 10102
rect -1820 9922 -1764 9978
rect -1696 9922 -1640 9978
rect -1572 9922 -1516 9978
rect -1448 9922 -1392 9978
rect -860 597156 -804 597212
rect -736 597156 -680 597212
rect -612 597156 -556 597212
rect -488 597156 -432 597212
rect -860 597032 -804 597088
rect -736 597032 -680 597088
rect -612 597032 -556 597088
rect -488 597032 -432 597088
rect -860 596908 -804 596964
rect -736 596908 -680 596964
rect -612 596908 -556 596964
rect -488 596908 -432 596964
rect -860 596784 -804 596840
rect -736 596784 -680 596840
rect -612 596784 -556 596840
rect -488 596784 -432 596840
rect -860 580294 -804 580350
rect -736 580294 -680 580350
rect -612 580294 -556 580350
rect -488 580294 -432 580350
rect -860 580170 -804 580226
rect -736 580170 -680 580226
rect -612 580170 -556 580226
rect -488 580170 -432 580226
rect -860 580046 -804 580102
rect -736 580046 -680 580102
rect -612 580046 -556 580102
rect -488 580046 -432 580102
rect -860 579922 -804 579978
rect -736 579922 -680 579978
rect -612 579922 -556 579978
rect -488 579922 -432 579978
rect -860 562294 -804 562350
rect -736 562294 -680 562350
rect -612 562294 -556 562350
rect -488 562294 -432 562350
rect -860 562170 -804 562226
rect -736 562170 -680 562226
rect -612 562170 -556 562226
rect -488 562170 -432 562226
rect -860 562046 -804 562102
rect -736 562046 -680 562102
rect -612 562046 -556 562102
rect -488 562046 -432 562102
rect -860 561922 -804 561978
rect -736 561922 -680 561978
rect -612 561922 -556 561978
rect -488 561922 -432 561978
rect -860 544294 -804 544350
rect -736 544294 -680 544350
rect -612 544294 -556 544350
rect -488 544294 -432 544350
rect -860 544170 -804 544226
rect -736 544170 -680 544226
rect -612 544170 -556 544226
rect -488 544170 -432 544226
rect -860 544046 -804 544102
rect -736 544046 -680 544102
rect -612 544046 -556 544102
rect -488 544046 -432 544102
rect -860 543922 -804 543978
rect -736 543922 -680 543978
rect -612 543922 -556 543978
rect -488 543922 -432 543978
rect -860 526294 -804 526350
rect -736 526294 -680 526350
rect -612 526294 -556 526350
rect -488 526294 -432 526350
rect -860 526170 -804 526226
rect -736 526170 -680 526226
rect -612 526170 -556 526226
rect -488 526170 -432 526226
rect -860 526046 -804 526102
rect -736 526046 -680 526102
rect -612 526046 -556 526102
rect -488 526046 -432 526102
rect -860 525922 -804 525978
rect -736 525922 -680 525978
rect -612 525922 -556 525978
rect -488 525922 -432 525978
rect -860 508294 -804 508350
rect -736 508294 -680 508350
rect -612 508294 -556 508350
rect -488 508294 -432 508350
rect -860 508170 -804 508226
rect -736 508170 -680 508226
rect -612 508170 -556 508226
rect -488 508170 -432 508226
rect -860 508046 -804 508102
rect -736 508046 -680 508102
rect -612 508046 -556 508102
rect -488 508046 -432 508102
rect -860 507922 -804 507978
rect -736 507922 -680 507978
rect -612 507922 -556 507978
rect -488 507922 -432 507978
rect -860 490294 -804 490350
rect -736 490294 -680 490350
rect -612 490294 -556 490350
rect -488 490294 -432 490350
rect -860 490170 -804 490226
rect -736 490170 -680 490226
rect -612 490170 -556 490226
rect -488 490170 -432 490226
rect -860 490046 -804 490102
rect -736 490046 -680 490102
rect -612 490046 -556 490102
rect -488 490046 -432 490102
rect -860 489922 -804 489978
rect -736 489922 -680 489978
rect -612 489922 -556 489978
rect -488 489922 -432 489978
rect -860 472294 -804 472350
rect -736 472294 -680 472350
rect -612 472294 -556 472350
rect -488 472294 -432 472350
rect -860 472170 -804 472226
rect -736 472170 -680 472226
rect -612 472170 -556 472226
rect -488 472170 -432 472226
rect -860 472046 -804 472102
rect -736 472046 -680 472102
rect -612 472046 -556 472102
rect -488 472046 -432 472102
rect -860 471922 -804 471978
rect -736 471922 -680 471978
rect -612 471922 -556 471978
rect -488 471922 -432 471978
rect -860 454294 -804 454350
rect -736 454294 -680 454350
rect -612 454294 -556 454350
rect -488 454294 -432 454350
rect -860 454170 -804 454226
rect -736 454170 -680 454226
rect -612 454170 -556 454226
rect -488 454170 -432 454226
rect -860 454046 -804 454102
rect -736 454046 -680 454102
rect -612 454046 -556 454102
rect -488 454046 -432 454102
rect -860 453922 -804 453978
rect -736 453922 -680 453978
rect -612 453922 -556 453978
rect -488 453922 -432 453978
rect -860 436294 -804 436350
rect -736 436294 -680 436350
rect -612 436294 -556 436350
rect -488 436294 -432 436350
rect -860 436170 -804 436226
rect -736 436170 -680 436226
rect -612 436170 -556 436226
rect -488 436170 -432 436226
rect -860 436046 -804 436102
rect -736 436046 -680 436102
rect -612 436046 -556 436102
rect -488 436046 -432 436102
rect -860 435922 -804 435978
rect -736 435922 -680 435978
rect -612 435922 -556 435978
rect -488 435922 -432 435978
rect -860 418294 -804 418350
rect -736 418294 -680 418350
rect -612 418294 -556 418350
rect -488 418294 -432 418350
rect -860 418170 -804 418226
rect -736 418170 -680 418226
rect -612 418170 -556 418226
rect -488 418170 -432 418226
rect -860 418046 -804 418102
rect -736 418046 -680 418102
rect -612 418046 -556 418102
rect -488 418046 -432 418102
rect -860 417922 -804 417978
rect -736 417922 -680 417978
rect -612 417922 -556 417978
rect -488 417922 -432 417978
rect -860 400294 -804 400350
rect -736 400294 -680 400350
rect -612 400294 -556 400350
rect -488 400294 -432 400350
rect -860 400170 -804 400226
rect -736 400170 -680 400226
rect -612 400170 -556 400226
rect -488 400170 -432 400226
rect -860 400046 -804 400102
rect -736 400046 -680 400102
rect -612 400046 -556 400102
rect -488 400046 -432 400102
rect -860 399922 -804 399978
rect -736 399922 -680 399978
rect -612 399922 -556 399978
rect -488 399922 -432 399978
rect -860 382294 -804 382350
rect -736 382294 -680 382350
rect -612 382294 -556 382350
rect -488 382294 -432 382350
rect -860 382170 -804 382226
rect -736 382170 -680 382226
rect -612 382170 -556 382226
rect -488 382170 -432 382226
rect -860 382046 -804 382102
rect -736 382046 -680 382102
rect -612 382046 -556 382102
rect -488 382046 -432 382102
rect -860 381922 -804 381978
rect -736 381922 -680 381978
rect -612 381922 -556 381978
rect -488 381922 -432 381978
rect -860 364294 -804 364350
rect -736 364294 -680 364350
rect -612 364294 -556 364350
rect -488 364294 -432 364350
rect -860 364170 -804 364226
rect -736 364170 -680 364226
rect -612 364170 -556 364226
rect -488 364170 -432 364226
rect -860 364046 -804 364102
rect -736 364046 -680 364102
rect -612 364046 -556 364102
rect -488 364046 -432 364102
rect -860 363922 -804 363978
rect -736 363922 -680 363978
rect -612 363922 -556 363978
rect -488 363922 -432 363978
rect -860 346294 -804 346350
rect -736 346294 -680 346350
rect -612 346294 -556 346350
rect -488 346294 -432 346350
rect -860 346170 -804 346226
rect -736 346170 -680 346226
rect -612 346170 -556 346226
rect -488 346170 -432 346226
rect -860 346046 -804 346102
rect -736 346046 -680 346102
rect -612 346046 -556 346102
rect -488 346046 -432 346102
rect -860 345922 -804 345978
rect -736 345922 -680 345978
rect -612 345922 -556 345978
rect -488 345922 -432 345978
rect -860 328294 -804 328350
rect -736 328294 -680 328350
rect -612 328294 -556 328350
rect -488 328294 -432 328350
rect -860 328170 -804 328226
rect -736 328170 -680 328226
rect -612 328170 -556 328226
rect -488 328170 -432 328226
rect -860 328046 -804 328102
rect -736 328046 -680 328102
rect -612 328046 -556 328102
rect -488 328046 -432 328102
rect -860 327922 -804 327978
rect -736 327922 -680 327978
rect -612 327922 -556 327978
rect -488 327922 -432 327978
rect -860 310294 -804 310350
rect -736 310294 -680 310350
rect -612 310294 -556 310350
rect -488 310294 -432 310350
rect -860 310170 -804 310226
rect -736 310170 -680 310226
rect -612 310170 -556 310226
rect -488 310170 -432 310226
rect -860 310046 -804 310102
rect -736 310046 -680 310102
rect -612 310046 -556 310102
rect -488 310046 -432 310102
rect -860 309922 -804 309978
rect -736 309922 -680 309978
rect -612 309922 -556 309978
rect -488 309922 -432 309978
rect -860 292294 -804 292350
rect -736 292294 -680 292350
rect -612 292294 -556 292350
rect -488 292294 -432 292350
rect -860 292170 -804 292226
rect -736 292170 -680 292226
rect -612 292170 -556 292226
rect -488 292170 -432 292226
rect -860 292046 -804 292102
rect -736 292046 -680 292102
rect -612 292046 -556 292102
rect -488 292046 -432 292102
rect -860 291922 -804 291978
rect -736 291922 -680 291978
rect -612 291922 -556 291978
rect -488 291922 -432 291978
rect -860 274294 -804 274350
rect -736 274294 -680 274350
rect -612 274294 -556 274350
rect -488 274294 -432 274350
rect -860 274170 -804 274226
rect -736 274170 -680 274226
rect -612 274170 -556 274226
rect -488 274170 -432 274226
rect -860 274046 -804 274102
rect -736 274046 -680 274102
rect -612 274046 -556 274102
rect -488 274046 -432 274102
rect -860 273922 -804 273978
rect -736 273922 -680 273978
rect -612 273922 -556 273978
rect -488 273922 -432 273978
rect -860 256294 -804 256350
rect -736 256294 -680 256350
rect -612 256294 -556 256350
rect -488 256294 -432 256350
rect -860 256170 -804 256226
rect -736 256170 -680 256226
rect -612 256170 -556 256226
rect -488 256170 -432 256226
rect -860 256046 -804 256102
rect -736 256046 -680 256102
rect -612 256046 -556 256102
rect -488 256046 -432 256102
rect -860 255922 -804 255978
rect -736 255922 -680 255978
rect -612 255922 -556 255978
rect -488 255922 -432 255978
rect -860 238294 -804 238350
rect -736 238294 -680 238350
rect -612 238294 -556 238350
rect -488 238294 -432 238350
rect -860 238170 -804 238226
rect -736 238170 -680 238226
rect -612 238170 -556 238226
rect -488 238170 -432 238226
rect -860 238046 -804 238102
rect -736 238046 -680 238102
rect -612 238046 -556 238102
rect -488 238046 -432 238102
rect -860 237922 -804 237978
rect -736 237922 -680 237978
rect -612 237922 -556 237978
rect -488 237922 -432 237978
rect -860 220294 -804 220350
rect -736 220294 -680 220350
rect -612 220294 -556 220350
rect -488 220294 -432 220350
rect -860 220170 -804 220226
rect -736 220170 -680 220226
rect -612 220170 -556 220226
rect -488 220170 -432 220226
rect -860 220046 -804 220102
rect -736 220046 -680 220102
rect -612 220046 -556 220102
rect -488 220046 -432 220102
rect -860 219922 -804 219978
rect -736 219922 -680 219978
rect -612 219922 -556 219978
rect -488 219922 -432 219978
rect -860 202294 -804 202350
rect -736 202294 -680 202350
rect -612 202294 -556 202350
rect -488 202294 -432 202350
rect -860 202170 -804 202226
rect -736 202170 -680 202226
rect -612 202170 -556 202226
rect -488 202170 -432 202226
rect -860 202046 -804 202102
rect -736 202046 -680 202102
rect -612 202046 -556 202102
rect -488 202046 -432 202102
rect -860 201922 -804 201978
rect -736 201922 -680 201978
rect -612 201922 -556 201978
rect -488 201922 -432 201978
rect -860 184294 -804 184350
rect -736 184294 -680 184350
rect -612 184294 -556 184350
rect -488 184294 -432 184350
rect -860 184170 -804 184226
rect -736 184170 -680 184226
rect -612 184170 -556 184226
rect -488 184170 -432 184226
rect -860 184046 -804 184102
rect -736 184046 -680 184102
rect -612 184046 -556 184102
rect -488 184046 -432 184102
rect -860 183922 -804 183978
rect -736 183922 -680 183978
rect -612 183922 -556 183978
rect -488 183922 -432 183978
rect -860 166294 -804 166350
rect -736 166294 -680 166350
rect -612 166294 -556 166350
rect -488 166294 -432 166350
rect -860 166170 -804 166226
rect -736 166170 -680 166226
rect -612 166170 -556 166226
rect -488 166170 -432 166226
rect -860 166046 -804 166102
rect -736 166046 -680 166102
rect -612 166046 -556 166102
rect -488 166046 -432 166102
rect -860 165922 -804 165978
rect -736 165922 -680 165978
rect -612 165922 -556 165978
rect -488 165922 -432 165978
rect -860 148294 -804 148350
rect -736 148294 -680 148350
rect -612 148294 -556 148350
rect -488 148294 -432 148350
rect -860 148170 -804 148226
rect -736 148170 -680 148226
rect -612 148170 -556 148226
rect -488 148170 -432 148226
rect -860 148046 -804 148102
rect -736 148046 -680 148102
rect -612 148046 -556 148102
rect -488 148046 -432 148102
rect -860 147922 -804 147978
rect -736 147922 -680 147978
rect -612 147922 -556 147978
rect -488 147922 -432 147978
rect -860 130294 -804 130350
rect -736 130294 -680 130350
rect -612 130294 -556 130350
rect -488 130294 -432 130350
rect -860 130170 -804 130226
rect -736 130170 -680 130226
rect -612 130170 -556 130226
rect -488 130170 -432 130226
rect -860 130046 -804 130102
rect -736 130046 -680 130102
rect -612 130046 -556 130102
rect -488 130046 -432 130102
rect -860 129922 -804 129978
rect -736 129922 -680 129978
rect -612 129922 -556 129978
rect -488 129922 -432 129978
rect -860 112294 -804 112350
rect -736 112294 -680 112350
rect -612 112294 -556 112350
rect -488 112294 -432 112350
rect -860 112170 -804 112226
rect -736 112170 -680 112226
rect -612 112170 -556 112226
rect -488 112170 -432 112226
rect -860 112046 -804 112102
rect -736 112046 -680 112102
rect -612 112046 -556 112102
rect -488 112046 -432 112102
rect -860 111922 -804 111978
rect -736 111922 -680 111978
rect -612 111922 -556 111978
rect -488 111922 -432 111978
rect -860 94294 -804 94350
rect -736 94294 -680 94350
rect -612 94294 -556 94350
rect -488 94294 -432 94350
rect -860 94170 -804 94226
rect -736 94170 -680 94226
rect -612 94170 -556 94226
rect -488 94170 -432 94226
rect -860 94046 -804 94102
rect -736 94046 -680 94102
rect -612 94046 -556 94102
rect -488 94046 -432 94102
rect -860 93922 -804 93978
rect -736 93922 -680 93978
rect -612 93922 -556 93978
rect -488 93922 -432 93978
rect -860 76294 -804 76350
rect -736 76294 -680 76350
rect -612 76294 -556 76350
rect -488 76294 -432 76350
rect -860 76170 -804 76226
rect -736 76170 -680 76226
rect -612 76170 -556 76226
rect -488 76170 -432 76226
rect -860 76046 -804 76102
rect -736 76046 -680 76102
rect -612 76046 -556 76102
rect -488 76046 -432 76102
rect -860 75922 -804 75978
rect -736 75922 -680 75978
rect -612 75922 -556 75978
rect -488 75922 -432 75978
rect -860 58294 -804 58350
rect -736 58294 -680 58350
rect -612 58294 -556 58350
rect -488 58294 -432 58350
rect -860 58170 -804 58226
rect -736 58170 -680 58226
rect -612 58170 -556 58226
rect -488 58170 -432 58226
rect -860 58046 -804 58102
rect -736 58046 -680 58102
rect -612 58046 -556 58102
rect -488 58046 -432 58102
rect -860 57922 -804 57978
rect -736 57922 -680 57978
rect -612 57922 -556 57978
rect -488 57922 -432 57978
rect -860 40294 -804 40350
rect -736 40294 -680 40350
rect -612 40294 -556 40350
rect -488 40294 -432 40350
rect -860 40170 -804 40226
rect -736 40170 -680 40226
rect -612 40170 -556 40226
rect -488 40170 -432 40226
rect -860 40046 -804 40102
rect -736 40046 -680 40102
rect -612 40046 -556 40102
rect -488 40046 -432 40102
rect -860 39922 -804 39978
rect -736 39922 -680 39978
rect -612 39922 -556 39978
rect -488 39922 -432 39978
rect -860 22294 -804 22350
rect -736 22294 -680 22350
rect -612 22294 -556 22350
rect -488 22294 -432 22350
rect -860 22170 -804 22226
rect -736 22170 -680 22226
rect -612 22170 -556 22226
rect -488 22170 -432 22226
rect -860 22046 -804 22102
rect -736 22046 -680 22102
rect -612 22046 -556 22102
rect -488 22046 -432 22102
rect -860 21922 -804 21978
rect -736 21922 -680 21978
rect -612 21922 -556 21978
rect -488 21922 -432 21978
rect -860 4294 -804 4350
rect -736 4294 -680 4350
rect -612 4294 -556 4350
rect -488 4294 -432 4350
rect -860 4170 -804 4226
rect -736 4170 -680 4226
rect -612 4170 -556 4226
rect -488 4170 -432 4226
rect -860 4046 -804 4102
rect -736 4046 -680 4102
rect -612 4046 -556 4102
rect -488 4046 -432 4102
rect -860 3922 -804 3978
rect -736 3922 -680 3978
rect -612 3922 -556 3978
rect -488 3922 -432 3978
rect -860 -216 -804 -160
rect -736 -216 -680 -160
rect -612 -216 -556 -160
rect -488 -216 -432 -160
rect -860 -340 -804 -284
rect -736 -340 -680 -284
rect -612 -340 -556 -284
rect -488 -340 -432 -284
rect -860 -464 -804 -408
rect -736 -464 -680 -408
rect -612 -464 -556 -408
rect -488 -464 -432 -408
rect -860 -588 -804 -532
rect -736 -588 -680 -532
rect -612 -588 -556 -532
rect -488 -588 -432 -532
rect 3250 597156 3306 597212
rect 3374 597156 3430 597212
rect 3498 597156 3554 597212
rect 3622 597156 3678 597212
rect 3250 597032 3306 597088
rect 3374 597032 3430 597088
rect 3498 597032 3554 597088
rect 3622 597032 3678 597088
rect 3250 596908 3306 596964
rect 3374 596908 3430 596964
rect 3498 596908 3554 596964
rect 3622 596908 3678 596964
rect 3250 596784 3306 596840
rect 3374 596784 3430 596840
rect 3498 596784 3554 596840
rect 3622 596784 3678 596840
rect 3250 580294 3306 580350
rect 3374 580294 3430 580350
rect 3498 580294 3554 580350
rect 3622 580294 3678 580350
rect 3250 580170 3306 580226
rect 3374 580170 3430 580226
rect 3498 580170 3554 580226
rect 3622 580170 3678 580226
rect 3250 580046 3306 580102
rect 3374 580046 3430 580102
rect 3498 580046 3554 580102
rect 3622 580046 3678 580102
rect 3250 579922 3306 579978
rect 3374 579922 3430 579978
rect 3498 579922 3554 579978
rect 3622 579922 3678 579978
rect 3250 562294 3306 562350
rect 3374 562294 3430 562350
rect 3498 562294 3554 562350
rect 3622 562294 3678 562350
rect 3250 562170 3306 562226
rect 3374 562170 3430 562226
rect 3498 562170 3554 562226
rect 3622 562170 3678 562226
rect 3250 562046 3306 562102
rect 3374 562046 3430 562102
rect 3498 562046 3554 562102
rect 3622 562046 3678 562102
rect 3250 561922 3306 561978
rect 3374 561922 3430 561978
rect 3498 561922 3554 561978
rect 3622 561922 3678 561978
rect 6970 598116 7026 598172
rect 7094 598116 7150 598172
rect 7218 598116 7274 598172
rect 7342 598116 7398 598172
rect 6970 597992 7026 598048
rect 7094 597992 7150 598048
rect 7218 597992 7274 598048
rect 7342 597992 7398 598048
rect 6970 597868 7026 597924
rect 7094 597868 7150 597924
rect 7218 597868 7274 597924
rect 7342 597868 7398 597924
rect 6970 597744 7026 597800
rect 7094 597744 7150 597800
rect 7218 597744 7274 597800
rect 7342 597744 7398 597800
rect 6970 586294 7026 586350
rect 7094 586294 7150 586350
rect 7218 586294 7274 586350
rect 7342 586294 7398 586350
rect 6970 586170 7026 586226
rect 7094 586170 7150 586226
rect 7218 586170 7274 586226
rect 7342 586170 7398 586226
rect 6970 586046 7026 586102
rect 7094 586046 7150 586102
rect 7218 586046 7274 586102
rect 7342 586046 7398 586102
rect 6970 585922 7026 585978
rect 7094 585922 7150 585978
rect 7218 585922 7274 585978
rect 7342 585922 7398 585978
rect 6970 568294 7026 568350
rect 7094 568294 7150 568350
rect 7218 568294 7274 568350
rect 7342 568294 7398 568350
rect 6970 568170 7026 568226
rect 7094 568170 7150 568226
rect 7218 568170 7274 568226
rect 7342 568170 7398 568226
rect 6970 568046 7026 568102
rect 7094 568046 7150 568102
rect 7218 568046 7274 568102
rect 7342 568046 7398 568102
rect 6970 567922 7026 567978
rect 7094 567922 7150 567978
rect 7218 567922 7274 567978
rect 7342 567922 7398 567978
rect 6970 550294 7026 550350
rect 7094 550294 7150 550350
rect 7218 550294 7274 550350
rect 7342 550294 7398 550350
rect 6970 550170 7026 550226
rect 7094 550170 7150 550226
rect 7218 550170 7274 550226
rect 7342 550170 7398 550226
rect 6970 550046 7026 550102
rect 7094 550046 7150 550102
rect 7218 550046 7274 550102
rect 7342 550046 7398 550102
rect 6970 549922 7026 549978
rect 7094 549922 7150 549978
rect 7218 549922 7274 549978
rect 7342 549922 7398 549978
rect 3250 544294 3306 544350
rect 3374 544294 3430 544350
rect 3498 544294 3554 544350
rect 3622 544294 3678 544350
rect 3250 544170 3306 544226
rect 3374 544170 3430 544226
rect 3498 544170 3554 544226
rect 3622 544170 3678 544226
rect 3250 544046 3306 544102
rect 3374 544046 3430 544102
rect 3498 544046 3554 544102
rect 3622 544046 3678 544102
rect 3250 543922 3306 543978
rect 3374 543922 3430 543978
rect 3498 543922 3554 543978
rect 3622 543922 3678 543978
rect 3250 526294 3306 526350
rect 3374 526294 3430 526350
rect 3498 526294 3554 526350
rect 3622 526294 3678 526350
rect 3250 526170 3306 526226
rect 3374 526170 3430 526226
rect 3498 526170 3554 526226
rect 3622 526170 3678 526226
rect 3250 526046 3306 526102
rect 3374 526046 3430 526102
rect 3498 526046 3554 526102
rect 3622 526046 3678 526102
rect 3250 525922 3306 525978
rect 3374 525922 3430 525978
rect 3498 525922 3554 525978
rect 3622 525922 3678 525978
rect 3250 508294 3306 508350
rect 3374 508294 3430 508350
rect 3498 508294 3554 508350
rect 3622 508294 3678 508350
rect 3250 508170 3306 508226
rect 3374 508170 3430 508226
rect 3498 508170 3554 508226
rect 3622 508170 3678 508226
rect 3250 508046 3306 508102
rect 3374 508046 3430 508102
rect 3498 508046 3554 508102
rect 3622 508046 3678 508102
rect 3250 507922 3306 507978
rect 3374 507922 3430 507978
rect 3498 507922 3554 507978
rect 3622 507922 3678 507978
rect 3250 490294 3306 490350
rect 3374 490294 3430 490350
rect 3498 490294 3554 490350
rect 3622 490294 3678 490350
rect 3250 490170 3306 490226
rect 3374 490170 3430 490226
rect 3498 490170 3554 490226
rect 3622 490170 3678 490226
rect 3250 490046 3306 490102
rect 3374 490046 3430 490102
rect 3498 490046 3554 490102
rect 3622 490046 3678 490102
rect 3250 489922 3306 489978
rect 3374 489922 3430 489978
rect 3498 489922 3554 489978
rect 3622 489922 3678 489978
rect 3250 472294 3306 472350
rect 3374 472294 3430 472350
rect 3498 472294 3554 472350
rect 3622 472294 3678 472350
rect 3250 472170 3306 472226
rect 3374 472170 3430 472226
rect 3498 472170 3554 472226
rect 3622 472170 3678 472226
rect 3250 472046 3306 472102
rect 3374 472046 3430 472102
rect 3498 472046 3554 472102
rect 3622 472046 3678 472102
rect 3250 471922 3306 471978
rect 3374 471922 3430 471978
rect 3498 471922 3554 471978
rect 3622 471922 3678 471978
rect 3250 454294 3306 454350
rect 3374 454294 3430 454350
rect 3498 454294 3554 454350
rect 3622 454294 3678 454350
rect 3250 454170 3306 454226
rect 3374 454170 3430 454226
rect 3498 454170 3554 454226
rect 3622 454170 3678 454226
rect 3250 454046 3306 454102
rect 3374 454046 3430 454102
rect 3498 454046 3554 454102
rect 3622 454046 3678 454102
rect 3250 453922 3306 453978
rect 3374 453922 3430 453978
rect 3498 453922 3554 453978
rect 3622 453922 3678 453978
rect 3250 436294 3306 436350
rect 3374 436294 3430 436350
rect 3498 436294 3554 436350
rect 3622 436294 3678 436350
rect 3250 436170 3306 436226
rect 3374 436170 3430 436226
rect 3498 436170 3554 436226
rect 3622 436170 3678 436226
rect 3250 436046 3306 436102
rect 3374 436046 3430 436102
rect 3498 436046 3554 436102
rect 3622 436046 3678 436102
rect 3250 435922 3306 435978
rect 3374 435922 3430 435978
rect 3498 435922 3554 435978
rect 3622 435922 3678 435978
rect 3250 418294 3306 418350
rect 3374 418294 3430 418350
rect 3498 418294 3554 418350
rect 3622 418294 3678 418350
rect 3250 418170 3306 418226
rect 3374 418170 3430 418226
rect 3498 418170 3554 418226
rect 3622 418170 3678 418226
rect 3250 418046 3306 418102
rect 3374 418046 3430 418102
rect 3498 418046 3554 418102
rect 3622 418046 3678 418102
rect 3250 417922 3306 417978
rect 3374 417922 3430 417978
rect 3498 417922 3554 417978
rect 3622 417922 3678 417978
rect 3250 400294 3306 400350
rect 3374 400294 3430 400350
rect 3498 400294 3554 400350
rect 3622 400294 3678 400350
rect 3250 400170 3306 400226
rect 3374 400170 3430 400226
rect 3498 400170 3554 400226
rect 3622 400170 3678 400226
rect 3250 400046 3306 400102
rect 3374 400046 3430 400102
rect 3498 400046 3554 400102
rect 3622 400046 3678 400102
rect 3250 399922 3306 399978
rect 3374 399922 3430 399978
rect 3498 399922 3554 399978
rect 3622 399922 3678 399978
rect 3250 382294 3306 382350
rect 3374 382294 3430 382350
rect 3498 382294 3554 382350
rect 3622 382294 3678 382350
rect 3250 382170 3306 382226
rect 3374 382170 3430 382226
rect 3498 382170 3554 382226
rect 3622 382170 3678 382226
rect 3250 382046 3306 382102
rect 3374 382046 3430 382102
rect 3498 382046 3554 382102
rect 3622 382046 3678 382102
rect 3250 381922 3306 381978
rect 3374 381922 3430 381978
rect 3498 381922 3554 381978
rect 3622 381922 3678 381978
rect 3250 364294 3306 364350
rect 3374 364294 3430 364350
rect 3498 364294 3554 364350
rect 3622 364294 3678 364350
rect 3250 364170 3306 364226
rect 3374 364170 3430 364226
rect 3498 364170 3554 364226
rect 3622 364170 3678 364226
rect 3250 364046 3306 364102
rect 3374 364046 3430 364102
rect 3498 364046 3554 364102
rect 3622 364046 3678 364102
rect 3250 363922 3306 363978
rect 3374 363922 3430 363978
rect 3498 363922 3554 363978
rect 3622 363922 3678 363978
rect 3250 346294 3306 346350
rect 3374 346294 3430 346350
rect 3498 346294 3554 346350
rect 3622 346294 3678 346350
rect 3250 346170 3306 346226
rect 3374 346170 3430 346226
rect 3498 346170 3554 346226
rect 3622 346170 3678 346226
rect 3250 346046 3306 346102
rect 3374 346046 3430 346102
rect 3498 346046 3554 346102
rect 3622 346046 3678 346102
rect 3250 345922 3306 345978
rect 3374 345922 3430 345978
rect 3498 345922 3554 345978
rect 3622 345922 3678 345978
rect 3250 328294 3306 328350
rect 3374 328294 3430 328350
rect 3498 328294 3554 328350
rect 3622 328294 3678 328350
rect 3250 328170 3306 328226
rect 3374 328170 3430 328226
rect 3498 328170 3554 328226
rect 3622 328170 3678 328226
rect 3250 328046 3306 328102
rect 3374 328046 3430 328102
rect 3498 328046 3554 328102
rect 3622 328046 3678 328102
rect 3250 327922 3306 327978
rect 3374 327922 3430 327978
rect 3498 327922 3554 327978
rect 3622 327922 3678 327978
rect 3250 310294 3306 310350
rect 3374 310294 3430 310350
rect 3498 310294 3554 310350
rect 3622 310294 3678 310350
rect 3250 310170 3306 310226
rect 3374 310170 3430 310226
rect 3498 310170 3554 310226
rect 3622 310170 3678 310226
rect 3250 310046 3306 310102
rect 3374 310046 3430 310102
rect 3498 310046 3554 310102
rect 3622 310046 3678 310102
rect 3250 309922 3306 309978
rect 3374 309922 3430 309978
rect 3498 309922 3554 309978
rect 3622 309922 3678 309978
rect 3250 292294 3306 292350
rect 3374 292294 3430 292350
rect 3498 292294 3554 292350
rect 3622 292294 3678 292350
rect 3250 292170 3306 292226
rect 3374 292170 3430 292226
rect 3498 292170 3554 292226
rect 3622 292170 3678 292226
rect 3250 292046 3306 292102
rect 3374 292046 3430 292102
rect 3498 292046 3554 292102
rect 3622 292046 3678 292102
rect 3250 291922 3306 291978
rect 3374 291922 3430 291978
rect 3498 291922 3554 291978
rect 3622 291922 3678 291978
rect 3250 274294 3306 274350
rect 3374 274294 3430 274350
rect 3498 274294 3554 274350
rect 3622 274294 3678 274350
rect 3250 274170 3306 274226
rect 3374 274170 3430 274226
rect 3498 274170 3554 274226
rect 3622 274170 3678 274226
rect 3250 274046 3306 274102
rect 3374 274046 3430 274102
rect 3498 274046 3554 274102
rect 3622 274046 3678 274102
rect 3250 273922 3306 273978
rect 3374 273922 3430 273978
rect 3498 273922 3554 273978
rect 3622 273922 3678 273978
rect 3250 256294 3306 256350
rect 3374 256294 3430 256350
rect 3498 256294 3554 256350
rect 3622 256294 3678 256350
rect 3250 256170 3306 256226
rect 3374 256170 3430 256226
rect 3498 256170 3554 256226
rect 3622 256170 3678 256226
rect 3250 256046 3306 256102
rect 3374 256046 3430 256102
rect 3498 256046 3554 256102
rect 3622 256046 3678 256102
rect 3250 255922 3306 255978
rect 3374 255922 3430 255978
rect 3498 255922 3554 255978
rect 3622 255922 3678 255978
rect 3250 238294 3306 238350
rect 3374 238294 3430 238350
rect 3498 238294 3554 238350
rect 3622 238294 3678 238350
rect 3250 238170 3306 238226
rect 3374 238170 3430 238226
rect 3498 238170 3554 238226
rect 3622 238170 3678 238226
rect 3250 238046 3306 238102
rect 3374 238046 3430 238102
rect 3498 238046 3554 238102
rect 3622 238046 3678 238102
rect 3250 237922 3306 237978
rect 3374 237922 3430 237978
rect 3498 237922 3554 237978
rect 3622 237922 3678 237978
rect 3250 220294 3306 220350
rect 3374 220294 3430 220350
rect 3498 220294 3554 220350
rect 3622 220294 3678 220350
rect 3250 220170 3306 220226
rect 3374 220170 3430 220226
rect 3498 220170 3554 220226
rect 3622 220170 3678 220226
rect 3250 220046 3306 220102
rect 3374 220046 3430 220102
rect 3498 220046 3554 220102
rect 3622 220046 3678 220102
rect 3250 219922 3306 219978
rect 3374 219922 3430 219978
rect 3498 219922 3554 219978
rect 3622 219922 3678 219978
rect 3250 202294 3306 202350
rect 3374 202294 3430 202350
rect 3498 202294 3554 202350
rect 3622 202294 3678 202350
rect 3250 202170 3306 202226
rect 3374 202170 3430 202226
rect 3498 202170 3554 202226
rect 3622 202170 3678 202226
rect 3250 202046 3306 202102
rect 3374 202046 3430 202102
rect 3498 202046 3554 202102
rect 3622 202046 3678 202102
rect 3250 201922 3306 201978
rect 3374 201922 3430 201978
rect 3498 201922 3554 201978
rect 3622 201922 3678 201978
rect 3250 184294 3306 184350
rect 3374 184294 3430 184350
rect 3498 184294 3554 184350
rect 3622 184294 3678 184350
rect 3250 184170 3306 184226
rect 3374 184170 3430 184226
rect 3498 184170 3554 184226
rect 3622 184170 3678 184226
rect 3250 184046 3306 184102
rect 3374 184046 3430 184102
rect 3498 184046 3554 184102
rect 3622 184046 3678 184102
rect 3250 183922 3306 183978
rect 3374 183922 3430 183978
rect 3498 183922 3554 183978
rect 3622 183922 3678 183978
rect 3250 166294 3306 166350
rect 3374 166294 3430 166350
rect 3498 166294 3554 166350
rect 3622 166294 3678 166350
rect 3250 166170 3306 166226
rect 3374 166170 3430 166226
rect 3498 166170 3554 166226
rect 3622 166170 3678 166226
rect 3250 166046 3306 166102
rect 3374 166046 3430 166102
rect 3498 166046 3554 166102
rect 3622 166046 3678 166102
rect 3250 165922 3306 165978
rect 3374 165922 3430 165978
rect 3498 165922 3554 165978
rect 3622 165922 3678 165978
rect 3250 148294 3306 148350
rect 3374 148294 3430 148350
rect 3498 148294 3554 148350
rect 3622 148294 3678 148350
rect 3250 148170 3306 148226
rect 3374 148170 3430 148226
rect 3498 148170 3554 148226
rect 3622 148170 3678 148226
rect 3250 148046 3306 148102
rect 3374 148046 3430 148102
rect 3498 148046 3554 148102
rect 3622 148046 3678 148102
rect 3250 147922 3306 147978
rect 3374 147922 3430 147978
rect 3498 147922 3554 147978
rect 3622 147922 3678 147978
rect 3250 130294 3306 130350
rect 3374 130294 3430 130350
rect 3498 130294 3554 130350
rect 3622 130294 3678 130350
rect 3250 130170 3306 130226
rect 3374 130170 3430 130226
rect 3498 130170 3554 130226
rect 3622 130170 3678 130226
rect 3250 130046 3306 130102
rect 3374 130046 3430 130102
rect 3498 130046 3554 130102
rect 3622 130046 3678 130102
rect 3250 129922 3306 129978
rect 3374 129922 3430 129978
rect 3498 129922 3554 129978
rect 3622 129922 3678 129978
rect 3250 112294 3306 112350
rect 3374 112294 3430 112350
rect 3498 112294 3554 112350
rect 3622 112294 3678 112350
rect 3250 112170 3306 112226
rect 3374 112170 3430 112226
rect 3498 112170 3554 112226
rect 3622 112170 3678 112226
rect 3250 112046 3306 112102
rect 3374 112046 3430 112102
rect 3498 112046 3554 112102
rect 3622 112046 3678 112102
rect 3250 111922 3306 111978
rect 3374 111922 3430 111978
rect 3498 111922 3554 111978
rect 3622 111922 3678 111978
rect 3250 94294 3306 94350
rect 3374 94294 3430 94350
rect 3498 94294 3554 94350
rect 3622 94294 3678 94350
rect 3250 94170 3306 94226
rect 3374 94170 3430 94226
rect 3498 94170 3554 94226
rect 3622 94170 3678 94226
rect 3250 94046 3306 94102
rect 3374 94046 3430 94102
rect 3498 94046 3554 94102
rect 3622 94046 3678 94102
rect 3250 93922 3306 93978
rect 3374 93922 3430 93978
rect 3498 93922 3554 93978
rect 3622 93922 3678 93978
rect 3250 76294 3306 76350
rect 3374 76294 3430 76350
rect 3498 76294 3554 76350
rect 3622 76294 3678 76350
rect 3250 76170 3306 76226
rect 3374 76170 3430 76226
rect 3498 76170 3554 76226
rect 3622 76170 3678 76226
rect 3250 76046 3306 76102
rect 3374 76046 3430 76102
rect 3498 76046 3554 76102
rect 3622 76046 3678 76102
rect 3250 75922 3306 75978
rect 3374 75922 3430 75978
rect 3498 75922 3554 75978
rect 3622 75922 3678 75978
rect 3250 58294 3306 58350
rect 3374 58294 3430 58350
rect 3498 58294 3554 58350
rect 3622 58294 3678 58350
rect 3250 58170 3306 58226
rect 3374 58170 3430 58226
rect 3498 58170 3554 58226
rect 3622 58170 3678 58226
rect 3250 58046 3306 58102
rect 3374 58046 3430 58102
rect 3498 58046 3554 58102
rect 3622 58046 3678 58102
rect 3250 57922 3306 57978
rect 3374 57922 3430 57978
rect 3498 57922 3554 57978
rect 3622 57922 3678 57978
rect 6970 532294 7026 532350
rect 7094 532294 7150 532350
rect 7218 532294 7274 532350
rect 7342 532294 7398 532350
rect 6970 532170 7026 532226
rect 7094 532170 7150 532226
rect 7218 532170 7274 532226
rect 7342 532170 7398 532226
rect 6970 532046 7026 532102
rect 7094 532046 7150 532102
rect 7218 532046 7274 532102
rect 7342 532046 7398 532102
rect 6970 531922 7026 531978
rect 7094 531922 7150 531978
rect 7218 531922 7274 531978
rect 7342 531922 7398 531978
rect 6970 514294 7026 514350
rect 7094 514294 7150 514350
rect 7218 514294 7274 514350
rect 7342 514294 7398 514350
rect 6970 514170 7026 514226
rect 7094 514170 7150 514226
rect 7218 514170 7274 514226
rect 7342 514170 7398 514226
rect 6970 514046 7026 514102
rect 7094 514046 7150 514102
rect 7218 514046 7274 514102
rect 7342 514046 7398 514102
rect 6970 513922 7026 513978
rect 7094 513922 7150 513978
rect 7218 513922 7274 513978
rect 7342 513922 7398 513978
rect 21250 597156 21306 597212
rect 21374 597156 21430 597212
rect 21498 597156 21554 597212
rect 21622 597156 21678 597212
rect 21250 597032 21306 597088
rect 21374 597032 21430 597088
rect 21498 597032 21554 597088
rect 21622 597032 21678 597088
rect 21250 596908 21306 596964
rect 21374 596908 21430 596964
rect 21498 596908 21554 596964
rect 21622 596908 21678 596964
rect 21250 596784 21306 596840
rect 21374 596784 21430 596840
rect 21498 596784 21554 596840
rect 21622 596784 21678 596840
rect 21250 580294 21306 580350
rect 21374 580294 21430 580350
rect 21498 580294 21554 580350
rect 21622 580294 21678 580350
rect 21250 580170 21306 580226
rect 21374 580170 21430 580226
rect 21498 580170 21554 580226
rect 21622 580170 21678 580226
rect 21250 580046 21306 580102
rect 21374 580046 21430 580102
rect 21498 580046 21554 580102
rect 21622 580046 21678 580102
rect 21250 579922 21306 579978
rect 21374 579922 21430 579978
rect 21498 579922 21554 579978
rect 21622 579922 21678 579978
rect 21250 562294 21306 562350
rect 21374 562294 21430 562350
rect 21498 562294 21554 562350
rect 21622 562294 21678 562350
rect 21250 562170 21306 562226
rect 21374 562170 21430 562226
rect 21498 562170 21554 562226
rect 21622 562170 21678 562226
rect 21250 562046 21306 562102
rect 21374 562046 21430 562102
rect 21498 562046 21554 562102
rect 21622 562046 21678 562102
rect 21250 561922 21306 561978
rect 21374 561922 21430 561978
rect 21498 561922 21554 561978
rect 21622 561922 21678 561978
rect 21250 544294 21306 544350
rect 21374 544294 21430 544350
rect 21498 544294 21554 544350
rect 21622 544294 21678 544350
rect 21250 544170 21306 544226
rect 21374 544170 21430 544226
rect 21498 544170 21554 544226
rect 21622 544170 21678 544226
rect 21250 544046 21306 544102
rect 21374 544046 21430 544102
rect 21498 544046 21554 544102
rect 21622 544046 21678 544102
rect 21250 543922 21306 543978
rect 21374 543922 21430 543978
rect 21498 543922 21554 543978
rect 21622 543922 21678 543978
rect 24970 598116 25026 598172
rect 25094 598116 25150 598172
rect 25218 598116 25274 598172
rect 25342 598116 25398 598172
rect 24970 597992 25026 598048
rect 25094 597992 25150 598048
rect 25218 597992 25274 598048
rect 25342 597992 25398 598048
rect 24970 597868 25026 597924
rect 25094 597868 25150 597924
rect 25218 597868 25274 597924
rect 25342 597868 25398 597924
rect 24970 597744 25026 597800
rect 25094 597744 25150 597800
rect 25218 597744 25274 597800
rect 25342 597744 25398 597800
rect 39250 597156 39306 597212
rect 39374 597156 39430 597212
rect 39498 597156 39554 597212
rect 39622 597156 39678 597212
rect 39250 597032 39306 597088
rect 39374 597032 39430 597088
rect 39498 597032 39554 597088
rect 39622 597032 39678 597088
rect 39250 596908 39306 596964
rect 39374 596908 39430 596964
rect 39498 596908 39554 596964
rect 39622 596908 39678 596964
rect 39250 596784 39306 596840
rect 39374 596784 39430 596840
rect 39498 596784 39554 596840
rect 39622 596784 39678 596840
rect 24970 586294 25026 586350
rect 25094 586294 25150 586350
rect 25218 586294 25274 586350
rect 25342 586294 25398 586350
rect 24970 586170 25026 586226
rect 25094 586170 25150 586226
rect 25218 586170 25274 586226
rect 25342 586170 25398 586226
rect 24970 586046 25026 586102
rect 25094 586046 25150 586102
rect 25218 586046 25274 586102
rect 25342 586046 25398 586102
rect 24970 585922 25026 585978
rect 25094 585922 25150 585978
rect 25218 585922 25274 585978
rect 25342 585922 25398 585978
rect 24970 568294 25026 568350
rect 25094 568294 25150 568350
rect 25218 568294 25274 568350
rect 25342 568294 25398 568350
rect 24970 568170 25026 568226
rect 25094 568170 25150 568226
rect 25218 568170 25274 568226
rect 25342 568170 25398 568226
rect 24970 568046 25026 568102
rect 25094 568046 25150 568102
rect 25218 568046 25274 568102
rect 25342 568046 25398 568102
rect 24970 567922 25026 567978
rect 25094 567922 25150 567978
rect 25218 567922 25274 567978
rect 25342 567922 25398 567978
rect 24970 550294 25026 550350
rect 25094 550294 25150 550350
rect 25218 550294 25274 550350
rect 25342 550294 25398 550350
rect 24970 550170 25026 550226
rect 25094 550170 25150 550226
rect 25218 550170 25274 550226
rect 25342 550170 25398 550226
rect 24970 550046 25026 550102
rect 25094 550046 25150 550102
rect 25218 550046 25274 550102
rect 25342 550046 25398 550102
rect 24970 549922 25026 549978
rect 25094 549922 25150 549978
rect 25218 549922 25274 549978
rect 25342 549922 25398 549978
rect 24970 532294 25026 532350
rect 25094 532294 25150 532350
rect 25218 532294 25274 532350
rect 25342 532294 25398 532350
rect 24970 532170 25026 532226
rect 25094 532170 25150 532226
rect 25218 532170 25274 532226
rect 25342 532170 25398 532226
rect 24970 532046 25026 532102
rect 25094 532046 25150 532102
rect 25218 532046 25274 532102
rect 25342 532046 25398 532102
rect 24970 531922 25026 531978
rect 25094 531922 25150 531978
rect 25218 531922 25274 531978
rect 25342 531922 25398 531978
rect 21250 526294 21306 526350
rect 21374 526294 21430 526350
rect 21498 526294 21554 526350
rect 21622 526294 21678 526350
rect 21250 526170 21306 526226
rect 21374 526170 21430 526226
rect 21498 526170 21554 526226
rect 21622 526170 21678 526226
rect 21250 526046 21306 526102
rect 21374 526046 21430 526102
rect 21498 526046 21554 526102
rect 21622 526046 21678 526102
rect 21250 525922 21306 525978
rect 21374 525922 21430 525978
rect 21498 525922 21554 525978
rect 21622 525922 21678 525978
rect 21250 508294 21306 508350
rect 21374 508294 21430 508350
rect 21498 508294 21554 508350
rect 21622 508294 21678 508350
rect 21250 508170 21306 508226
rect 21374 508170 21430 508226
rect 21498 508170 21554 508226
rect 21622 508170 21678 508226
rect 21250 508046 21306 508102
rect 21374 508046 21430 508102
rect 21498 508046 21554 508102
rect 21622 508046 21678 508102
rect 21250 507922 21306 507978
rect 21374 507922 21430 507978
rect 21498 507922 21554 507978
rect 21622 507922 21678 507978
rect 6970 496294 7026 496350
rect 7094 496294 7150 496350
rect 7218 496294 7274 496350
rect 7342 496294 7398 496350
rect 6970 496170 7026 496226
rect 7094 496170 7150 496226
rect 7218 496170 7274 496226
rect 7342 496170 7398 496226
rect 6970 496046 7026 496102
rect 7094 496046 7150 496102
rect 7218 496046 7274 496102
rect 7342 496046 7398 496102
rect 6970 495922 7026 495978
rect 7094 495922 7150 495978
rect 7218 495922 7274 495978
rect 7342 495922 7398 495978
rect 6970 478294 7026 478350
rect 7094 478294 7150 478350
rect 7218 478294 7274 478350
rect 7342 478294 7398 478350
rect 6970 478170 7026 478226
rect 7094 478170 7150 478226
rect 7218 478170 7274 478226
rect 7342 478170 7398 478226
rect 6970 478046 7026 478102
rect 7094 478046 7150 478102
rect 7218 478046 7274 478102
rect 7342 478046 7398 478102
rect 6970 477922 7026 477978
rect 7094 477922 7150 477978
rect 7218 477922 7274 477978
rect 7342 477922 7398 477978
rect 6970 460294 7026 460350
rect 7094 460294 7150 460350
rect 7218 460294 7274 460350
rect 7342 460294 7398 460350
rect 6970 460170 7026 460226
rect 7094 460170 7150 460226
rect 7218 460170 7274 460226
rect 7342 460170 7398 460226
rect 6970 460046 7026 460102
rect 7094 460046 7150 460102
rect 7218 460046 7274 460102
rect 7342 460046 7398 460102
rect 6970 459922 7026 459978
rect 7094 459922 7150 459978
rect 7218 459922 7274 459978
rect 7342 459922 7398 459978
rect 6970 442294 7026 442350
rect 7094 442294 7150 442350
rect 7218 442294 7274 442350
rect 7342 442294 7398 442350
rect 6970 442170 7026 442226
rect 7094 442170 7150 442226
rect 7218 442170 7274 442226
rect 7342 442170 7398 442226
rect 6970 442046 7026 442102
rect 7094 442046 7150 442102
rect 7218 442046 7274 442102
rect 7342 442046 7398 442102
rect 6970 441922 7026 441978
rect 7094 441922 7150 441978
rect 7218 441922 7274 441978
rect 7342 441922 7398 441978
rect 6970 424294 7026 424350
rect 7094 424294 7150 424350
rect 7218 424294 7274 424350
rect 7342 424294 7398 424350
rect 6970 424170 7026 424226
rect 7094 424170 7150 424226
rect 7218 424170 7274 424226
rect 7342 424170 7398 424226
rect 6970 424046 7026 424102
rect 7094 424046 7150 424102
rect 7218 424046 7274 424102
rect 7342 424046 7398 424102
rect 6970 423922 7026 423978
rect 7094 423922 7150 423978
rect 7218 423922 7274 423978
rect 7342 423922 7398 423978
rect 6970 406294 7026 406350
rect 7094 406294 7150 406350
rect 7218 406294 7274 406350
rect 7342 406294 7398 406350
rect 6970 406170 7026 406226
rect 7094 406170 7150 406226
rect 7218 406170 7274 406226
rect 7342 406170 7398 406226
rect 6970 406046 7026 406102
rect 7094 406046 7150 406102
rect 7218 406046 7274 406102
rect 7342 406046 7398 406102
rect 6970 405922 7026 405978
rect 7094 405922 7150 405978
rect 7218 405922 7274 405978
rect 7342 405922 7398 405978
rect 6970 388294 7026 388350
rect 7094 388294 7150 388350
rect 7218 388294 7274 388350
rect 7342 388294 7398 388350
rect 6970 388170 7026 388226
rect 7094 388170 7150 388226
rect 7218 388170 7274 388226
rect 7342 388170 7398 388226
rect 6970 388046 7026 388102
rect 7094 388046 7150 388102
rect 7218 388046 7274 388102
rect 7342 388046 7398 388102
rect 6970 387922 7026 387978
rect 7094 387922 7150 387978
rect 7218 387922 7274 387978
rect 7342 387922 7398 387978
rect 6970 370294 7026 370350
rect 7094 370294 7150 370350
rect 7218 370294 7274 370350
rect 7342 370294 7398 370350
rect 6970 370170 7026 370226
rect 7094 370170 7150 370226
rect 7218 370170 7274 370226
rect 7342 370170 7398 370226
rect 6970 370046 7026 370102
rect 7094 370046 7150 370102
rect 7218 370046 7274 370102
rect 7342 370046 7398 370102
rect 6970 369922 7026 369978
rect 7094 369922 7150 369978
rect 7218 369922 7274 369978
rect 7342 369922 7398 369978
rect 6970 352294 7026 352350
rect 7094 352294 7150 352350
rect 7218 352294 7274 352350
rect 7342 352294 7398 352350
rect 6970 352170 7026 352226
rect 7094 352170 7150 352226
rect 7218 352170 7274 352226
rect 7342 352170 7398 352226
rect 6970 352046 7026 352102
rect 7094 352046 7150 352102
rect 7218 352046 7274 352102
rect 7342 352046 7398 352102
rect 6970 351922 7026 351978
rect 7094 351922 7150 351978
rect 7218 351922 7274 351978
rect 7342 351922 7398 351978
rect 6970 334294 7026 334350
rect 7094 334294 7150 334350
rect 7218 334294 7274 334350
rect 7342 334294 7398 334350
rect 6970 334170 7026 334226
rect 7094 334170 7150 334226
rect 7218 334170 7274 334226
rect 7342 334170 7398 334226
rect 6970 334046 7026 334102
rect 7094 334046 7150 334102
rect 7218 334046 7274 334102
rect 7342 334046 7398 334102
rect 6970 333922 7026 333978
rect 7094 333922 7150 333978
rect 7218 333922 7274 333978
rect 7342 333922 7398 333978
rect 6970 316294 7026 316350
rect 7094 316294 7150 316350
rect 7218 316294 7274 316350
rect 7342 316294 7398 316350
rect 6970 316170 7026 316226
rect 7094 316170 7150 316226
rect 7218 316170 7274 316226
rect 7342 316170 7398 316226
rect 6970 316046 7026 316102
rect 7094 316046 7150 316102
rect 7218 316046 7274 316102
rect 7342 316046 7398 316102
rect 6970 315922 7026 315978
rect 7094 315922 7150 315978
rect 7218 315922 7274 315978
rect 7342 315922 7398 315978
rect 6970 298294 7026 298350
rect 7094 298294 7150 298350
rect 7218 298294 7274 298350
rect 7342 298294 7398 298350
rect 6970 298170 7026 298226
rect 7094 298170 7150 298226
rect 7218 298170 7274 298226
rect 7342 298170 7398 298226
rect 6970 298046 7026 298102
rect 7094 298046 7150 298102
rect 7218 298046 7274 298102
rect 7342 298046 7398 298102
rect 6970 297922 7026 297978
rect 7094 297922 7150 297978
rect 7218 297922 7274 297978
rect 7342 297922 7398 297978
rect 6970 280294 7026 280350
rect 7094 280294 7150 280350
rect 7218 280294 7274 280350
rect 7342 280294 7398 280350
rect 6970 280170 7026 280226
rect 7094 280170 7150 280226
rect 7218 280170 7274 280226
rect 7342 280170 7398 280226
rect 6970 280046 7026 280102
rect 7094 280046 7150 280102
rect 7218 280046 7274 280102
rect 7342 280046 7398 280102
rect 6970 279922 7026 279978
rect 7094 279922 7150 279978
rect 7218 279922 7274 279978
rect 7342 279922 7398 279978
rect 6970 262294 7026 262350
rect 7094 262294 7150 262350
rect 7218 262294 7274 262350
rect 7342 262294 7398 262350
rect 6970 262170 7026 262226
rect 7094 262170 7150 262226
rect 7218 262170 7274 262226
rect 7342 262170 7398 262226
rect 6970 262046 7026 262102
rect 7094 262046 7150 262102
rect 7218 262046 7274 262102
rect 7342 262046 7398 262102
rect 6970 261922 7026 261978
rect 7094 261922 7150 261978
rect 7218 261922 7274 261978
rect 7342 261922 7398 261978
rect 6970 244294 7026 244350
rect 7094 244294 7150 244350
rect 7218 244294 7274 244350
rect 7342 244294 7398 244350
rect 6970 244170 7026 244226
rect 7094 244170 7150 244226
rect 7218 244170 7274 244226
rect 7342 244170 7398 244226
rect 6970 244046 7026 244102
rect 7094 244046 7150 244102
rect 7218 244046 7274 244102
rect 7342 244046 7398 244102
rect 6970 243922 7026 243978
rect 7094 243922 7150 243978
rect 7218 243922 7274 243978
rect 7342 243922 7398 243978
rect 6970 226294 7026 226350
rect 7094 226294 7150 226350
rect 7218 226294 7274 226350
rect 7342 226294 7398 226350
rect 6970 226170 7026 226226
rect 7094 226170 7150 226226
rect 7218 226170 7274 226226
rect 7342 226170 7398 226226
rect 6970 226046 7026 226102
rect 7094 226046 7150 226102
rect 7218 226046 7274 226102
rect 7342 226046 7398 226102
rect 6970 225922 7026 225978
rect 7094 225922 7150 225978
rect 7218 225922 7274 225978
rect 7342 225922 7398 225978
rect 6970 208294 7026 208350
rect 7094 208294 7150 208350
rect 7218 208294 7274 208350
rect 7342 208294 7398 208350
rect 6970 208170 7026 208226
rect 7094 208170 7150 208226
rect 7218 208170 7274 208226
rect 7342 208170 7398 208226
rect 6970 208046 7026 208102
rect 7094 208046 7150 208102
rect 7218 208046 7274 208102
rect 7342 208046 7398 208102
rect 6970 207922 7026 207978
rect 7094 207922 7150 207978
rect 7218 207922 7274 207978
rect 7342 207922 7398 207978
rect 6970 190294 7026 190350
rect 7094 190294 7150 190350
rect 7218 190294 7274 190350
rect 7342 190294 7398 190350
rect 6970 190170 7026 190226
rect 7094 190170 7150 190226
rect 7218 190170 7274 190226
rect 7342 190170 7398 190226
rect 6970 190046 7026 190102
rect 7094 190046 7150 190102
rect 7218 190046 7274 190102
rect 7342 190046 7398 190102
rect 6970 189922 7026 189978
rect 7094 189922 7150 189978
rect 7218 189922 7274 189978
rect 7342 189922 7398 189978
rect 6970 172294 7026 172350
rect 7094 172294 7150 172350
rect 7218 172294 7274 172350
rect 7342 172294 7398 172350
rect 6970 172170 7026 172226
rect 7094 172170 7150 172226
rect 7218 172170 7274 172226
rect 7342 172170 7398 172226
rect 6970 172046 7026 172102
rect 7094 172046 7150 172102
rect 7218 172046 7274 172102
rect 7342 172046 7398 172102
rect 6970 171922 7026 171978
rect 7094 171922 7150 171978
rect 7218 171922 7274 171978
rect 7342 171922 7398 171978
rect 6970 154294 7026 154350
rect 7094 154294 7150 154350
rect 7218 154294 7274 154350
rect 7342 154294 7398 154350
rect 6970 154170 7026 154226
rect 7094 154170 7150 154226
rect 7218 154170 7274 154226
rect 7342 154170 7398 154226
rect 6970 154046 7026 154102
rect 7094 154046 7150 154102
rect 7218 154046 7274 154102
rect 7342 154046 7398 154102
rect 6970 153922 7026 153978
rect 7094 153922 7150 153978
rect 7218 153922 7274 153978
rect 7342 153922 7398 153978
rect 6970 136294 7026 136350
rect 7094 136294 7150 136350
rect 7218 136294 7274 136350
rect 7342 136294 7398 136350
rect 6970 136170 7026 136226
rect 7094 136170 7150 136226
rect 7218 136170 7274 136226
rect 7342 136170 7398 136226
rect 6970 136046 7026 136102
rect 7094 136046 7150 136102
rect 7218 136046 7274 136102
rect 7342 136046 7398 136102
rect 6970 135922 7026 135978
rect 7094 135922 7150 135978
rect 7218 135922 7274 135978
rect 7342 135922 7398 135978
rect 6970 118294 7026 118350
rect 7094 118294 7150 118350
rect 7218 118294 7274 118350
rect 7342 118294 7398 118350
rect 6970 118170 7026 118226
rect 7094 118170 7150 118226
rect 7218 118170 7274 118226
rect 7342 118170 7398 118226
rect 6970 118046 7026 118102
rect 7094 118046 7150 118102
rect 7218 118046 7274 118102
rect 7342 118046 7398 118102
rect 6970 117922 7026 117978
rect 7094 117922 7150 117978
rect 7218 117922 7274 117978
rect 7342 117922 7398 117978
rect 6970 100294 7026 100350
rect 7094 100294 7150 100350
rect 7218 100294 7274 100350
rect 7342 100294 7398 100350
rect 6970 100170 7026 100226
rect 7094 100170 7150 100226
rect 7218 100170 7274 100226
rect 7342 100170 7398 100226
rect 6970 100046 7026 100102
rect 7094 100046 7150 100102
rect 7218 100046 7274 100102
rect 7342 100046 7398 100102
rect 6970 99922 7026 99978
rect 7094 99922 7150 99978
rect 7218 99922 7274 99978
rect 7342 99922 7398 99978
rect 6970 82294 7026 82350
rect 7094 82294 7150 82350
rect 7218 82294 7274 82350
rect 7342 82294 7398 82350
rect 6970 82170 7026 82226
rect 7094 82170 7150 82226
rect 7218 82170 7274 82226
rect 7342 82170 7398 82226
rect 6970 82046 7026 82102
rect 7094 82046 7150 82102
rect 7218 82046 7274 82102
rect 7342 82046 7398 82102
rect 6970 81922 7026 81978
rect 7094 81922 7150 81978
rect 7218 81922 7274 81978
rect 7342 81922 7398 81978
rect 21250 490294 21306 490350
rect 21374 490294 21430 490350
rect 21498 490294 21554 490350
rect 21622 490294 21678 490350
rect 21250 490170 21306 490226
rect 21374 490170 21430 490226
rect 21498 490170 21554 490226
rect 21622 490170 21678 490226
rect 21250 490046 21306 490102
rect 21374 490046 21430 490102
rect 21498 490046 21554 490102
rect 21622 490046 21678 490102
rect 21250 489922 21306 489978
rect 21374 489922 21430 489978
rect 21498 489922 21554 489978
rect 21622 489922 21678 489978
rect 21250 472294 21306 472350
rect 21374 472294 21430 472350
rect 21498 472294 21554 472350
rect 21622 472294 21678 472350
rect 21250 472170 21306 472226
rect 21374 472170 21430 472226
rect 21498 472170 21554 472226
rect 21622 472170 21678 472226
rect 21250 472046 21306 472102
rect 21374 472046 21430 472102
rect 21498 472046 21554 472102
rect 21622 472046 21678 472102
rect 21250 471922 21306 471978
rect 21374 471922 21430 471978
rect 21498 471922 21554 471978
rect 21622 471922 21678 471978
rect 21250 454294 21306 454350
rect 21374 454294 21430 454350
rect 21498 454294 21554 454350
rect 21622 454294 21678 454350
rect 21250 454170 21306 454226
rect 21374 454170 21430 454226
rect 21498 454170 21554 454226
rect 21622 454170 21678 454226
rect 21250 454046 21306 454102
rect 21374 454046 21430 454102
rect 21498 454046 21554 454102
rect 21622 454046 21678 454102
rect 21250 453922 21306 453978
rect 21374 453922 21430 453978
rect 21498 453922 21554 453978
rect 21622 453922 21678 453978
rect 21250 436294 21306 436350
rect 21374 436294 21430 436350
rect 21498 436294 21554 436350
rect 21622 436294 21678 436350
rect 21250 436170 21306 436226
rect 21374 436170 21430 436226
rect 21498 436170 21554 436226
rect 21622 436170 21678 436226
rect 21250 436046 21306 436102
rect 21374 436046 21430 436102
rect 21498 436046 21554 436102
rect 21622 436046 21678 436102
rect 21250 435922 21306 435978
rect 21374 435922 21430 435978
rect 21498 435922 21554 435978
rect 21622 435922 21678 435978
rect 21250 418294 21306 418350
rect 21374 418294 21430 418350
rect 21498 418294 21554 418350
rect 21622 418294 21678 418350
rect 21250 418170 21306 418226
rect 21374 418170 21430 418226
rect 21498 418170 21554 418226
rect 21622 418170 21678 418226
rect 21250 418046 21306 418102
rect 21374 418046 21430 418102
rect 21498 418046 21554 418102
rect 21622 418046 21678 418102
rect 21250 417922 21306 417978
rect 21374 417922 21430 417978
rect 21498 417922 21554 417978
rect 21622 417922 21678 417978
rect 21250 400294 21306 400350
rect 21374 400294 21430 400350
rect 21498 400294 21554 400350
rect 21622 400294 21678 400350
rect 21250 400170 21306 400226
rect 21374 400170 21430 400226
rect 21498 400170 21554 400226
rect 21622 400170 21678 400226
rect 21250 400046 21306 400102
rect 21374 400046 21430 400102
rect 21498 400046 21554 400102
rect 21622 400046 21678 400102
rect 21250 399922 21306 399978
rect 21374 399922 21430 399978
rect 21498 399922 21554 399978
rect 21622 399922 21678 399978
rect 21250 382294 21306 382350
rect 21374 382294 21430 382350
rect 21498 382294 21554 382350
rect 21622 382294 21678 382350
rect 21250 382170 21306 382226
rect 21374 382170 21430 382226
rect 21498 382170 21554 382226
rect 21622 382170 21678 382226
rect 21250 382046 21306 382102
rect 21374 382046 21430 382102
rect 21498 382046 21554 382102
rect 21622 382046 21678 382102
rect 21250 381922 21306 381978
rect 21374 381922 21430 381978
rect 21498 381922 21554 381978
rect 21622 381922 21678 381978
rect 21250 364294 21306 364350
rect 21374 364294 21430 364350
rect 21498 364294 21554 364350
rect 21622 364294 21678 364350
rect 21250 364170 21306 364226
rect 21374 364170 21430 364226
rect 21498 364170 21554 364226
rect 21622 364170 21678 364226
rect 21250 364046 21306 364102
rect 21374 364046 21430 364102
rect 21498 364046 21554 364102
rect 21622 364046 21678 364102
rect 21250 363922 21306 363978
rect 21374 363922 21430 363978
rect 21498 363922 21554 363978
rect 21622 363922 21678 363978
rect 21250 346294 21306 346350
rect 21374 346294 21430 346350
rect 21498 346294 21554 346350
rect 21622 346294 21678 346350
rect 21250 346170 21306 346226
rect 21374 346170 21430 346226
rect 21498 346170 21554 346226
rect 21622 346170 21678 346226
rect 21250 346046 21306 346102
rect 21374 346046 21430 346102
rect 21498 346046 21554 346102
rect 21622 346046 21678 346102
rect 21250 345922 21306 345978
rect 21374 345922 21430 345978
rect 21498 345922 21554 345978
rect 21622 345922 21678 345978
rect 21250 328294 21306 328350
rect 21374 328294 21430 328350
rect 21498 328294 21554 328350
rect 21622 328294 21678 328350
rect 21250 328170 21306 328226
rect 21374 328170 21430 328226
rect 21498 328170 21554 328226
rect 21622 328170 21678 328226
rect 21250 328046 21306 328102
rect 21374 328046 21430 328102
rect 21498 328046 21554 328102
rect 21622 328046 21678 328102
rect 21250 327922 21306 327978
rect 21374 327922 21430 327978
rect 21498 327922 21554 327978
rect 21622 327922 21678 327978
rect 21250 310294 21306 310350
rect 21374 310294 21430 310350
rect 21498 310294 21554 310350
rect 21622 310294 21678 310350
rect 21250 310170 21306 310226
rect 21374 310170 21430 310226
rect 21498 310170 21554 310226
rect 21622 310170 21678 310226
rect 21250 310046 21306 310102
rect 21374 310046 21430 310102
rect 21498 310046 21554 310102
rect 21622 310046 21678 310102
rect 21250 309922 21306 309978
rect 21374 309922 21430 309978
rect 21498 309922 21554 309978
rect 21622 309922 21678 309978
rect 21250 292294 21306 292350
rect 21374 292294 21430 292350
rect 21498 292294 21554 292350
rect 21622 292294 21678 292350
rect 21250 292170 21306 292226
rect 21374 292170 21430 292226
rect 21498 292170 21554 292226
rect 21622 292170 21678 292226
rect 21250 292046 21306 292102
rect 21374 292046 21430 292102
rect 21498 292046 21554 292102
rect 21622 292046 21678 292102
rect 21250 291922 21306 291978
rect 21374 291922 21430 291978
rect 21498 291922 21554 291978
rect 21622 291922 21678 291978
rect 21250 274294 21306 274350
rect 21374 274294 21430 274350
rect 21498 274294 21554 274350
rect 21622 274294 21678 274350
rect 21250 274170 21306 274226
rect 21374 274170 21430 274226
rect 21498 274170 21554 274226
rect 21622 274170 21678 274226
rect 21250 274046 21306 274102
rect 21374 274046 21430 274102
rect 21498 274046 21554 274102
rect 21622 274046 21678 274102
rect 21250 273922 21306 273978
rect 21374 273922 21430 273978
rect 21498 273922 21554 273978
rect 21622 273922 21678 273978
rect 21250 256294 21306 256350
rect 21374 256294 21430 256350
rect 21498 256294 21554 256350
rect 21622 256294 21678 256350
rect 21250 256170 21306 256226
rect 21374 256170 21430 256226
rect 21498 256170 21554 256226
rect 21622 256170 21678 256226
rect 21250 256046 21306 256102
rect 21374 256046 21430 256102
rect 21498 256046 21554 256102
rect 21622 256046 21678 256102
rect 21250 255922 21306 255978
rect 21374 255922 21430 255978
rect 21498 255922 21554 255978
rect 21622 255922 21678 255978
rect 21250 238294 21306 238350
rect 21374 238294 21430 238350
rect 21498 238294 21554 238350
rect 21622 238294 21678 238350
rect 21250 238170 21306 238226
rect 21374 238170 21430 238226
rect 21498 238170 21554 238226
rect 21622 238170 21678 238226
rect 21250 238046 21306 238102
rect 21374 238046 21430 238102
rect 21498 238046 21554 238102
rect 21622 238046 21678 238102
rect 21250 237922 21306 237978
rect 21374 237922 21430 237978
rect 21498 237922 21554 237978
rect 21622 237922 21678 237978
rect 21250 220294 21306 220350
rect 21374 220294 21430 220350
rect 21498 220294 21554 220350
rect 21622 220294 21678 220350
rect 21250 220170 21306 220226
rect 21374 220170 21430 220226
rect 21498 220170 21554 220226
rect 21622 220170 21678 220226
rect 21250 220046 21306 220102
rect 21374 220046 21430 220102
rect 21498 220046 21554 220102
rect 21622 220046 21678 220102
rect 21250 219922 21306 219978
rect 21374 219922 21430 219978
rect 21498 219922 21554 219978
rect 21622 219922 21678 219978
rect 21250 202294 21306 202350
rect 21374 202294 21430 202350
rect 21498 202294 21554 202350
rect 21622 202294 21678 202350
rect 21250 202170 21306 202226
rect 21374 202170 21430 202226
rect 21498 202170 21554 202226
rect 21622 202170 21678 202226
rect 21250 202046 21306 202102
rect 21374 202046 21430 202102
rect 21498 202046 21554 202102
rect 21622 202046 21678 202102
rect 21250 201922 21306 201978
rect 21374 201922 21430 201978
rect 21498 201922 21554 201978
rect 21622 201922 21678 201978
rect 21250 184294 21306 184350
rect 21374 184294 21430 184350
rect 21498 184294 21554 184350
rect 21622 184294 21678 184350
rect 21250 184170 21306 184226
rect 21374 184170 21430 184226
rect 21498 184170 21554 184226
rect 21622 184170 21678 184226
rect 21250 184046 21306 184102
rect 21374 184046 21430 184102
rect 21498 184046 21554 184102
rect 21622 184046 21678 184102
rect 21250 183922 21306 183978
rect 21374 183922 21430 183978
rect 21498 183922 21554 183978
rect 21622 183922 21678 183978
rect 24970 514294 25026 514350
rect 25094 514294 25150 514350
rect 25218 514294 25274 514350
rect 25342 514294 25398 514350
rect 24970 514170 25026 514226
rect 25094 514170 25150 514226
rect 25218 514170 25274 514226
rect 25342 514170 25398 514226
rect 24970 514046 25026 514102
rect 25094 514046 25150 514102
rect 25218 514046 25274 514102
rect 25342 514046 25398 514102
rect 24970 513922 25026 513978
rect 25094 513922 25150 513978
rect 25218 513922 25274 513978
rect 25342 513922 25398 513978
rect 24970 496294 25026 496350
rect 25094 496294 25150 496350
rect 25218 496294 25274 496350
rect 25342 496294 25398 496350
rect 24970 496170 25026 496226
rect 25094 496170 25150 496226
rect 25218 496170 25274 496226
rect 25342 496170 25398 496226
rect 24970 496046 25026 496102
rect 25094 496046 25150 496102
rect 25218 496046 25274 496102
rect 25342 496046 25398 496102
rect 24970 495922 25026 495978
rect 25094 495922 25150 495978
rect 25218 495922 25274 495978
rect 25342 495922 25398 495978
rect 24970 478294 25026 478350
rect 25094 478294 25150 478350
rect 25218 478294 25274 478350
rect 25342 478294 25398 478350
rect 24970 478170 25026 478226
rect 25094 478170 25150 478226
rect 25218 478170 25274 478226
rect 25342 478170 25398 478226
rect 24970 478046 25026 478102
rect 25094 478046 25150 478102
rect 25218 478046 25274 478102
rect 25342 478046 25398 478102
rect 24970 477922 25026 477978
rect 25094 477922 25150 477978
rect 25218 477922 25274 477978
rect 25342 477922 25398 477978
rect 24970 460294 25026 460350
rect 25094 460294 25150 460350
rect 25218 460294 25274 460350
rect 25342 460294 25398 460350
rect 24970 460170 25026 460226
rect 25094 460170 25150 460226
rect 25218 460170 25274 460226
rect 25342 460170 25398 460226
rect 24970 460046 25026 460102
rect 25094 460046 25150 460102
rect 25218 460046 25274 460102
rect 25342 460046 25398 460102
rect 24970 459922 25026 459978
rect 25094 459922 25150 459978
rect 25218 459922 25274 459978
rect 25342 459922 25398 459978
rect 24970 442294 25026 442350
rect 25094 442294 25150 442350
rect 25218 442294 25274 442350
rect 25342 442294 25398 442350
rect 24970 442170 25026 442226
rect 25094 442170 25150 442226
rect 25218 442170 25274 442226
rect 25342 442170 25398 442226
rect 24970 442046 25026 442102
rect 25094 442046 25150 442102
rect 25218 442046 25274 442102
rect 25342 442046 25398 442102
rect 24970 441922 25026 441978
rect 25094 441922 25150 441978
rect 25218 441922 25274 441978
rect 25342 441922 25398 441978
rect 24970 424294 25026 424350
rect 25094 424294 25150 424350
rect 25218 424294 25274 424350
rect 25342 424294 25398 424350
rect 24970 424170 25026 424226
rect 25094 424170 25150 424226
rect 25218 424170 25274 424226
rect 25342 424170 25398 424226
rect 24970 424046 25026 424102
rect 25094 424046 25150 424102
rect 25218 424046 25274 424102
rect 25342 424046 25398 424102
rect 24970 423922 25026 423978
rect 25094 423922 25150 423978
rect 25218 423922 25274 423978
rect 25342 423922 25398 423978
rect 24970 406294 25026 406350
rect 25094 406294 25150 406350
rect 25218 406294 25274 406350
rect 25342 406294 25398 406350
rect 24970 406170 25026 406226
rect 25094 406170 25150 406226
rect 25218 406170 25274 406226
rect 25342 406170 25398 406226
rect 24970 406046 25026 406102
rect 25094 406046 25150 406102
rect 25218 406046 25274 406102
rect 25342 406046 25398 406102
rect 24970 405922 25026 405978
rect 25094 405922 25150 405978
rect 25218 405922 25274 405978
rect 25342 405922 25398 405978
rect 24970 388294 25026 388350
rect 25094 388294 25150 388350
rect 25218 388294 25274 388350
rect 25342 388294 25398 388350
rect 24970 388170 25026 388226
rect 25094 388170 25150 388226
rect 25218 388170 25274 388226
rect 25342 388170 25398 388226
rect 24970 388046 25026 388102
rect 25094 388046 25150 388102
rect 25218 388046 25274 388102
rect 25342 388046 25398 388102
rect 24970 387922 25026 387978
rect 25094 387922 25150 387978
rect 25218 387922 25274 387978
rect 25342 387922 25398 387978
rect 24970 370294 25026 370350
rect 25094 370294 25150 370350
rect 25218 370294 25274 370350
rect 25342 370294 25398 370350
rect 24970 370170 25026 370226
rect 25094 370170 25150 370226
rect 25218 370170 25274 370226
rect 25342 370170 25398 370226
rect 24970 370046 25026 370102
rect 25094 370046 25150 370102
rect 25218 370046 25274 370102
rect 25342 370046 25398 370102
rect 24970 369922 25026 369978
rect 25094 369922 25150 369978
rect 25218 369922 25274 369978
rect 25342 369922 25398 369978
rect 24970 352294 25026 352350
rect 25094 352294 25150 352350
rect 25218 352294 25274 352350
rect 25342 352294 25398 352350
rect 24970 352170 25026 352226
rect 25094 352170 25150 352226
rect 25218 352170 25274 352226
rect 25342 352170 25398 352226
rect 24970 352046 25026 352102
rect 25094 352046 25150 352102
rect 25218 352046 25274 352102
rect 25342 352046 25398 352102
rect 24970 351922 25026 351978
rect 25094 351922 25150 351978
rect 25218 351922 25274 351978
rect 25342 351922 25398 351978
rect 24970 334294 25026 334350
rect 25094 334294 25150 334350
rect 25218 334294 25274 334350
rect 25342 334294 25398 334350
rect 24970 334170 25026 334226
rect 25094 334170 25150 334226
rect 25218 334170 25274 334226
rect 25342 334170 25398 334226
rect 24970 334046 25026 334102
rect 25094 334046 25150 334102
rect 25218 334046 25274 334102
rect 25342 334046 25398 334102
rect 24970 333922 25026 333978
rect 25094 333922 25150 333978
rect 25218 333922 25274 333978
rect 25342 333922 25398 333978
rect 24970 316294 25026 316350
rect 25094 316294 25150 316350
rect 25218 316294 25274 316350
rect 25342 316294 25398 316350
rect 24970 316170 25026 316226
rect 25094 316170 25150 316226
rect 25218 316170 25274 316226
rect 25342 316170 25398 316226
rect 24970 316046 25026 316102
rect 25094 316046 25150 316102
rect 25218 316046 25274 316102
rect 25342 316046 25398 316102
rect 24970 315922 25026 315978
rect 25094 315922 25150 315978
rect 25218 315922 25274 315978
rect 25342 315922 25398 315978
rect 24970 298294 25026 298350
rect 25094 298294 25150 298350
rect 25218 298294 25274 298350
rect 25342 298294 25398 298350
rect 24970 298170 25026 298226
rect 25094 298170 25150 298226
rect 25218 298170 25274 298226
rect 25342 298170 25398 298226
rect 24970 298046 25026 298102
rect 25094 298046 25150 298102
rect 25218 298046 25274 298102
rect 25342 298046 25398 298102
rect 24970 297922 25026 297978
rect 25094 297922 25150 297978
rect 25218 297922 25274 297978
rect 25342 297922 25398 297978
rect 21250 166294 21306 166350
rect 21374 166294 21430 166350
rect 21498 166294 21554 166350
rect 21622 166294 21678 166350
rect 21250 166170 21306 166226
rect 21374 166170 21430 166226
rect 21498 166170 21554 166226
rect 21622 166170 21678 166226
rect 21250 166046 21306 166102
rect 21374 166046 21430 166102
rect 21498 166046 21554 166102
rect 21622 166046 21678 166102
rect 21250 165922 21306 165978
rect 21374 165922 21430 165978
rect 21498 165922 21554 165978
rect 21622 165922 21678 165978
rect 21250 148294 21306 148350
rect 21374 148294 21430 148350
rect 21498 148294 21554 148350
rect 21622 148294 21678 148350
rect 21250 148170 21306 148226
rect 21374 148170 21430 148226
rect 21498 148170 21554 148226
rect 21622 148170 21678 148226
rect 21250 148046 21306 148102
rect 21374 148046 21430 148102
rect 21498 148046 21554 148102
rect 21622 148046 21678 148102
rect 21250 147922 21306 147978
rect 21374 147922 21430 147978
rect 21498 147922 21554 147978
rect 21622 147922 21678 147978
rect 21250 130294 21306 130350
rect 21374 130294 21430 130350
rect 21498 130294 21554 130350
rect 21622 130294 21678 130350
rect 21250 130170 21306 130226
rect 21374 130170 21430 130226
rect 21498 130170 21554 130226
rect 21622 130170 21678 130226
rect 21250 130046 21306 130102
rect 21374 130046 21430 130102
rect 21498 130046 21554 130102
rect 21622 130046 21678 130102
rect 21250 129922 21306 129978
rect 21374 129922 21430 129978
rect 21498 129922 21554 129978
rect 21622 129922 21678 129978
rect 24970 280294 25026 280350
rect 25094 280294 25150 280350
rect 25218 280294 25274 280350
rect 25342 280294 25398 280350
rect 24970 280170 25026 280226
rect 25094 280170 25150 280226
rect 25218 280170 25274 280226
rect 25342 280170 25398 280226
rect 24970 280046 25026 280102
rect 25094 280046 25150 280102
rect 25218 280046 25274 280102
rect 25342 280046 25398 280102
rect 24970 279922 25026 279978
rect 25094 279922 25150 279978
rect 25218 279922 25274 279978
rect 25342 279922 25398 279978
rect 24970 262294 25026 262350
rect 25094 262294 25150 262350
rect 25218 262294 25274 262350
rect 25342 262294 25398 262350
rect 24970 262170 25026 262226
rect 25094 262170 25150 262226
rect 25218 262170 25274 262226
rect 25342 262170 25398 262226
rect 24970 262046 25026 262102
rect 25094 262046 25150 262102
rect 25218 262046 25274 262102
rect 25342 262046 25398 262102
rect 24970 261922 25026 261978
rect 25094 261922 25150 261978
rect 25218 261922 25274 261978
rect 25342 261922 25398 261978
rect 24970 244294 25026 244350
rect 25094 244294 25150 244350
rect 25218 244294 25274 244350
rect 25342 244294 25398 244350
rect 24970 244170 25026 244226
rect 25094 244170 25150 244226
rect 25218 244170 25274 244226
rect 25342 244170 25398 244226
rect 24970 244046 25026 244102
rect 25094 244046 25150 244102
rect 25218 244046 25274 244102
rect 25342 244046 25398 244102
rect 24970 243922 25026 243978
rect 25094 243922 25150 243978
rect 25218 243922 25274 243978
rect 25342 243922 25398 243978
rect 24970 226294 25026 226350
rect 25094 226294 25150 226350
rect 25218 226294 25274 226350
rect 25342 226294 25398 226350
rect 24970 226170 25026 226226
rect 25094 226170 25150 226226
rect 25218 226170 25274 226226
rect 25342 226170 25398 226226
rect 24970 226046 25026 226102
rect 25094 226046 25150 226102
rect 25218 226046 25274 226102
rect 25342 226046 25398 226102
rect 24970 225922 25026 225978
rect 25094 225922 25150 225978
rect 25218 225922 25274 225978
rect 25342 225922 25398 225978
rect 24970 208294 25026 208350
rect 25094 208294 25150 208350
rect 25218 208294 25274 208350
rect 25342 208294 25398 208350
rect 24970 208170 25026 208226
rect 25094 208170 25150 208226
rect 25218 208170 25274 208226
rect 25342 208170 25398 208226
rect 24970 208046 25026 208102
rect 25094 208046 25150 208102
rect 25218 208046 25274 208102
rect 25342 208046 25398 208102
rect 24970 207922 25026 207978
rect 25094 207922 25150 207978
rect 25218 207922 25274 207978
rect 25342 207922 25398 207978
rect 24970 190294 25026 190350
rect 25094 190294 25150 190350
rect 25218 190294 25274 190350
rect 25342 190294 25398 190350
rect 24970 190170 25026 190226
rect 25094 190170 25150 190226
rect 25218 190170 25274 190226
rect 25342 190170 25398 190226
rect 24970 190046 25026 190102
rect 25094 190046 25150 190102
rect 25218 190046 25274 190102
rect 25342 190046 25398 190102
rect 24970 189922 25026 189978
rect 25094 189922 25150 189978
rect 25218 189922 25274 189978
rect 25342 189922 25398 189978
rect 24970 172294 25026 172350
rect 25094 172294 25150 172350
rect 25218 172294 25274 172350
rect 25342 172294 25398 172350
rect 24970 172170 25026 172226
rect 25094 172170 25150 172226
rect 25218 172170 25274 172226
rect 25342 172170 25398 172226
rect 24970 172046 25026 172102
rect 25094 172046 25150 172102
rect 25218 172046 25274 172102
rect 25342 172046 25398 172102
rect 24970 171922 25026 171978
rect 25094 171922 25150 171978
rect 25218 171922 25274 171978
rect 25342 171922 25398 171978
rect 24970 154294 25026 154350
rect 25094 154294 25150 154350
rect 25218 154294 25274 154350
rect 25342 154294 25398 154350
rect 24970 154170 25026 154226
rect 25094 154170 25150 154226
rect 25218 154170 25274 154226
rect 25342 154170 25398 154226
rect 24970 154046 25026 154102
rect 25094 154046 25150 154102
rect 25218 154046 25274 154102
rect 25342 154046 25398 154102
rect 24970 153922 25026 153978
rect 25094 153922 25150 153978
rect 25218 153922 25274 153978
rect 25342 153922 25398 153978
rect 24970 136294 25026 136350
rect 25094 136294 25150 136350
rect 25218 136294 25274 136350
rect 25342 136294 25398 136350
rect 24970 136170 25026 136226
rect 25094 136170 25150 136226
rect 25218 136170 25274 136226
rect 25342 136170 25398 136226
rect 24970 136046 25026 136102
rect 25094 136046 25150 136102
rect 25218 136046 25274 136102
rect 25342 136046 25398 136102
rect 24970 135922 25026 135978
rect 25094 135922 25150 135978
rect 25218 135922 25274 135978
rect 25342 135922 25398 135978
rect 24970 118294 25026 118350
rect 25094 118294 25150 118350
rect 25218 118294 25274 118350
rect 25342 118294 25398 118350
rect 24970 118170 25026 118226
rect 25094 118170 25150 118226
rect 25218 118170 25274 118226
rect 25342 118170 25398 118226
rect 24970 118046 25026 118102
rect 25094 118046 25150 118102
rect 25218 118046 25274 118102
rect 25342 118046 25398 118102
rect 24970 117922 25026 117978
rect 25094 117922 25150 117978
rect 25218 117922 25274 117978
rect 25342 117922 25398 117978
rect 21250 112294 21306 112350
rect 21374 112294 21430 112350
rect 21498 112294 21554 112350
rect 21622 112294 21678 112350
rect 21250 112170 21306 112226
rect 21374 112170 21430 112226
rect 21498 112170 21554 112226
rect 21622 112170 21678 112226
rect 21250 112046 21306 112102
rect 21374 112046 21430 112102
rect 21498 112046 21554 112102
rect 21622 112046 21678 112102
rect 21250 111922 21306 111978
rect 21374 111922 21430 111978
rect 21498 111922 21554 111978
rect 21622 111922 21678 111978
rect 21250 94294 21306 94350
rect 21374 94294 21430 94350
rect 21498 94294 21554 94350
rect 21622 94294 21678 94350
rect 21250 94170 21306 94226
rect 21374 94170 21430 94226
rect 21498 94170 21554 94226
rect 21622 94170 21678 94226
rect 21250 94046 21306 94102
rect 21374 94046 21430 94102
rect 21498 94046 21554 94102
rect 21622 94046 21678 94102
rect 21250 93922 21306 93978
rect 21374 93922 21430 93978
rect 21498 93922 21554 93978
rect 21622 93922 21678 93978
rect 21250 76294 21306 76350
rect 21374 76294 21430 76350
rect 21498 76294 21554 76350
rect 21622 76294 21678 76350
rect 21250 76170 21306 76226
rect 21374 76170 21430 76226
rect 21498 76170 21554 76226
rect 21622 76170 21678 76226
rect 21250 76046 21306 76102
rect 21374 76046 21430 76102
rect 21498 76046 21554 76102
rect 21622 76046 21678 76102
rect 21250 75922 21306 75978
rect 21374 75922 21430 75978
rect 21498 75922 21554 75978
rect 21622 75922 21678 75978
rect 6970 64294 7026 64350
rect 7094 64294 7150 64350
rect 7218 64294 7274 64350
rect 7342 64294 7398 64350
rect 6970 64170 7026 64226
rect 7094 64170 7150 64226
rect 7218 64170 7274 64226
rect 7342 64170 7398 64226
rect 6970 64046 7026 64102
rect 7094 64046 7150 64102
rect 7218 64046 7274 64102
rect 7342 64046 7398 64102
rect 6970 63922 7026 63978
rect 7094 63922 7150 63978
rect 7218 63922 7274 63978
rect 7342 63922 7398 63978
rect 6970 46294 7026 46350
rect 7094 46294 7150 46350
rect 7218 46294 7274 46350
rect 7342 46294 7398 46350
rect 6970 46170 7026 46226
rect 7094 46170 7150 46226
rect 7218 46170 7274 46226
rect 7342 46170 7398 46226
rect 6970 46046 7026 46102
rect 7094 46046 7150 46102
rect 7218 46046 7274 46102
rect 7342 46046 7398 46102
rect 6970 45922 7026 45978
rect 7094 45922 7150 45978
rect 7218 45922 7274 45978
rect 7342 45922 7398 45978
rect 3250 40294 3306 40350
rect 3374 40294 3430 40350
rect 3498 40294 3554 40350
rect 3622 40294 3678 40350
rect 3250 40170 3306 40226
rect 3374 40170 3430 40226
rect 3498 40170 3554 40226
rect 3622 40170 3678 40226
rect 3250 40046 3306 40102
rect 3374 40046 3430 40102
rect 3498 40046 3554 40102
rect 3622 40046 3678 40102
rect 3250 39922 3306 39978
rect 3374 39922 3430 39978
rect 3498 39922 3554 39978
rect 3622 39922 3678 39978
rect 3250 22294 3306 22350
rect 3374 22294 3430 22350
rect 3498 22294 3554 22350
rect 3622 22294 3678 22350
rect 3250 22170 3306 22226
rect 3374 22170 3430 22226
rect 3498 22170 3554 22226
rect 3622 22170 3678 22226
rect 3250 22046 3306 22102
rect 3374 22046 3430 22102
rect 3498 22046 3554 22102
rect 3622 22046 3678 22102
rect 3250 21922 3306 21978
rect 3374 21922 3430 21978
rect 3498 21922 3554 21978
rect 3622 21922 3678 21978
rect 6970 28294 7026 28350
rect 7094 28294 7150 28350
rect 7218 28294 7274 28350
rect 7342 28294 7398 28350
rect 6970 28170 7026 28226
rect 7094 28170 7150 28226
rect 7218 28170 7274 28226
rect 7342 28170 7398 28226
rect 6970 28046 7026 28102
rect 7094 28046 7150 28102
rect 7218 28046 7274 28102
rect 7342 28046 7398 28102
rect 6970 27922 7026 27978
rect 7094 27922 7150 27978
rect 7218 27922 7274 27978
rect 7342 27922 7398 27978
rect 6970 10294 7026 10350
rect 7094 10294 7150 10350
rect 7218 10294 7274 10350
rect 7342 10294 7398 10350
rect 6970 10170 7026 10226
rect 7094 10170 7150 10226
rect 7218 10170 7274 10226
rect 7342 10170 7398 10226
rect 6970 10046 7026 10102
rect 7094 10046 7150 10102
rect 7218 10046 7274 10102
rect 7342 10046 7398 10102
rect 6970 9922 7026 9978
rect 7094 9922 7150 9978
rect 7218 9922 7274 9978
rect 7342 9922 7398 9978
rect 3250 4294 3306 4350
rect 3374 4294 3430 4350
rect 3498 4294 3554 4350
rect 3622 4294 3678 4350
rect 3250 4170 3306 4226
rect 3374 4170 3430 4226
rect 3498 4170 3554 4226
rect 3622 4170 3678 4226
rect 3250 4046 3306 4102
rect 3374 4046 3430 4102
rect 3498 4046 3554 4102
rect 3622 4046 3678 4102
rect 3250 3922 3306 3978
rect 3374 3922 3430 3978
rect 3498 3922 3554 3978
rect 3622 3922 3678 3978
rect 3250 -216 3306 -160
rect 3374 -216 3430 -160
rect 3498 -216 3554 -160
rect 3622 -216 3678 -160
rect 3250 -340 3306 -284
rect 3374 -340 3430 -284
rect 3498 -340 3554 -284
rect 3622 -340 3678 -284
rect 3250 -464 3306 -408
rect 3374 -464 3430 -408
rect 3498 -464 3554 -408
rect 3622 -464 3678 -408
rect 3250 -588 3306 -532
rect 3374 -588 3430 -532
rect 3498 -588 3554 -532
rect 3622 -588 3678 -532
rect -1820 -1176 -1764 -1120
rect -1696 -1176 -1640 -1120
rect -1572 -1176 -1516 -1120
rect -1448 -1176 -1392 -1120
rect -1820 -1300 -1764 -1244
rect -1696 -1300 -1640 -1244
rect -1572 -1300 -1516 -1244
rect -1448 -1300 -1392 -1244
rect -1820 -1424 -1764 -1368
rect -1696 -1424 -1640 -1368
rect -1572 -1424 -1516 -1368
rect -1448 -1424 -1392 -1368
rect -1820 -1548 -1764 -1492
rect -1696 -1548 -1640 -1492
rect -1572 -1548 -1516 -1492
rect -1448 -1548 -1392 -1492
rect 6970 -1176 7026 -1120
rect 7094 -1176 7150 -1120
rect 7218 -1176 7274 -1120
rect 7342 -1176 7398 -1120
rect 6970 -1300 7026 -1244
rect 7094 -1300 7150 -1244
rect 7218 -1300 7274 -1244
rect 7342 -1300 7398 -1244
rect 6970 -1424 7026 -1368
rect 7094 -1424 7150 -1368
rect 7218 -1424 7274 -1368
rect 7342 -1424 7398 -1368
rect 6970 -1548 7026 -1492
rect 7094 -1548 7150 -1492
rect 7218 -1548 7274 -1492
rect 7342 -1548 7398 -1492
rect 21250 58294 21306 58350
rect 21374 58294 21430 58350
rect 21498 58294 21554 58350
rect 21622 58294 21678 58350
rect 21250 58170 21306 58226
rect 21374 58170 21430 58226
rect 21498 58170 21554 58226
rect 21622 58170 21678 58226
rect 21250 58046 21306 58102
rect 21374 58046 21430 58102
rect 21498 58046 21554 58102
rect 21622 58046 21678 58102
rect 21250 57922 21306 57978
rect 21374 57922 21430 57978
rect 21498 57922 21554 57978
rect 21622 57922 21678 57978
rect 21250 40294 21306 40350
rect 21374 40294 21430 40350
rect 21498 40294 21554 40350
rect 21622 40294 21678 40350
rect 21250 40170 21306 40226
rect 21374 40170 21430 40226
rect 21498 40170 21554 40226
rect 21622 40170 21678 40226
rect 21250 40046 21306 40102
rect 21374 40046 21430 40102
rect 21498 40046 21554 40102
rect 21622 40046 21678 40102
rect 21250 39922 21306 39978
rect 21374 39922 21430 39978
rect 21498 39922 21554 39978
rect 21622 39922 21678 39978
rect 21250 22294 21306 22350
rect 21374 22294 21430 22350
rect 21498 22294 21554 22350
rect 21622 22294 21678 22350
rect 21250 22170 21306 22226
rect 21374 22170 21430 22226
rect 21498 22170 21554 22226
rect 21622 22170 21678 22226
rect 21250 22046 21306 22102
rect 21374 22046 21430 22102
rect 21498 22046 21554 22102
rect 21622 22046 21678 22102
rect 21250 21922 21306 21978
rect 21374 21922 21430 21978
rect 21498 21922 21554 21978
rect 21622 21922 21678 21978
rect 21250 4294 21306 4350
rect 21374 4294 21430 4350
rect 21498 4294 21554 4350
rect 21622 4294 21678 4350
rect 21250 4170 21306 4226
rect 21374 4170 21430 4226
rect 21498 4170 21554 4226
rect 21622 4170 21678 4226
rect 21250 4046 21306 4102
rect 21374 4046 21430 4102
rect 21498 4046 21554 4102
rect 21622 4046 21678 4102
rect 21250 3922 21306 3978
rect 21374 3922 21430 3978
rect 21498 3922 21554 3978
rect 21622 3922 21678 3978
rect 21250 -216 21306 -160
rect 21374 -216 21430 -160
rect 21498 -216 21554 -160
rect 21622 -216 21678 -160
rect 21250 -340 21306 -284
rect 21374 -340 21430 -284
rect 21498 -340 21554 -284
rect 21622 -340 21678 -284
rect 21250 -464 21306 -408
rect 21374 -464 21430 -408
rect 21498 -464 21554 -408
rect 21622 -464 21678 -408
rect 21250 -588 21306 -532
rect 21374 -588 21430 -532
rect 21498 -588 21554 -532
rect 21622 -588 21678 -532
rect 24970 100294 25026 100350
rect 25094 100294 25150 100350
rect 25218 100294 25274 100350
rect 25342 100294 25398 100350
rect 24970 100170 25026 100226
rect 25094 100170 25150 100226
rect 25218 100170 25274 100226
rect 25342 100170 25398 100226
rect 24970 100046 25026 100102
rect 25094 100046 25150 100102
rect 25218 100046 25274 100102
rect 25342 100046 25398 100102
rect 24970 99922 25026 99978
rect 25094 99922 25150 99978
rect 25218 99922 25274 99978
rect 25342 99922 25398 99978
rect 39250 580294 39306 580350
rect 39374 580294 39430 580350
rect 39498 580294 39554 580350
rect 39622 580294 39678 580350
rect 39250 580170 39306 580226
rect 39374 580170 39430 580226
rect 39498 580170 39554 580226
rect 39622 580170 39678 580226
rect 39250 580046 39306 580102
rect 39374 580046 39430 580102
rect 39498 580046 39554 580102
rect 39622 580046 39678 580102
rect 39250 579922 39306 579978
rect 39374 579922 39430 579978
rect 39498 579922 39554 579978
rect 39622 579922 39678 579978
rect 39250 562294 39306 562350
rect 39374 562294 39430 562350
rect 39498 562294 39554 562350
rect 39622 562294 39678 562350
rect 39250 562170 39306 562226
rect 39374 562170 39430 562226
rect 39498 562170 39554 562226
rect 39622 562170 39678 562226
rect 39250 562046 39306 562102
rect 39374 562046 39430 562102
rect 39498 562046 39554 562102
rect 39622 562046 39678 562102
rect 39250 561922 39306 561978
rect 39374 561922 39430 561978
rect 39498 561922 39554 561978
rect 39622 561922 39678 561978
rect 39250 544294 39306 544350
rect 39374 544294 39430 544350
rect 39498 544294 39554 544350
rect 39622 544294 39678 544350
rect 39250 544170 39306 544226
rect 39374 544170 39430 544226
rect 39498 544170 39554 544226
rect 39622 544170 39678 544226
rect 39250 544046 39306 544102
rect 39374 544046 39430 544102
rect 39498 544046 39554 544102
rect 39622 544046 39678 544102
rect 39250 543922 39306 543978
rect 39374 543922 39430 543978
rect 39498 543922 39554 543978
rect 39622 543922 39678 543978
rect 39250 526294 39306 526350
rect 39374 526294 39430 526350
rect 39498 526294 39554 526350
rect 39622 526294 39678 526350
rect 39250 526170 39306 526226
rect 39374 526170 39430 526226
rect 39498 526170 39554 526226
rect 39622 526170 39678 526226
rect 39250 526046 39306 526102
rect 39374 526046 39430 526102
rect 39498 526046 39554 526102
rect 39622 526046 39678 526102
rect 39250 525922 39306 525978
rect 39374 525922 39430 525978
rect 39498 525922 39554 525978
rect 39622 525922 39678 525978
rect 39250 508294 39306 508350
rect 39374 508294 39430 508350
rect 39498 508294 39554 508350
rect 39622 508294 39678 508350
rect 39250 508170 39306 508226
rect 39374 508170 39430 508226
rect 39498 508170 39554 508226
rect 39622 508170 39678 508226
rect 39250 508046 39306 508102
rect 39374 508046 39430 508102
rect 39498 508046 39554 508102
rect 39622 508046 39678 508102
rect 39250 507922 39306 507978
rect 39374 507922 39430 507978
rect 39498 507922 39554 507978
rect 39622 507922 39678 507978
rect 39250 490294 39306 490350
rect 39374 490294 39430 490350
rect 39498 490294 39554 490350
rect 39622 490294 39678 490350
rect 39250 490170 39306 490226
rect 39374 490170 39430 490226
rect 39498 490170 39554 490226
rect 39622 490170 39678 490226
rect 39250 490046 39306 490102
rect 39374 490046 39430 490102
rect 39498 490046 39554 490102
rect 39622 490046 39678 490102
rect 39250 489922 39306 489978
rect 39374 489922 39430 489978
rect 39498 489922 39554 489978
rect 39622 489922 39678 489978
rect 39250 472294 39306 472350
rect 39374 472294 39430 472350
rect 39498 472294 39554 472350
rect 39622 472294 39678 472350
rect 39250 472170 39306 472226
rect 39374 472170 39430 472226
rect 39498 472170 39554 472226
rect 39622 472170 39678 472226
rect 39250 472046 39306 472102
rect 39374 472046 39430 472102
rect 39498 472046 39554 472102
rect 39622 472046 39678 472102
rect 39250 471922 39306 471978
rect 39374 471922 39430 471978
rect 39498 471922 39554 471978
rect 39622 471922 39678 471978
rect 39250 454294 39306 454350
rect 39374 454294 39430 454350
rect 39498 454294 39554 454350
rect 39622 454294 39678 454350
rect 39250 454170 39306 454226
rect 39374 454170 39430 454226
rect 39498 454170 39554 454226
rect 39622 454170 39678 454226
rect 39250 454046 39306 454102
rect 39374 454046 39430 454102
rect 39498 454046 39554 454102
rect 39622 454046 39678 454102
rect 39250 453922 39306 453978
rect 39374 453922 39430 453978
rect 39498 453922 39554 453978
rect 39622 453922 39678 453978
rect 39250 436294 39306 436350
rect 39374 436294 39430 436350
rect 39498 436294 39554 436350
rect 39622 436294 39678 436350
rect 39250 436170 39306 436226
rect 39374 436170 39430 436226
rect 39498 436170 39554 436226
rect 39622 436170 39678 436226
rect 39250 436046 39306 436102
rect 39374 436046 39430 436102
rect 39498 436046 39554 436102
rect 39622 436046 39678 436102
rect 39250 435922 39306 435978
rect 39374 435922 39430 435978
rect 39498 435922 39554 435978
rect 39622 435922 39678 435978
rect 39250 418294 39306 418350
rect 39374 418294 39430 418350
rect 39498 418294 39554 418350
rect 39622 418294 39678 418350
rect 39250 418170 39306 418226
rect 39374 418170 39430 418226
rect 39498 418170 39554 418226
rect 39622 418170 39678 418226
rect 39250 418046 39306 418102
rect 39374 418046 39430 418102
rect 39498 418046 39554 418102
rect 39622 418046 39678 418102
rect 39250 417922 39306 417978
rect 39374 417922 39430 417978
rect 39498 417922 39554 417978
rect 39622 417922 39678 417978
rect 39250 400294 39306 400350
rect 39374 400294 39430 400350
rect 39498 400294 39554 400350
rect 39622 400294 39678 400350
rect 39250 400170 39306 400226
rect 39374 400170 39430 400226
rect 39498 400170 39554 400226
rect 39622 400170 39678 400226
rect 39250 400046 39306 400102
rect 39374 400046 39430 400102
rect 39498 400046 39554 400102
rect 39622 400046 39678 400102
rect 39250 399922 39306 399978
rect 39374 399922 39430 399978
rect 39498 399922 39554 399978
rect 39622 399922 39678 399978
rect 39250 382294 39306 382350
rect 39374 382294 39430 382350
rect 39498 382294 39554 382350
rect 39622 382294 39678 382350
rect 39250 382170 39306 382226
rect 39374 382170 39430 382226
rect 39498 382170 39554 382226
rect 39622 382170 39678 382226
rect 39250 382046 39306 382102
rect 39374 382046 39430 382102
rect 39498 382046 39554 382102
rect 39622 382046 39678 382102
rect 39250 381922 39306 381978
rect 39374 381922 39430 381978
rect 39498 381922 39554 381978
rect 39622 381922 39678 381978
rect 39250 364294 39306 364350
rect 39374 364294 39430 364350
rect 39498 364294 39554 364350
rect 39622 364294 39678 364350
rect 39250 364170 39306 364226
rect 39374 364170 39430 364226
rect 39498 364170 39554 364226
rect 39622 364170 39678 364226
rect 39250 364046 39306 364102
rect 39374 364046 39430 364102
rect 39498 364046 39554 364102
rect 39622 364046 39678 364102
rect 39250 363922 39306 363978
rect 39374 363922 39430 363978
rect 39498 363922 39554 363978
rect 39622 363922 39678 363978
rect 39250 346294 39306 346350
rect 39374 346294 39430 346350
rect 39498 346294 39554 346350
rect 39622 346294 39678 346350
rect 39250 346170 39306 346226
rect 39374 346170 39430 346226
rect 39498 346170 39554 346226
rect 39622 346170 39678 346226
rect 39250 346046 39306 346102
rect 39374 346046 39430 346102
rect 39498 346046 39554 346102
rect 39622 346046 39678 346102
rect 39250 345922 39306 345978
rect 39374 345922 39430 345978
rect 39498 345922 39554 345978
rect 39622 345922 39678 345978
rect 39250 328294 39306 328350
rect 39374 328294 39430 328350
rect 39498 328294 39554 328350
rect 39622 328294 39678 328350
rect 39250 328170 39306 328226
rect 39374 328170 39430 328226
rect 39498 328170 39554 328226
rect 39622 328170 39678 328226
rect 39250 328046 39306 328102
rect 39374 328046 39430 328102
rect 39498 328046 39554 328102
rect 39622 328046 39678 328102
rect 39250 327922 39306 327978
rect 39374 327922 39430 327978
rect 39498 327922 39554 327978
rect 39622 327922 39678 327978
rect 39250 310294 39306 310350
rect 39374 310294 39430 310350
rect 39498 310294 39554 310350
rect 39622 310294 39678 310350
rect 39250 310170 39306 310226
rect 39374 310170 39430 310226
rect 39498 310170 39554 310226
rect 39622 310170 39678 310226
rect 39250 310046 39306 310102
rect 39374 310046 39430 310102
rect 39498 310046 39554 310102
rect 39622 310046 39678 310102
rect 39250 309922 39306 309978
rect 39374 309922 39430 309978
rect 39498 309922 39554 309978
rect 39622 309922 39678 309978
rect 39250 292294 39306 292350
rect 39374 292294 39430 292350
rect 39498 292294 39554 292350
rect 39622 292294 39678 292350
rect 39250 292170 39306 292226
rect 39374 292170 39430 292226
rect 39498 292170 39554 292226
rect 39622 292170 39678 292226
rect 39250 292046 39306 292102
rect 39374 292046 39430 292102
rect 39498 292046 39554 292102
rect 39622 292046 39678 292102
rect 39250 291922 39306 291978
rect 39374 291922 39430 291978
rect 39498 291922 39554 291978
rect 39622 291922 39678 291978
rect 39250 274294 39306 274350
rect 39374 274294 39430 274350
rect 39498 274294 39554 274350
rect 39622 274294 39678 274350
rect 39250 274170 39306 274226
rect 39374 274170 39430 274226
rect 39498 274170 39554 274226
rect 39622 274170 39678 274226
rect 39250 274046 39306 274102
rect 39374 274046 39430 274102
rect 39498 274046 39554 274102
rect 39622 274046 39678 274102
rect 39250 273922 39306 273978
rect 39374 273922 39430 273978
rect 39498 273922 39554 273978
rect 39622 273922 39678 273978
rect 39250 256294 39306 256350
rect 39374 256294 39430 256350
rect 39498 256294 39554 256350
rect 39622 256294 39678 256350
rect 39250 256170 39306 256226
rect 39374 256170 39430 256226
rect 39498 256170 39554 256226
rect 39622 256170 39678 256226
rect 39250 256046 39306 256102
rect 39374 256046 39430 256102
rect 39498 256046 39554 256102
rect 39622 256046 39678 256102
rect 39250 255922 39306 255978
rect 39374 255922 39430 255978
rect 39498 255922 39554 255978
rect 39622 255922 39678 255978
rect 39250 238294 39306 238350
rect 39374 238294 39430 238350
rect 39498 238294 39554 238350
rect 39622 238294 39678 238350
rect 39250 238170 39306 238226
rect 39374 238170 39430 238226
rect 39498 238170 39554 238226
rect 39622 238170 39678 238226
rect 39250 238046 39306 238102
rect 39374 238046 39430 238102
rect 39498 238046 39554 238102
rect 39622 238046 39678 238102
rect 39250 237922 39306 237978
rect 39374 237922 39430 237978
rect 39498 237922 39554 237978
rect 39622 237922 39678 237978
rect 39250 220294 39306 220350
rect 39374 220294 39430 220350
rect 39498 220294 39554 220350
rect 39622 220294 39678 220350
rect 39250 220170 39306 220226
rect 39374 220170 39430 220226
rect 39498 220170 39554 220226
rect 39622 220170 39678 220226
rect 39250 220046 39306 220102
rect 39374 220046 39430 220102
rect 39498 220046 39554 220102
rect 39622 220046 39678 220102
rect 39250 219922 39306 219978
rect 39374 219922 39430 219978
rect 39498 219922 39554 219978
rect 39622 219922 39678 219978
rect 39250 202294 39306 202350
rect 39374 202294 39430 202350
rect 39498 202294 39554 202350
rect 39622 202294 39678 202350
rect 39250 202170 39306 202226
rect 39374 202170 39430 202226
rect 39498 202170 39554 202226
rect 39622 202170 39678 202226
rect 39250 202046 39306 202102
rect 39374 202046 39430 202102
rect 39498 202046 39554 202102
rect 39622 202046 39678 202102
rect 39250 201922 39306 201978
rect 39374 201922 39430 201978
rect 39498 201922 39554 201978
rect 39622 201922 39678 201978
rect 42970 598116 43026 598172
rect 43094 598116 43150 598172
rect 43218 598116 43274 598172
rect 43342 598116 43398 598172
rect 42970 597992 43026 598048
rect 43094 597992 43150 598048
rect 43218 597992 43274 598048
rect 43342 597992 43398 598048
rect 42970 597868 43026 597924
rect 43094 597868 43150 597924
rect 43218 597868 43274 597924
rect 43342 597868 43398 597924
rect 42970 597744 43026 597800
rect 43094 597744 43150 597800
rect 43218 597744 43274 597800
rect 43342 597744 43398 597800
rect 42970 586294 43026 586350
rect 43094 586294 43150 586350
rect 43218 586294 43274 586350
rect 43342 586294 43398 586350
rect 42970 586170 43026 586226
rect 43094 586170 43150 586226
rect 43218 586170 43274 586226
rect 43342 586170 43398 586226
rect 42970 586046 43026 586102
rect 43094 586046 43150 586102
rect 43218 586046 43274 586102
rect 43342 586046 43398 586102
rect 42970 585922 43026 585978
rect 43094 585922 43150 585978
rect 43218 585922 43274 585978
rect 43342 585922 43398 585978
rect 42970 568294 43026 568350
rect 43094 568294 43150 568350
rect 43218 568294 43274 568350
rect 43342 568294 43398 568350
rect 42970 568170 43026 568226
rect 43094 568170 43150 568226
rect 43218 568170 43274 568226
rect 43342 568170 43398 568226
rect 42970 568046 43026 568102
rect 43094 568046 43150 568102
rect 43218 568046 43274 568102
rect 43342 568046 43398 568102
rect 42970 567922 43026 567978
rect 43094 567922 43150 567978
rect 43218 567922 43274 567978
rect 43342 567922 43398 567978
rect 42970 550294 43026 550350
rect 43094 550294 43150 550350
rect 43218 550294 43274 550350
rect 43342 550294 43398 550350
rect 42970 550170 43026 550226
rect 43094 550170 43150 550226
rect 43218 550170 43274 550226
rect 43342 550170 43398 550226
rect 42970 550046 43026 550102
rect 43094 550046 43150 550102
rect 43218 550046 43274 550102
rect 43342 550046 43398 550102
rect 42970 549922 43026 549978
rect 43094 549922 43150 549978
rect 43218 549922 43274 549978
rect 43342 549922 43398 549978
rect 42970 532294 43026 532350
rect 43094 532294 43150 532350
rect 43218 532294 43274 532350
rect 43342 532294 43398 532350
rect 42970 532170 43026 532226
rect 43094 532170 43150 532226
rect 43218 532170 43274 532226
rect 43342 532170 43398 532226
rect 42970 532046 43026 532102
rect 43094 532046 43150 532102
rect 43218 532046 43274 532102
rect 43342 532046 43398 532102
rect 42970 531922 43026 531978
rect 43094 531922 43150 531978
rect 43218 531922 43274 531978
rect 43342 531922 43398 531978
rect 42970 514294 43026 514350
rect 43094 514294 43150 514350
rect 43218 514294 43274 514350
rect 43342 514294 43398 514350
rect 42970 514170 43026 514226
rect 43094 514170 43150 514226
rect 43218 514170 43274 514226
rect 43342 514170 43398 514226
rect 42970 514046 43026 514102
rect 43094 514046 43150 514102
rect 43218 514046 43274 514102
rect 43342 514046 43398 514102
rect 42970 513922 43026 513978
rect 43094 513922 43150 513978
rect 43218 513922 43274 513978
rect 43342 513922 43398 513978
rect 42970 496294 43026 496350
rect 43094 496294 43150 496350
rect 43218 496294 43274 496350
rect 43342 496294 43398 496350
rect 42970 496170 43026 496226
rect 43094 496170 43150 496226
rect 43218 496170 43274 496226
rect 43342 496170 43398 496226
rect 42970 496046 43026 496102
rect 43094 496046 43150 496102
rect 43218 496046 43274 496102
rect 43342 496046 43398 496102
rect 42970 495922 43026 495978
rect 43094 495922 43150 495978
rect 43218 495922 43274 495978
rect 43342 495922 43398 495978
rect 42970 478294 43026 478350
rect 43094 478294 43150 478350
rect 43218 478294 43274 478350
rect 43342 478294 43398 478350
rect 42970 478170 43026 478226
rect 43094 478170 43150 478226
rect 43218 478170 43274 478226
rect 43342 478170 43398 478226
rect 42970 478046 43026 478102
rect 43094 478046 43150 478102
rect 43218 478046 43274 478102
rect 43342 478046 43398 478102
rect 42970 477922 43026 477978
rect 43094 477922 43150 477978
rect 43218 477922 43274 477978
rect 43342 477922 43398 477978
rect 42970 460294 43026 460350
rect 43094 460294 43150 460350
rect 43218 460294 43274 460350
rect 43342 460294 43398 460350
rect 42970 460170 43026 460226
rect 43094 460170 43150 460226
rect 43218 460170 43274 460226
rect 43342 460170 43398 460226
rect 42970 460046 43026 460102
rect 43094 460046 43150 460102
rect 43218 460046 43274 460102
rect 43342 460046 43398 460102
rect 42970 459922 43026 459978
rect 43094 459922 43150 459978
rect 43218 459922 43274 459978
rect 43342 459922 43398 459978
rect 42970 442294 43026 442350
rect 43094 442294 43150 442350
rect 43218 442294 43274 442350
rect 43342 442294 43398 442350
rect 42970 442170 43026 442226
rect 43094 442170 43150 442226
rect 43218 442170 43274 442226
rect 43342 442170 43398 442226
rect 42970 442046 43026 442102
rect 43094 442046 43150 442102
rect 43218 442046 43274 442102
rect 43342 442046 43398 442102
rect 42970 441922 43026 441978
rect 43094 441922 43150 441978
rect 43218 441922 43274 441978
rect 43342 441922 43398 441978
rect 42970 424294 43026 424350
rect 43094 424294 43150 424350
rect 43218 424294 43274 424350
rect 43342 424294 43398 424350
rect 42970 424170 43026 424226
rect 43094 424170 43150 424226
rect 43218 424170 43274 424226
rect 43342 424170 43398 424226
rect 42970 424046 43026 424102
rect 43094 424046 43150 424102
rect 43218 424046 43274 424102
rect 43342 424046 43398 424102
rect 42970 423922 43026 423978
rect 43094 423922 43150 423978
rect 43218 423922 43274 423978
rect 43342 423922 43398 423978
rect 42970 406294 43026 406350
rect 43094 406294 43150 406350
rect 43218 406294 43274 406350
rect 43342 406294 43398 406350
rect 42970 406170 43026 406226
rect 43094 406170 43150 406226
rect 43218 406170 43274 406226
rect 43342 406170 43398 406226
rect 42970 406046 43026 406102
rect 43094 406046 43150 406102
rect 43218 406046 43274 406102
rect 43342 406046 43398 406102
rect 42970 405922 43026 405978
rect 43094 405922 43150 405978
rect 43218 405922 43274 405978
rect 43342 405922 43398 405978
rect 42970 388294 43026 388350
rect 43094 388294 43150 388350
rect 43218 388294 43274 388350
rect 43342 388294 43398 388350
rect 42970 388170 43026 388226
rect 43094 388170 43150 388226
rect 43218 388170 43274 388226
rect 43342 388170 43398 388226
rect 42970 388046 43026 388102
rect 43094 388046 43150 388102
rect 43218 388046 43274 388102
rect 43342 388046 43398 388102
rect 42970 387922 43026 387978
rect 43094 387922 43150 387978
rect 43218 387922 43274 387978
rect 43342 387922 43398 387978
rect 42970 370294 43026 370350
rect 43094 370294 43150 370350
rect 43218 370294 43274 370350
rect 43342 370294 43398 370350
rect 42970 370170 43026 370226
rect 43094 370170 43150 370226
rect 43218 370170 43274 370226
rect 43342 370170 43398 370226
rect 42970 370046 43026 370102
rect 43094 370046 43150 370102
rect 43218 370046 43274 370102
rect 43342 370046 43398 370102
rect 42970 369922 43026 369978
rect 43094 369922 43150 369978
rect 43218 369922 43274 369978
rect 43342 369922 43398 369978
rect 42970 352294 43026 352350
rect 43094 352294 43150 352350
rect 43218 352294 43274 352350
rect 43342 352294 43398 352350
rect 42970 352170 43026 352226
rect 43094 352170 43150 352226
rect 43218 352170 43274 352226
rect 43342 352170 43398 352226
rect 42970 352046 43026 352102
rect 43094 352046 43150 352102
rect 43218 352046 43274 352102
rect 43342 352046 43398 352102
rect 42970 351922 43026 351978
rect 43094 351922 43150 351978
rect 43218 351922 43274 351978
rect 43342 351922 43398 351978
rect 42970 334294 43026 334350
rect 43094 334294 43150 334350
rect 43218 334294 43274 334350
rect 43342 334294 43398 334350
rect 42970 334170 43026 334226
rect 43094 334170 43150 334226
rect 43218 334170 43274 334226
rect 43342 334170 43398 334226
rect 42970 334046 43026 334102
rect 43094 334046 43150 334102
rect 43218 334046 43274 334102
rect 43342 334046 43398 334102
rect 42970 333922 43026 333978
rect 43094 333922 43150 333978
rect 43218 333922 43274 333978
rect 43342 333922 43398 333978
rect 42970 316294 43026 316350
rect 43094 316294 43150 316350
rect 43218 316294 43274 316350
rect 43342 316294 43398 316350
rect 42970 316170 43026 316226
rect 43094 316170 43150 316226
rect 43218 316170 43274 316226
rect 43342 316170 43398 316226
rect 42970 316046 43026 316102
rect 43094 316046 43150 316102
rect 43218 316046 43274 316102
rect 43342 316046 43398 316102
rect 42970 315922 43026 315978
rect 43094 315922 43150 315978
rect 43218 315922 43274 315978
rect 43342 315922 43398 315978
rect 42970 298294 43026 298350
rect 43094 298294 43150 298350
rect 43218 298294 43274 298350
rect 43342 298294 43398 298350
rect 42970 298170 43026 298226
rect 43094 298170 43150 298226
rect 43218 298170 43274 298226
rect 43342 298170 43398 298226
rect 42970 298046 43026 298102
rect 43094 298046 43150 298102
rect 43218 298046 43274 298102
rect 43342 298046 43398 298102
rect 42970 297922 43026 297978
rect 43094 297922 43150 297978
rect 43218 297922 43274 297978
rect 43342 297922 43398 297978
rect 42970 280294 43026 280350
rect 43094 280294 43150 280350
rect 43218 280294 43274 280350
rect 43342 280294 43398 280350
rect 42970 280170 43026 280226
rect 43094 280170 43150 280226
rect 43218 280170 43274 280226
rect 43342 280170 43398 280226
rect 42970 280046 43026 280102
rect 43094 280046 43150 280102
rect 43218 280046 43274 280102
rect 43342 280046 43398 280102
rect 42970 279922 43026 279978
rect 43094 279922 43150 279978
rect 43218 279922 43274 279978
rect 43342 279922 43398 279978
rect 42970 262294 43026 262350
rect 43094 262294 43150 262350
rect 43218 262294 43274 262350
rect 43342 262294 43398 262350
rect 42970 262170 43026 262226
rect 43094 262170 43150 262226
rect 43218 262170 43274 262226
rect 43342 262170 43398 262226
rect 42970 262046 43026 262102
rect 43094 262046 43150 262102
rect 43218 262046 43274 262102
rect 43342 262046 43398 262102
rect 42970 261922 43026 261978
rect 43094 261922 43150 261978
rect 43218 261922 43274 261978
rect 43342 261922 43398 261978
rect 42970 244294 43026 244350
rect 43094 244294 43150 244350
rect 43218 244294 43274 244350
rect 43342 244294 43398 244350
rect 42970 244170 43026 244226
rect 43094 244170 43150 244226
rect 43218 244170 43274 244226
rect 43342 244170 43398 244226
rect 42970 244046 43026 244102
rect 43094 244046 43150 244102
rect 43218 244046 43274 244102
rect 43342 244046 43398 244102
rect 42970 243922 43026 243978
rect 43094 243922 43150 243978
rect 43218 243922 43274 243978
rect 43342 243922 43398 243978
rect 57250 597156 57306 597212
rect 57374 597156 57430 597212
rect 57498 597156 57554 597212
rect 57622 597156 57678 597212
rect 57250 597032 57306 597088
rect 57374 597032 57430 597088
rect 57498 597032 57554 597088
rect 57622 597032 57678 597088
rect 57250 596908 57306 596964
rect 57374 596908 57430 596964
rect 57498 596908 57554 596964
rect 57622 596908 57678 596964
rect 57250 596784 57306 596840
rect 57374 596784 57430 596840
rect 57498 596784 57554 596840
rect 57622 596784 57678 596840
rect 57250 580294 57306 580350
rect 57374 580294 57430 580350
rect 57498 580294 57554 580350
rect 57622 580294 57678 580350
rect 57250 580170 57306 580226
rect 57374 580170 57430 580226
rect 57498 580170 57554 580226
rect 57622 580170 57678 580226
rect 57250 580046 57306 580102
rect 57374 580046 57430 580102
rect 57498 580046 57554 580102
rect 57622 580046 57678 580102
rect 57250 579922 57306 579978
rect 57374 579922 57430 579978
rect 57498 579922 57554 579978
rect 57622 579922 57678 579978
rect 57250 562294 57306 562350
rect 57374 562294 57430 562350
rect 57498 562294 57554 562350
rect 57622 562294 57678 562350
rect 57250 562170 57306 562226
rect 57374 562170 57430 562226
rect 57498 562170 57554 562226
rect 57622 562170 57678 562226
rect 57250 562046 57306 562102
rect 57374 562046 57430 562102
rect 57498 562046 57554 562102
rect 57622 562046 57678 562102
rect 57250 561922 57306 561978
rect 57374 561922 57430 561978
rect 57498 561922 57554 561978
rect 57622 561922 57678 561978
rect 57250 544294 57306 544350
rect 57374 544294 57430 544350
rect 57498 544294 57554 544350
rect 57622 544294 57678 544350
rect 57250 544170 57306 544226
rect 57374 544170 57430 544226
rect 57498 544170 57554 544226
rect 57622 544170 57678 544226
rect 57250 544046 57306 544102
rect 57374 544046 57430 544102
rect 57498 544046 57554 544102
rect 57622 544046 57678 544102
rect 57250 543922 57306 543978
rect 57374 543922 57430 543978
rect 57498 543922 57554 543978
rect 57622 543922 57678 543978
rect 57250 526294 57306 526350
rect 57374 526294 57430 526350
rect 57498 526294 57554 526350
rect 57622 526294 57678 526350
rect 57250 526170 57306 526226
rect 57374 526170 57430 526226
rect 57498 526170 57554 526226
rect 57622 526170 57678 526226
rect 57250 526046 57306 526102
rect 57374 526046 57430 526102
rect 57498 526046 57554 526102
rect 57622 526046 57678 526102
rect 57250 525922 57306 525978
rect 57374 525922 57430 525978
rect 57498 525922 57554 525978
rect 57622 525922 57678 525978
rect 57250 508294 57306 508350
rect 57374 508294 57430 508350
rect 57498 508294 57554 508350
rect 57622 508294 57678 508350
rect 57250 508170 57306 508226
rect 57374 508170 57430 508226
rect 57498 508170 57554 508226
rect 57622 508170 57678 508226
rect 57250 508046 57306 508102
rect 57374 508046 57430 508102
rect 57498 508046 57554 508102
rect 57622 508046 57678 508102
rect 57250 507922 57306 507978
rect 57374 507922 57430 507978
rect 57498 507922 57554 507978
rect 57622 507922 57678 507978
rect 57250 490294 57306 490350
rect 57374 490294 57430 490350
rect 57498 490294 57554 490350
rect 57622 490294 57678 490350
rect 57250 490170 57306 490226
rect 57374 490170 57430 490226
rect 57498 490170 57554 490226
rect 57622 490170 57678 490226
rect 57250 490046 57306 490102
rect 57374 490046 57430 490102
rect 57498 490046 57554 490102
rect 57622 490046 57678 490102
rect 57250 489922 57306 489978
rect 57374 489922 57430 489978
rect 57498 489922 57554 489978
rect 57622 489922 57678 489978
rect 57250 472294 57306 472350
rect 57374 472294 57430 472350
rect 57498 472294 57554 472350
rect 57622 472294 57678 472350
rect 57250 472170 57306 472226
rect 57374 472170 57430 472226
rect 57498 472170 57554 472226
rect 57622 472170 57678 472226
rect 57250 472046 57306 472102
rect 57374 472046 57430 472102
rect 57498 472046 57554 472102
rect 57622 472046 57678 472102
rect 57250 471922 57306 471978
rect 57374 471922 57430 471978
rect 57498 471922 57554 471978
rect 57622 471922 57678 471978
rect 57250 454294 57306 454350
rect 57374 454294 57430 454350
rect 57498 454294 57554 454350
rect 57622 454294 57678 454350
rect 57250 454170 57306 454226
rect 57374 454170 57430 454226
rect 57498 454170 57554 454226
rect 57622 454170 57678 454226
rect 57250 454046 57306 454102
rect 57374 454046 57430 454102
rect 57498 454046 57554 454102
rect 57622 454046 57678 454102
rect 57250 453922 57306 453978
rect 57374 453922 57430 453978
rect 57498 453922 57554 453978
rect 57622 453922 57678 453978
rect 57250 436294 57306 436350
rect 57374 436294 57430 436350
rect 57498 436294 57554 436350
rect 57622 436294 57678 436350
rect 57250 436170 57306 436226
rect 57374 436170 57430 436226
rect 57498 436170 57554 436226
rect 57622 436170 57678 436226
rect 57250 436046 57306 436102
rect 57374 436046 57430 436102
rect 57498 436046 57554 436102
rect 57622 436046 57678 436102
rect 57250 435922 57306 435978
rect 57374 435922 57430 435978
rect 57498 435922 57554 435978
rect 57622 435922 57678 435978
rect 57250 418294 57306 418350
rect 57374 418294 57430 418350
rect 57498 418294 57554 418350
rect 57622 418294 57678 418350
rect 57250 418170 57306 418226
rect 57374 418170 57430 418226
rect 57498 418170 57554 418226
rect 57622 418170 57678 418226
rect 57250 418046 57306 418102
rect 57374 418046 57430 418102
rect 57498 418046 57554 418102
rect 57622 418046 57678 418102
rect 57250 417922 57306 417978
rect 57374 417922 57430 417978
rect 57498 417922 57554 417978
rect 57622 417922 57678 417978
rect 57250 400294 57306 400350
rect 57374 400294 57430 400350
rect 57498 400294 57554 400350
rect 57622 400294 57678 400350
rect 57250 400170 57306 400226
rect 57374 400170 57430 400226
rect 57498 400170 57554 400226
rect 57622 400170 57678 400226
rect 57250 400046 57306 400102
rect 57374 400046 57430 400102
rect 57498 400046 57554 400102
rect 57622 400046 57678 400102
rect 57250 399922 57306 399978
rect 57374 399922 57430 399978
rect 57498 399922 57554 399978
rect 57622 399922 57678 399978
rect 57250 382294 57306 382350
rect 57374 382294 57430 382350
rect 57498 382294 57554 382350
rect 57622 382294 57678 382350
rect 57250 382170 57306 382226
rect 57374 382170 57430 382226
rect 57498 382170 57554 382226
rect 57622 382170 57678 382226
rect 57250 382046 57306 382102
rect 57374 382046 57430 382102
rect 57498 382046 57554 382102
rect 57622 382046 57678 382102
rect 57250 381922 57306 381978
rect 57374 381922 57430 381978
rect 57498 381922 57554 381978
rect 57622 381922 57678 381978
rect 57250 364294 57306 364350
rect 57374 364294 57430 364350
rect 57498 364294 57554 364350
rect 57622 364294 57678 364350
rect 57250 364170 57306 364226
rect 57374 364170 57430 364226
rect 57498 364170 57554 364226
rect 57622 364170 57678 364226
rect 57250 364046 57306 364102
rect 57374 364046 57430 364102
rect 57498 364046 57554 364102
rect 57622 364046 57678 364102
rect 57250 363922 57306 363978
rect 57374 363922 57430 363978
rect 57498 363922 57554 363978
rect 57622 363922 57678 363978
rect 57250 346294 57306 346350
rect 57374 346294 57430 346350
rect 57498 346294 57554 346350
rect 57622 346294 57678 346350
rect 57250 346170 57306 346226
rect 57374 346170 57430 346226
rect 57498 346170 57554 346226
rect 57622 346170 57678 346226
rect 57250 346046 57306 346102
rect 57374 346046 57430 346102
rect 57498 346046 57554 346102
rect 57622 346046 57678 346102
rect 57250 345922 57306 345978
rect 57374 345922 57430 345978
rect 57498 345922 57554 345978
rect 57622 345922 57678 345978
rect 57250 328294 57306 328350
rect 57374 328294 57430 328350
rect 57498 328294 57554 328350
rect 57622 328294 57678 328350
rect 57250 328170 57306 328226
rect 57374 328170 57430 328226
rect 57498 328170 57554 328226
rect 57622 328170 57678 328226
rect 57250 328046 57306 328102
rect 57374 328046 57430 328102
rect 57498 328046 57554 328102
rect 57622 328046 57678 328102
rect 57250 327922 57306 327978
rect 57374 327922 57430 327978
rect 57498 327922 57554 327978
rect 57622 327922 57678 327978
rect 57250 310294 57306 310350
rect 57374 310294 57430 310350
rect 57498 310294 57554 310350
rect 57622 310294 57678 310350
rect 57250 310170 57306 310226
rect 57374 310170 57430 310226
rect 57498 310170 57554 310226
rect 57622 310170 57678 310226
rect 57250 310046 57306 310102
rect 57374 310046 57430 310102
rect 57498 310046 57554 310102
rect 57622 310046 57678 310102
rect 57250 309922 57306 309978
rect 57374 309922 57430 309978
rect 57498 309922 57554 309978
rect 57622 309922 57678 309978
rect 57250 292294 57306 292350
rect 57374 292294 57430 292350
rect 57498 292294 57554 292350
rect 57622 292294 57678 292350
rect 57250 292170 57306 292226
rect 57374 292170 57430 292226
rect 57498 292170 57554 292226
rect 57622 292170 57678 292226
rect 57250 292046 57306 292102
rect 57374 292046 57430 292102
rect 57498 292046 57554 292102
rect 57622 292046 57678 292102
rect 57250 291922 57306 291978
rect 57374 291922 57430 291978
rect 57498 291922 57554 291978
rect 57622 291922 57678 291978
rect 57250 274294 57306 274350
rect 57374 274294 57430 274350
rect 57498 274294 57554 274350
rect 57622 274294 57678 274350
rect 57250 274170 57306 274226
rect 57374 274170 57430 274226
rect 57498 274170 57554 274226
rect 57622 274170 57678 274226
rect 57250 274046 57306 274102
rect 57374 274046 57430 274102
rect 57498 274046 57554 274102
rect 57622 274046 57678 274102
rect 57250 273922 57306 273978
rect 57374 273922 57430 273978
rect 57498 273922 57554 273978
rect 57622 273922 57678 273978
rect 57250 256294 57306 256350
rect 57374 256294 57430 256350
rect 57498 256294 57554 256350
rect 57622 256294 57678 256350
rect 57250 256170 57306 256226
rect 57374 256170 57430 256226
rect 57498 256170 57554 256226
rect 57622 256170 57678 256226
rect 57250 256046 57306 256102
rect 57374 256046 57430 256102
rect 57498 256046 57554 256102
rect 57622 256046 57678 256102
rect 57250 255922 57306 255978
rect 57374 255922 57430 255978
rect 57498 255922 57554 255978
rect 57622 255922 57678 255978
rect 57250 238294 57306 238350
rect 57374 238294 57430 238350
rect 57498 238294 57554 238350
rect 57622 238294 57678 238350
rect 57250 238170 57306 238226
rect 57374 238170 57430 238226
rect 57498 238170 57554 238226
rect 57622 238170 57678 238226
rect 57250 238046 57306 238102
rect 57374 238046 57430 238102
rect 57498 238046 57554 238102
rect 57622 238046 57678 238102
rect 57250 237922 57306 237978
rect 57374 237922 57430 237978
rect 57498 237922 57554 237978
rect 57622 237922 57678 237978
rect 42970 226294 43026 226350
rect 43094 226294 43150 226350
rect 43218 226294 43274 226350
rect 43342 226294 43398 226350
rect 42970 226170 43026 226226
rect 43094 226170 43150 226226
rect 43218 226170 43274 226226
rect 43342 226170 43398 226226
rect 42970 226046 43026 226102
rect 43094 226046 43150 226102
rect 43218 226046 43274 226102
rect 43342 226046 43398 226102
rect 42970 225922 43026 225978
rect 43094 225922 43150 225978
rect 43218 225922 43274 225978
rect 43342 225922 43398 225978
rect 42970 208294 43026 208350
rect 43094 208294 43150 208350
rect 43218 208294 43274 208350
rect 43342 208294 43398 208350
rect 42970 208170 43026 208226
rect 43094 208170 43150 208226
rect 43218 208170 43274 208226
rect 43342 208170 43398 208226
rect 42970 208046 43026 208102
rect 43094 208046 43150 208102
rect 43218 208046 43274 208102
rect 43342 208046 43398 208102
rect 42970 207922 43026 207978
rect 43094 207922 43150 207978
rect 43218 207922 43274 207978
rect 43342 207922 43398 207978
rect 39250 184294 39306 184350
rect 39374 184294 39430 184350
rect 39498 184294 39554 184350
rect 39622 184294 39678 184350
rect 39250 184170 39306 184226
rect 39374 184170 39430 184226
rect 39498 184170 39554 184226
rect 39622 184170 39678 184226
rect 39250 184046 39306 184102
rect 39374 184046 39430 184102
rect 39498 184046 39554 184102
rect 39622 184046 39678 184102
rect 39250 183922 39306 183978
rect 39374 183922 39430 183978
rect 39498 183922 39554 183978
rect 39622 183922 39678 183978
rect 39250 166294 39306 166350
rect 39374 166294 39430 166350
rect 39498 166294 39554 166350
rect 39622 166294 39678 166350
rect 39250 166170 39306 166226
rect 39374 166170 39430 166226
rect 39498 166170 39554 166226
rect 39622 166170 39678 166226
rect 39250 166046 39306 166102
rect 39374 166046 39430 166102
rect 39498 166046 39554 166102
rect 39622 166046 39678 166102
rect 39250 165922 39306 165978
rect 39374 165922 39430 165978
rect 39498 165922 39554 165978
rect 39622 165922 39678 165978
rect 39250 148294 39306 148350
rect 39374 148294 39430 148350
rect 39498 148294 39554 148350
rect 39622 148294 39678 148350
rect 39250 148170 39306 148226
rect 39374 148170 39430 148226
rect 39498 148170 39554 148226
rect 39622 148170 39678 148226
rect 39250 148046 39306 148102
rect 39374 148046 39430 148102
rect 39498 148046 39554 148102
rect 39622 148046 39678 148102
rect 39250 147922 39306 147978
rect 39374 147922 39430 147978
rect 39498 147922 39554 147978
rect 39622 147922 39678 147978
rect 39250 130294 39306 130350
rect 39374 130294 39430 130350
rect 39498 130294 39554 130350
rect 39622 130294 39678 130350
rect 39250 130170 39306 130226
rect 39374 130170 39430 130226
rect 39498 130170 39554 130226
rect 39622 130170 39678 130226
rect 39250 130046 39306 130102
rect 39374 130046 39430 130102
rect 39498 130046 39554 130102
rect 39622 130046 39678 130102
rect 39250 129922 39306 129978
rect 39374 129922 39430 129978
rect 39498 129922 39554 129978
rect 39622 129922 39678 129978
rect 39250 112294 39306 112350
rect 39374 112294 39430 112350
rect 39498 112294 39554 112350
rect 39622 112294 39678 112350
rect 39250 112170 39306 112226
rect 39374 112170 39430 112226
rect 39498 112170 39554 112226
rect 39622 112170 39678 112226
rect 39250 112046 39306 112102
rect 39374 112046 39430 112102
rect 39498 112046 39554 112102
rect 39622 112046 39678 112102
rect 39250 111922 39306 111978
rect 39374 111922 39430 111978
rect 39498 111922 39554 111978
rect 39622 111922 39678 111978
rect 39250 94294 39306 94350
rect 39374 94294 39430 94350
rect 39498 94294 39554 94350
rect 39622 94294 39678 94350
rect 39250 94170 39306 94226
rect 39374 94170 39430 94226
rect 39498 94170 39554 94226
rect 39622 94170 39678 94226
rect 39250 94046 39306 94102
rect 39374 94046 39430 94102
rect 39498 94046 39554 94102
rect 39622 94046 39678 94102
rect 39250 93922 39306 93978
rect 39374 93922 39430 93978
rect 39498 93922 39554 93978
rect 39622 93922 39678 93978
rect 24970 82294 25026 82350
rect 25094 82294 25150 82350
rect 25218 82294 25274 82350
rect 25342 82294 25398 82350
rect 24970 82170 25026 82226
rect 25094 82170 25150 82226
rect 25218 82170 25274 82226
rect 25342 82170 25398 82226
rect 24970 82046 25026 82102
rect 25094 82046 25150 82102
rect 25218 82046 25274 82102
rect 25342 82046 25398 82102
rect 24970 81922 25026 81978
rect 25094 81922 25150 81978
rect 25218 81922 25274 81978
rect 25342 81922 25398 81978
rect 24970 64294 25026 64350
rect 25094 64294 25150 64350
rect 25218 64294 25274 64350
rect 25342 64294 25398 64350
rect 24970 64170 25026 64226
rect 25094 64170 25150 64226
rect 25218 64170 25274 64226
rect 25342 64170 25398 64226
rect 24970 64046 25026 64102
rect 25094 64046 25150 64102
rect 25218 64046 25274 64102
rect 25342 64046 25398 64102
rect 24970 63922 25026 63978
rect 25094 63922 25150 63978
rect 25218 63922 25274 63978
rect 25342 63922 25398 63978
rect 24970 46294 25026 46350
rect 25094 46294 25150 46350
rect 25218 46294 25274 46350
rect 25342 46294 25398 46350
rect 24970 46170 25026 46226
rect 25094 46170 25150 46226
rect 25218 46170 25274 46226
rect 25342 46170 25398 46226
rect 24970 46046 25026 46102
rect 25094 46046 25150 46102
rect 25218 46046 25274 46102
rect 25342 46046 25398 46102
rect 24970 45922 25026 45978
rect 25094 45922 25150 45978
rect 25218 45922 25274 45978
rect 25342 45922 25398 45978
rect 24970 28294 25026 28350
rect 25094 28294 25150 28350
rect 25218 28294 25274 28350
rect 25342 28294 25398 28350
rect 24970 28170 25026 28226
rect 25094 28170 25150 28226
rect 25218 28170 25274 28226
rect 25342 28170 25398 28226
rect 24970 28046 25026 28102
rect 25094 28046 25150 28102
rect 25218 28046 25274 28102
rect 25342 28046 25398 28102
rect 24970 27922 25026 27978
rect 25094 27922 25150 27978
rect 25218 27922 25274 27978
rect 25342 27922 25398 27978
rect 24970 10294 25026 10350
rect 25094 10294 25150 10350
rect 25218 10294 25274 10350
rect 25342 10294 25398 10350
rect 24970 10170 25026 10226
rect 25094 10170 25150 10226
rect 25218 10170 25274 10226
rect 25342 10170 25398 10226
rect 24970 10046 25026 10102
rect 25094 10046 25150 10102
rect 25218 10046 25274 10102
rect 25342 10046 25398 10102
rect 24970 9922 25026 9978
rect 25094 9922 25150 9978
rect 25218 9922 25274 9978
rect 25342 9922 25398 9978
rect 24970 -1176 25026 -1120
rect 25094 -1176 25150 -1120
rect 25218 -1176 25274 -1120
rect 25342 -1176 25398 -1120
rect 24970 -1300 25026 -1244
rect 25094 -1300 25150 -1244
rect 25218 -1300 25274 -1244
rect 25342 -1300 25398 -1244
rect 24970 -1424 25026 -1368
rect 25094 -1424 25150 -1368
rect 25218 -1424 25274 -1368
rect 25342 -1424 25398 -1368
rect 24970 -1548 25026 -1492
rect 25094 -1548 25150 -1492
rect 25218 -1548 25274 -1492
rect 25342 -1548 25398 -1492
rect 42970 190294 43026 190350
rect 43094 190294 43150 190350
rect 43218 190294 43274 190350
rect 43342 190294 43398 190350
rect 42970 190170 43026 190226
rect 43094 190170 43150 190226
rect 43218 190170 43274 190226
rect 43342 190170 43398 190226
rect 42970 190046 43026 190102
rect 43094 190046 43150 190102
rect 43218 190046 43274 190102
rect 43342 190046 43398 190102
rect 42970 189922 43026 189978
rect 43094 189922 43150 189978
rect 43218 189922 43274 189978
rect 43342 189922 43398 189978
rect 42970 172294 43026 172350
rect 43094 172294 43150 172350
rect 43218 172294 43274 172350
rect 43342 172294 43398 172350
rect 42970 172170 43026 172226
rect 43094 172170 43150 172226
rect 43218 172170 43274 172226
rect 43342 172170 43398 172226
rect 42970 172046 43026 172102
rect 43094 172046 43150 172102
rect 43218 172046 43274 172102
rect 43342 172046 43398 172102
rect 42970 171922 43026 171978
rect 43094 171922 43150 171978
rect 43218 171922 43274 171978
rect 43342 171922 43398 171978
rect 42970 154294 43026 154350
rect 43094 154294 43150 154350
rect 43218 154294 43274 154350
rect 43342 154294 43398 154350
rect 42970 154170 43026 154226
rect 43094 154170 43150 154226
rect 43218 154170 43274 154226
rect 43342 154170 43398 154226
rect 42970 154046 43026 154102
rect 43094 154046 43150 154102
rect 43218 154046 43274 154102
rect 43342 154046 43398 154102
rect 42970 153922 43026 153978
rect 43094 153922 43150 153978
rect 43218 153922 43274 153978
rect 43342 153922 43398 153978
rect 42970 136294 43026 136350
rect 43094 136294 43150 136350
rect 43218 136294 43274 136350
rect 43342 136294 43398 136350
rect 42970 136170 43026 136226
rect 43094 136170 43150 136226
rect 43218 136170 43274 136226
rect 43342 136170 43398 136226
rect 42970 136046 43026 136102
rect 43094 136046 43150 136102
rect 43218 136046 43274 136102
rect 43342 136046 43398 136102
rect 42970 135922 43026 135978
rect 43094 135922 43150 135978
rect 43218 135922 43274 135978
rect 43342 135922 43398 135978
rect 42970 118294 43026 118350
rect 43094 118294 43150 118350
rect 43218 118294 43274 118350
rect 43342 118294 43398 118350
rect 42970 118170 43026 118226
rect 43094 118170 43150 118226
rect 43218 118170 43274 118226
rect 43342 118170 43398 118226
rect 42970 118046 43026 118102
rect 43094 118046 43150 118102
rect 43218 118046 43274 118102
rect 43342 118046 43398 118102
rect 42970 117922 43026 117978
rect 43094 117922 43150 117978
rect 43218 117922 43274 117978
rect 43342 117922 43398 117978
rect 42970 100294 43026 100350
rect 43094 100294 43150 100350
rect 43218 100294 43274 100350
rect 43342 100294 43398 100350
rect 42970 100170 43026 100226
rect 43094 100170 43150 100226
rect 43218 100170 43274 100226
rect 43342 100170 43398 100226
rect 42970 100046 43026 100102
rect 43094 100046 43150 100102
rect 43218 100046 43274 100102
rect 43342 100046 43398 100102
rect 42970 99922 43026 99978
rect 43094 99922 43150 99978
rect 43218 99922 43274 99978
rect 43342 99922 43398 99978
rect 39250 76294 39306 76350
rect 39374 76294 39430 76350
rect 39498 76294 39554 76350
rect 39622 76294 39678 76350
rect 39250 76170 39306 76226
rect 39374 76170 39430 76226
rect 39498 76170 39554 76226
rect 39622 76170 39678 76226
rect 39250 76046 39306 76102
rect 39374 76046 39430 76102
rect 39498 76046 39554 76102
rect 39622 76046 39678 76102
rect 39250 75922 39306 75978
rect 39374 75922 39430 75978
rect 39498 75922 39554 75978
rect 39622 75922 39678 75978
rect 39250 58294 39306 58350
rect 39374 58294 39430 58350
rect 39498 58294 39554 58350
rect 39622 58294 39678 58350
rect 39250 58170 39306 58226
rect 39374 58170 39430 58226
rect 39498 58170 39554 58226
rect 39622 58170 39678 58226
rect 39250 58046 39306 58102
rect 39374 58046 39430 58102
rect 39498 58046 39554 58102
rect 39622 58046 39678 58102
rect 39250 57922 39306 57978
rect 39374 57922 39430 57978
rect 39498 57922 39554 57978
rect 39622 57922 39678 57978
rect 39250 40294 39306 40350
rect 39374 40294 39430 40350
rect 39498 40294 39554 40350
rect 39622 40294 39678 40350
rect 39250 40170 39306 40226
rect 39374 40170 39430 40226
rect 39498 40170 39554 40226
rect 39622 40170 39678 40226
rect 39250 40046 39306 40102
rect 39374 40046 39430 40102
rect 39498 40046 39554 40102
rect 39622 40046 39678 40102
rect 39250 39922 39306 39978
rect 39374 39922 39430 39978
rect 39498 39922 39554 39978
rect 39622 39922 39678 39978
rect 39250 22294 39306 22350
rect 39374 22294 39430 22350
rect 39498 22294 39554 22350
rect 39622 22294 39678 22350
rect 39250 22170 39306 22226
rect 39374 22170 39430 22226
rect 39498 22170 39554 22226
rect 39622 22170 39678 22226
rect 39250 22046 39306 22102
rect 39374 22046 39430 22102
rect 39498 22046 39554 22102
rect 39622 22046 39678 22102
rect 39250 21922 39306 21978
rect 39374 21922 39430 21978
rect 39498 21922 39554 21978
rect 39622 21922 39678 21978
rect 39250 4294 39306 4350
rect 39374 4294 39430 4350
rect 39498 4294 39554 4350
rect 39622 4294 39678 4350
rect 39250 4170 39306 4226
rect 39374 4170 39430 4226
rect 39498 4170 39554 4226
rect 39622 4170 39678 4226
rect 39250 4046 39306 4102
rect 39374 4046 39430 4102
rect 39498 4046 39554 4102
rect 39622 4046 39678 4102
rect 39250 3922 39306 3978
rect 39374 3922 39430 3978
rect 39498 3922 39554 3978
rect 39622 3922 39678 3978
rect 39250 -216 39306 -160
rect 39374 -216 39430 -160
rect 39498 -216 39554 -160
rect 39622 -216 39678 -160
rect 39250 -340 39306 -284
rect 39374 -340 39430 -284
rect 39498 -340 39554 -284
rect 39622 -340 39678 -284
rect 39250 -464 39306 -408
rect 39374 -464 39430 -408
rect 39498 -464 39554 -408
rect 39622 -464 39678 -408
rect 39250 -588 39306 -532
rect 39374 -588 39430 -532
rect 39498 -588 39554 -532
rect 39622 -588 39678 -532
rect 57250 220294 57306 220350
rect 57374 220294 57430 220350
rect 57498 220294 57554 220350
rect 57622 220294 57678 220350
rect 57250 220170 57306 220226
rect 57374 220170 57430 220226
rect 57498 220170 57554 220226
rect 57622 220170 57678 220226
rect 57250 220046 57306 220102
rect 57374 220046 57430 220102
rect 57498 220046 57554 220102
rect 57622 220046 57678 220102
rect 57250 219922 57306 219978
rect 57374 219922 57430 219978
rect 57498 219922 57554 219978
rect 57622 219922 57678 219978
rect 60970 598116 61026 598172
rect 61094 598116 61150 598172
rect 61218 598116 61274 598172
rect 61342 598116 61398 598172
rect 60970 597992 61026 598048
rect 61094 597992 61150 598048
rect 61218 597992 61274 598048
rect 61342 597992 61398 598048
rect 60970 597868 61026 597924
rect 61094 597868 61150 597924
rect 61218 597868 61274 597924
rect 61342 597868 61398 597924
rect 60970 597744 61026 597800
rect 61094 597744 61150 597800
rect 61218 597744 61274 597800
rect 61342 597744 61398 597800
rect 78970 598116 79026 598172
rect 79094 598116 79150 598172
rect 79218 598116 79274 598172
rect 79342 598116 79398 598172
rect 78970 597992 79026 598048
rect 79094 597992 79150 598048
rect 79218 597992 79274 598048
rect 79342 597992 79398 598048
rect 78970 597868 79026 597924
rect 79094 597868 79150 597924
rect 79218 597868 79274 597924
rect 79342 597868 79398 597924
rect 78970 597744 79026 597800
rect 79094 597744 79150 597800
rect 79218 597744 79274 597800
rect 79342 597744 79398 597800
rect 60970 586294 61026 586350
rect 61094 586294 61150 586350
rect 61218 586294 61274 586350
rect 61342 586294 61398 586350
rect 60970 586170 61026 586226
rect 61094 586170 61150 586226
rect 61218 586170 61274 586226
rect 61342 586170 61398 586226
rect 60970 586046 61026 586102
rect 61094 586046 61150 586102
rect 61218 586046 61274 586102
rect 61342 586046 61398 586102
rect 60970 585922 61026 585978
rect 61094 585922 61150 585978
rect 61218 585922 61274 585978
rect 61342 585922 61398 585978
rect 60970 568294 61026 568350
rect 61094 568294 61150 568350
rect 61218 568294 61274 568350
rect 61342 568294 61398 568350
rect 60970 568170 61026 568226
rect 61094 568170 61150 568226
rect 61218 568170 61274 568226
rect 61342 568170 61398 568226
rect 60970 568046 61026 568102
rect 61094 568046 61150 568102
rect 61218 568046 61274 568102
rect 61342 568046 61398 568102
rect 60970 567922 61026 567978
rect 61094 567922 61150 567978
rect 61218 567922 61274 567978
rect 61342 567922 61398 567978
rect 60970 550294 61026 550350
rect 61094 550294 61150 550350
rect 61218 550294 61274 550350
rect 61342 550294 61398 550350
rect 60970 550170 61026 550226
rect 61094 550170 61150 550226
rect 61218 550170 61274 550226
rect 61342 550170 61398 550226
rect 60970 550046 61026 550102
rect 61094 550046 61150 550102
rect 61218 550046 61274 550102
rect 61342 550046 61398 550102
rect 60970 549922 61026 549978
rect 61094 549922 61150 549978
rect 61218 549922 61274 549978
rect 61342 549922 61398 549978
rect 60970 532294 61026 532350
rect 61094 532294 61150 532350
rect 61218 532294 61274 532350
rect 61342 532294 61398 532350
rect 60970 532170 61026 532226
rect 61094 532170 61150 532226
rect 61218 532170 61274 532226
rect 61342 532170 61398 532226
rect 60970 532046 61026 532102
rect 61094 532046 61150 532102
rect 61218 532046 61274 532102
rect 61342 532046 61398 532102
rect 60970 531922 61026 531978
rect 61094 531922 61150 531978
rect 61218 531922 61274 531978
rect 61342 531922 61398 531978
rect 60970 514294 61026 514350
rect 61094 514294 61150 514350
rect 61218 514294 61274 514350
rect 61342 514294 61398 514350
rect 60970 514170 61026 514226
rect 61094 514170 61150 514226
rect 61218 514170 61274 514226
rect 61342 514170 61398 514226
rect 60970 514046 61026 514102
rect 61094 514046 61150 514102
rect 61218 514046 61274 514102
rect 61342 514046 61398 514102
rect 60970 513922 61026 513978
rect 61094 513922 61150 513978
rect 61218 513922 61274 513978
rect 61342 513922 61398 513978
rect 60970 496294 61026 496350
rect 61094 496294 61150 496350
rect 61218 496294 61274 496350
rect 61342 496294 61398 496350
rect 60970 496170 61026 496226
rect 61094 496170 61150 496226
rect 61218 496170 61274 496226
rect 61342 496170 61398 496226
rect 60970 496046 61026 496102
rect 61094 496046 61150 496102
rect 61218 496046 61274 496102
rect 61342 496046 61398 496102
rect 60970 495922 61026 495978
rect 61094 495922 61150 495978
rect 61218 495922 61274 495978
rect 61342 495922 61398 495978
rect 60970 478294 61026 478350
rect 61094 478294 61150 478350
rect 61218 478294 61274 478350
rect 61342 478294 61398 478350
rect 60970 478170 61026 478226
rect 61094 478170 61150 478226
rect 61218 478170 61274 478226
rect 61342 478170 61398 478226
rect 60970 478046 61026 478102
rect 61094 478046 61150 478102
rect 61218 478046 61274 478102
rect 61342 478046 61398 478102
rect 60970 477922 61026 477978
rect 61094 477922 61150 477978
rect 61218 477922 61274 477978
rect 61342 477922 61398 477978
rect 60970 460294 61026 460350
rect 61094 460294 61150 460350
rect 61218 460294 61274 460350
rect 61342 460294 61398 460350
rect 60970 460170 61026 460226
rect 61094 460170 61150 460226
rect 61218 460170 61274 460226
rect 61342 460170 61398 460226
rect 60970 460046 61026 460102
rect 61094 460046 61150 460102
rect 61218 460046 61274 460102
rect 61342 460046 61398 460102
rect 60970 459922 61026 459978
rect 61094 459922 61150 459978
rect 61218 459922 61274 459978
rect 61342 459922 61398 459978
rect 60970 442294 61026 442350
rect 61094 442294 61150 442350
rect 61218 442294 61274 442350
rect 61342 442294 61398 442350
rect 60970 442170 61026 442226
rect 61094 442170 61150 442226
rect 61218 442170 61274 442226
rect 61342 442170 61398 442226
rect 60970 442046 61026 442102
rect 61094 442046 61150 442102
rect 61218 442046 61274 442102
rect 61342 442046 61398 442102
rect 60970 441922 61026 441978
rect 61094 441922 61150 441978
rect 61218 441922 61274 441978
rect 61342 441922 61398 441978
rect 60970 424294 61026 424350
rect 61094 424294 61150 424350
rect 61218 424294 61274 424350
rect 61342 424294 61398 424350
rect 60970 424170 61026 424226
rect 61094 424170 61150 424226
rect 61218 424170 61274 424226
rect 61342 424170 61398 424226
rect 60970 424046 61026 424102
rect 61094 424046 61150 424102
rect 61218 424046 61274 424102
rect 61342 424046 61398 424102
rect 60970 423922 61026 423978
rect 61094 423922 61150 423978
rect 61218 423922 61274 423978
rect 61342 423922 61398 423978
rect 60970 406294 61026 406350
rect 61094 406294 61150 406350
rect 61218 406294 61274 406350
rect 61342 406294 61398 406350
rect 60970 406170 61026 406226
rect 61094 406170 61150 406226
rect 61218 406170 61274 406226
rect 61342 406170 61398 406226
rect 60970 406046 61026 406102
rect 61094 406046 61150 406102
rect 61218 406046 61274 406102
rect 61342 406046 61398 406102
rect 60970 405922 61026 405978
rect 61094 405922 61150 405978
rect 61218 405922 61274 405978
rect 61342 405922 61398 405978
rect 60970 388294 61026 388350
rect 61094 388294 61150 388350
rect 61218 388294 61274 388350
rect 61342 388294 61398 388350
rect 60970 388170 61026 388226
rect 61094 388170 61150 388226
rect 61218 388170 61274 388226
rect 61342 388170 61398 388226
rect 60970 388046 61026 388102
rect 61094 388046 61150 388102
rect 61218 388046 61274 388102
rect 61342 388046 61398 388102
rect 60970 387922 61026 387978
rect 61094 387922 61150 387978
rect 61218 387922 61274 387978
rect 61342 387922 61398 387978
rect 60970 370294 61026 370350
rect 61094 370294 61150 370350
rect 61218 370294 61274 370350
rect 61342 370294 61398 370350
rect 60970 370170 61026 370226
rect 61094 370170 61150 370226
rect 61218 370170 61274 370226
rect 61342 370170 61398 370226
rect 60970 370046 61026 370102
rect 61094 370046 61150 370102
rect 61218 370046 61274 370102
rect 61342 370046 61398 370102
rect 60970 369922 61026 369978
rect 61094 369922 61150 369978
rect 61218 369922 61274 369978
rect 61342 369922 61398 369978
rect 60970 352294 61026 352350
rect 61094 352294 61150 352350
rect 61218 352294 61274 352350
rect 61342 352294 61398 352350
rect 60970 352170 61026 352226
rect 61094 352170 61150 352226
rect 61218 352170 61274 352226
rect 61342 352170 61398 352226
rect 60970 352046 61026 352102
rect 61094 352046 61150 352102
rect 61218 352046 61274 352102
rect 61342 352046 61398 352102
rect 60970 351922 61026 351978
rect 61094 351922 61150 351978
rect 61218 351922 61274 351978
rect 61342 351922 61398 351978
rect 60970 334294 61026 334350
rect 61094 334294 61150 334350
rect 61218 334294 61274 334350
rect 61342 334294 61398 334350
rect 60970 334170 61026 334226
rect 61094 334170 61150 334226
rect 61218 334170 61274 334226
rect 61342 334170 61398 334226
rect 60970 334046 61026 334102
rect 61094 334046 61150 334102
rect 61218 334046 61274 334102
rect 61342 334046 61398 334102
rect 60970 333922 61026 333978
rect 61094 333922 61150 333978
rect 61218 333922 61274 333978
rect 61342 333922 61398 333978
rect 60970 316294 61026 316350
rect 61094 316294 61150 316350
rect 61218 316294 61274 316350
rect 61342 316294 61398 316350
rect 60970 316170 61026 316226
rect 61094 316170 61150 316226
rect 61218 316170 61274 316226
rect 61342 316170 61398 316226
rect 60970 316046 61026 316102
rect 61094 316046 61150 316102
rect 61218 316046 61274 316102
rect 61342 316046 61398 316102
rect 60970 315922 61026 315978
rect 61094 315922 61150 315978
rect 61218 315922 61274 315978
rect 61342 315922 61398 315978
rect 60970 298294 61026 298350
rect 61094 298294 61150 298350
rect 61218 298294 61274 298350
rect 61342 298294 61398 298350
rect 60970 298170 61026 298226
rect 61094 298170 61150 298226
rect 61218 298170 61274 298226
rect 61342 298170 61398 298226
rect 60970 298046 61026 298102
rect 61094 298046 61150 298102
rect 61218 298046 61274 298102
rect 61342 298046 61398 298102
rect 60970 297922 61026 297978
rect 61094 297922 61150 297978
rect 61218 297922 61274 297978
rect 61342 297922 61398 297978
rect 60970 280294 61026 280350
rect 61094 280294 61150 280350
rect 61218 280294 61274 280350
rect 61342 280294 61398 280350
rect 60970 280170 61026 280226
rect 61094 280170 61150 280226
rect 61218 280170 61274 280226
rect 61342 280170 61398 280226
rect 60970 280046 61026 280102
rect 61094 280046 61150 280102
rect 61218 280046 61274 280102
rect 61342 280046 61398 280102
rect 60970 279922 61026 279978
rect 61094 279922 61150 279978
rect 61218 279922 61274 279978
rect 61342 279922 61398 279978
rect 60970 262294 61026 262350
rect 61094 262294 61150 262350
rect 61218 262294 61274 262350
rect 61342 262294 61398 262350
rect 60970 262170 61026 262226
rect 61094 262170 61150 262226
rect 61218 262170 61274 262226
rect 61342 262170 61398 262226
rect 60970 262046 61026 262102
rect 61094 262046 61150 262102
rect 61218 262046 61274 262102
rect 61342 262046 61398 262102
rect 60970 261922 61026 261978
rect 61094 261922 61150 261978
rect 61218 261922 61274 261978
rect 61342 261922 61398 261978
rect 60970 244294 61026 244350
rect 61094 244294 61150 244350
rect 61218 244294 61274 244350
rect 61342 244294 61398 244350
rect 60970 244170 61026 244226
rect 61094 244170 61150 244226
rect 61218 244170 61274 244226
rect 61342 244170 61398 244226
rect 60970 244046 61026 244102
rect 61094 244046 61150 244102
rect 61218 244046 61274 244102
rect 61342 244046 61398 244102
rect 60970 243922 61026 243978
rect 61094 243922 61150 243978
rect 61218 243922 61274 243978
rect 61342 243922 61398 243978
rect 78970 586294 79026 586350
rect 79094 586294 79150 586350
rect 79218 586294 79274 586350
rect 79342 586294 79398 586350
rect 78970 586170 79026 586226
rect 79094 586170 79150 586226
rect 79218 586170 79274 586226
rect 79342 586170 79398 586226
rect 78970 586046 79026 586102
rect 79094 586046 79150 586102
rect 79218 586046 79274 586102
rect 79342 586046 79398 586102
rect 78970 585922 79026 585978
rect 79094 585922 79150 585978
rect 79218 585922 79274 585978
rect 79342 585922 79398 585978
rect 78970 568294 79026 568350
rect 79094 568294 79150 568350
rect 79218 568294 79274 568350
rect 79342 568294 79398 568350
rect 78970 568170 79026 568226
rect 79094 568170 79150 568226
rect 79218 568170 79274 568226
rect 79342 568170 79398 568226
rect 78970 568046 79026 568102
rect 79094 568046 79150 568102
rect 79218 568046 79274 568102
rect 79342 568046 79398 568102
rect 78970 567922 79026 567978
rect 79094 567922 79150 567978
rect 79218 567922 79274 567978
rect 79342 567922 79398 567978
rect 78970 550294 79026 550350
rect 79094 550294 79150 550350
rect 79218 550294 79274 550350
rect 79342 550294 79398 550350
rect 78970 550170 79026 550226
rect 79094 550170 79150 550226
rect 79218 550170 79274 550226
rect 79342 550170 79398 550226
rect 78970 550046 79026 550102
rect 79094 550046 79150 550102
rect 79218 550046 79274 550102
rect 79342 550046 79398 550102
rect 78970 549922 79026 549978
rect 79094 549922 79150 549978
rect 79218 549922 79274 549978
rect 79342 549922 79398 549978
rect 78970 532294 79026 532350
rect 79094 532294 79150 532350
rect 79218 532294 79274 532350
rect 79342 532294 79398 532350
rect 78970 532170 79026 532226
rect 79094 532170 79150 532226
rect 79218 532170 79274 532226
rect 79342 532170 79398 532226
rect 78970 532046 79026 532102
rect 79094 532046 79150 532102
rect 79218 532046 79274 532102
rect 79342 532046 79398 532102
rect 78970 531922 79026 531978
rect 79094 531922 79150 531978
rect 79218 531922 79274 531978
rect 79342 531922 79398 531978
rect 78970 514294 79026 514350
rect 79094 514294 79150 514350
rect 79218 514294 79274 514350
rect 79342 514294 79398 514350
rect 78970 514170 79026 514226
rect 79094 514170 79150 514226
rect 79218 514170 79274 514226
rect 79342 514170 79398 514226
rect 78970 514046 79026 514102
rect 79094 514046 79150 514102
rect 79218 514046 79274 514102
rect 79342 514046 79398 514102
rect 78970 513922 79026 513978
rect 79094 513922 79150 513978
rect 79218 513922 79274 513978
rect 79342 513922 79398 513978
rect 78970 496294 79026 496350
rect 79094 496294 79150 496350
rect 79218 496294 79274 496350
rect 79342 496294 79398 496350
rect 78970 496170 79026 496226
rect 79094 496170 79150 496226
rect 79218 496170 79274 496226
rect 79342 496170 79398 496226
rect 78970 496046 79026 496102
rect 79094 496046 79150 496102
rect 79218 496046 79274 496102
rect 79342 496046 79398 496102
rect 78970 495922 79026 495978
rect 79094 495922 79150 495978
rect 79218 495922 79274 495978
rect 79342 495922 79398 495978
rect 78970 478294 79026 478350
rect 79094 478294 79150 478350
rect 79218 478294 79274 478350
rect 79342 478294 79398 478350
rect 78970 478170 79026 478226
rect 79094 478170 79150 478226
rect 79218 478170 79274 478226
rect 79342 478170 79398 478226
rect 78970 478046 79026 478102
rect 79094 478046 79150 478102
rect 79218 478046 79274 478102
rect 79342 478046 79398 478102
rect 78970 477922 79026 477978
rect 79094 477922 79150 477978
rect 79218 477922 79274 477978
rect 79342 477922 79398 477978
rect 78970 460294 79026 460350
rect 79094 460294 79150 460350
rect 79218 460294 79274 460350
rect 79342 460294 79398 460350
rect 78970 460170 79026 460226
rect 79094 460170 79150 460226
rect 79218 460170 79274 460226
rect 79342 460170 79398 460226
rect 78970 460046 79026 460102
rect 79094 460046 79150 460102
rect 79218 460046 79274 460102
rect 79342 460046 79398 460102
rect 78970 459922 79026 459978
rect 79094 459922 79150 459978
rect 79218 459922 79274 459978
rect 79342 459922 79398 459978
rect 78970 442294 79026 442350
rect 79094 442294 79150 442350
rect 79218 442294 79274 442350
rect 79342 442294 79398 442350
rect 78970 442170 79026 442226
rect 79094 442170 79150 442226
rect 79218 442170 79274 442226
rect 79342 442170 79398 442226
rect 78970 442046 79026 442102
rect 79094 442046 79150 442102
rect 79218 442046 79274 442102
rect 79342 442046 79398 442102
rect 78970 441922 79026 441978
rect 79094 441922 79150 441978
rect 79218 441922 79274 441978
rect 79342 441922 79398 441978
rect 78970 424294 79026 424350
rect 79094 424294 79150 424350
rect 79218 424294 79274 424350
rect 79342 424294 79398 424350
rect 78970 424170 79026 424226
rect 79094 424170 79150 424226
rect 79218 424170 79274 424226
rect 79342 424170 79398 424226
rect 78970 424046 79026 424102
rect 79094 424046 79150 424102
rect 79218 424046 79274 424102
rect 79342 424046 79398 424102
rect 78970 423922 79026 423978
rect 79094 423922 79150 423978
rect 79218 423922 79274 423978
rect 79342 423922 79398 423978
rect 78970 406294 79026 406350
rect 79094 406294 79150 406350
rect 79218 406294 79274 406350
rect 79342 406294 79398 406350
rect 78970 406170 79026 406226
rect 79094 406170 79150 406226
rect 79218 406170 79274 406226
rect 79342 406170 79398 406226
rect 78970 406046 79026 406102
rect 79094 406046 79150 406102
rect 79218 406046 79274 406102
rect 79342 406046 79398 406102
rect 78970 405922 79026 405978
rect 79094 405922 79150 405978
rect 79218 405922 79274 405978
rect 79342 405922 79398 405978
rect 78970 388294 79026 388350
rect 79094 388294 79150 388350
rect 79218 388294 79274 388350
rect 79342 388294 79398 388350
rect 78970 388170 79026 388226
rect 79094 388170 79150 388226
rect 79218 388170 79274 388226
rect 79342 388170 79398 388226
rect 78970 388046 79026 388102
rect 79094 388046 79150 388102
rect 79218 388046 79274 388102
rect 79342 388046 79398 388102
rect 78970 387922 79026 387978
rect 79094 387922 79150 387978
rect 79218 387922 79274 387978
rect 79342 387922 79398 387978
rect 78970 370294 79026 370350
rect 79094 370294 79150 370350
rect 79218 370294 79274 370350
rect 79342 370294 79398 370350
rect 78970 370170 79026 370226
rect 79094 370170 79150 370226
rect 79218 370170 79274 370226
rect 79342 370170 79398 370226
rect 78970 370046 79026 370102
rect 79094 370046 79150 370102
rect 79218 370046 79274 370102
rect 79342 370046 79398 370102
rect 78970 369922 79026 369978
rect 79094 369922 79150 369978
rect 79218 369922 79274 369978
rect 79342 369922 79398 369978
rect 78970 352294 79026 352350
rect 79094 352294 79150 352350
rect 79218 352294 79274 352350
rect 79342 352294 79398 352350
rect 78970 352170 79026 352226
rect 79094 352170 79150 352226
rect 79218 352170 79274 352226
rect 79342 352170 79398 352226
rect 78970 352046 79026 352102
rect 79094 352046 79150 352102
rect 79218 352046 79274 352102
rect 79342 352046 79398 352102
rect 78970 351922 79026 351978
rect 79094 351922 79150 351978
rect 79218 351922 79274 351978
rect 79342 351922 79398 351978
rect 78970 334294 79026 334350
rect 79094 334294 79150 334350
rect 79218 334294 79274 334350
rect 79342 334294 79398 334350
rect 78970 334170 79026 334226
rect 79094 334170 79150 334226
rect 79218 334170 79274 334226
rect 79342 334170 79398 334226
rect 78970 334046 79026 334102
rect 79094 334046 79150 334102
rect 79218 334046 79274 334102
rect 79342 334046 79398 334102
rect 78970 333922 79026 333978
rect 79094 333922 79150 333978
rect 79218 333922 79274 333978
rect 79342 333922 79398 333978
rect 78970 316294 79026 316350
rect 79094 316294 79150 316350
rect 79218 316294 79274 316350
rect 79342 316294 79398 316350
rect 78970 316170 79026 316226
rect 79094 316170 79150 316226
rect 79218 316170 79274 316226
rect 79342 316170 79398 316226
rect 78970 316046 79026 316102
rect 79094 316046 79150 316102
rect 79218 316046 79274 316102
rect 79342 316046 79398 316102
rect 78970 315922 79026 315978
rect 79094 315922 79150 315978
rect 79218 315922 79274 315978
rect 79342 315922 79398 315978
rect 78970 298294 79026 298350
rect 79094 298294 79150 298350
rect 79218 298294 79274 298350
rect 79342 298294 79398 298350
rect 78970 298170 79026 298226
rect 79094 298170 79150 298226
rect 79218 298170 79274 298226
rect 79342 298170 79398 298226
rect 78970 298046 79026 298102
rect 79094 298046 79150 298102
rect 79218 298046 79274 298102
rect 79342 298046 79398 298102
rect 78970 297922 79026 297978
rect 79094 297922 79150 297978
rect 79218 297922 79274 297978
rect 79342 297922 79398 297978
rect 78970 280294 79026 280350
rect 79094 280294 79150 280350
rect 79218 280294 79274 280350
rect 79342 280294 79398 280350
rect 78970 280170 79026 280226
rect 79094 280170 79150 280226
rect 79218 280170 79274 280226
rect 79342 280170 79398 280226
rect 78970 280046 79026 280102
rect 79094 280046 79150 280102
rect 79218 280046 79274 280102
rect 79342 280046 79398 280102
rect 78970 279922 79026 279978
rect 79094 279922 79150 279978
rect 79218 279922 79274 279978
rect 79342 279922 79398 279978
rect 78970 262294 79026 262350
rect 79094 262294 79150 262350
rect 79218 262294 79274 262350
rect 79342 262294 79398 262350
rect 78970 262170 79026 262226
rect 79094 262170 79150 262226
rect 79218 262170 79274 262226
rect 79342 262170 79398 262226
rect 78970 262046 79026 262102
rect 79094 262046 79150 262102
rect 79218 262046 79274 262102
rect 79342 262046 79398 262102
rect 78970 261922 79026 261978
rect 79094 261922 79150 261978
rect 79218 261922 79274 261978
rect 79342 261922 79398 261978
rect 78970 244294 79026 244350
rect 79094 244294 79150 244350
rect 79218 244294 79274 244350
rect 79342 244294 79398 244350
rect 78970 244170 79026 244226
rect 79094 244170 79150 244226
rect 79218 244170 79274 244226
rect 79342 244170 79398 244226
rect 78970 244046 79026 244102
rect 79094 244046 79150 244102
rect 79218 244046 79274 244102
rect 79342 244046 79398 244102
rect 78970 243922 79026 243978
rect 79094 243922 79150 243978
rect 79218 243922 79274 243978
rect 79342 243922 79398 243978
rect 75250 238294 75306 238350
rect 75374 238294 75430 238350
rect 75498 238294 75554 238350
rect 75622 238294 75678 238350
rect 75250 238170 75306 238226
rect 75374 238170 75430 238226
rect 75498 238170 75554 238226
rect 75622 238170 75678 238226
rect 75250 238046 75306 238102
rect 75374 238046 75430 238102
rect 75498 238046 75554 238102
rect 75622 238046 75678 238102
rect 75250 237922 75306 237978
rect 75374 237922 75430 237978
rect 75498 237922 75554 237978
rect 75622 237922 75678 237978
rect 60970 226294 61026 226350
rect 61094 226294 61150 226350
rect 61218 226294 61274 226350
rect 61342 226294 61398 226350
rect 60970 226170 61026 226226
rect 61094 226170 61150 226226
rect 61218 226170 61274 226226
rect 61342 226170 61398 226226
rect 60970 226046 61026 226102
rect 61094 226046 61150 226102
rect 61218 226046 61274 226102
rect 61342 226046 61398 226102
rect 60970 225922 61026 225978
rect 61094 225922 61150 225978
rect 61218 225922 61274 225978
rect 61342 225922 61398 225978
rect 64518 220294 64574 220350
rect 64642 220294 64698 220350
rect 64518 220170 64574 220226
rect 64642 220170 64698 220226
rect 64518 220046 64574 220102
rect 64642 220046 64698 220102
rect 64518 219922 64574 219978
rect 64642 219922 64698 219978
rect 75250 220294 75306 220350
rect 75374 220294 75430 220350
rect 75498 220294 75554 220350
rect 75622 220294 75678 220350
rect 75250 220170 75306 220226
rect 75374 220170 75430 220226
rect 75498 220170 75554 220226
rect 75622 220170 75678 220226
rect 75250 220046 75306 220102
rect 75374 220046 75430 220102
rect 75498 220046 75554 220102
rect 75622 220046 75678 220102
rect 75250 219922 75306 219978
rect 75374 219922 75430 219978
rect 75498 219922 75554 219978
rect 75622 219922 75678 219978
rect 93250 597156 93306 597212
rect 93374 597156 93430 597212
rect 93498 597156 93554 597212
rect 93622 597156 93678 597212
rect 93250 597032 93306 597088
rect 93374 597032 93430 597088
rect 93498 597032 93554 597088
rect 93622 597032 93678 597088
rect 93250 596908 93306 596964
rect 93374 596908 93430 596964
rect 93498 596908 93554 596964
rect 93622 596908 93678 596964
rect 93250 596784 93306 596840
rect 93374 596784 93430 596840
rect 93498 596784 93554 596840
rect 93622 596784 93678 596840
rect 93250 580294 93306 580350
rect 93374 580294 93430 580350
rect 93498 580294 93554 580350
rect 93622 580294 93678 580350
rect 93250 580170 93306 580226
rect 93374 580170 93430 580226
rect 93498 580170 93554 580226
rect 93622 580170 93678 580226
rect 93250 580046 93306 580102
rect 93374 580046 93430 580102
rect 93498 580046 93554 580102
rect 93622 580046 93678 580102
rect 93250 579922 93306 579978
rect 93374 579922 93430 579978
rect 93498 579922 93554 579978
rect 93622 579922 93678 579978
rect 93250 562294 93306 562350
rect 93374 562294 93430 562350
rect 93498 562294 93554 562350
rect 93622 562294 93678 562350
rect 93250 562170 93306 562226
rect 93374 562170 93430 562226
rect 93498 562170 93554 562226
rect 93622 562170 93678 562226
rect 93250 562046 93306 562102
rect 93374 562046 93430 562102
rect 93498 562046 93554 562102
rect 93622 562046 93678 562102
rect 93250 561922 93306 561978
rect 93374 561922 93430 561978
rect 93498 561922 93554 561978
rect 93622 561922 93678 561978
rect 93250 544294 93306 544350
rect 93374 544294 93430 544350
rect 93498 544294 93554 544350
rect 93622 544294 93678 544350
rect 93250 544170 93306 544226
rect 93374 544170 93430 544226
rect 93498 544170 93554 544226
rect 93622 544170 93678 544226
rect 93250 544046 93306 544102
rect 93374 544046 93430 544102
rect 93498 544046 93554 544102
rect 93622 544046 93678 544102
rect 93250 543922 93306 543978
rect 93374 543922 93430 543978
rect 93498 543922 93554 543978
rect 93622 543922 93678 543978
rect 93250 526294 93306 526350
rect 93374 526294 93430 526350
rect 93498 526294 93554 526350
rect 93622 526294 93678 526350
rect 93250 526170 93306 526226
rect 93374 526170 93430 526226
rect 93498 526170 93554 526226
rect 93622 526170 93678 526226
rect 93250 526046 93306 526102
rect 93374 526046 93430 526102
rect 93498 526046 93554 526102
rect 93622 526046 93678 526102
rect 93250 525922 93306 525978
rect 93374 525922 93430 525978
rect 93498 525922 93554 525978
rect 93622 525922 93678 525978
rect 93250 508294 93306 508350
rect 93374 508294 93430 508350
rect 93498 508294 93554 508350
rect 93622 508294 93678 508350
rect 93250 508170 93306 508226
rect 93374 508170 93430 508226
rect 93498 508170 93554 508226
rect 93622 508170 93678 508226
rect 93250 508046 93306 508102
rect 93374 508046 93430 508102
rect 93498 508046 93554 508102
rect 93622 508046 93678 508102
rect 93250 507922 93306 507978
rect 93374 507922 93430 507978
rect 93498 507922 93554 507978
rect 93622 507922 93678 507978
rect 93250 490294 93306 490350
rect 93374 490294 93430 490350
rect 93498 490294 93554 490350
rect 93622 490294 93678 490350
rect 93250 490170 93306 490226
rect 93374 490170 93430 490226
rect 93498 490170 93554 490226
rect 93622 490170 93678 490226
rect 93250 490046 93306 490102
rect 93374 490046 93430 490102
rect 93498 490046 93554 490102
rect 93622 490046 93678 490102
rect 93250 489922 93306 489978
rect 93374 489922 93430 489978
rect 93498 489922 93554 489978
rect 93622 489922 93678 489978
rect 93250 472294 93306 472350
rect 93374 472294 93430 472350
rect 93498 472294 93554 472350
rect 93622 472294 93678 472350
rect 93250 472170 93306 472226
rect 93374 472170 93430 472226
rect 93498 472170 93554 472226
rect 93622 472170 93678 472226
rect 93250 472046 93306 472102
rect 93374 472046 93430 472102
rect 93498 472046 93554 472102
rect 93622 472046 93678 472102
rect 93250 471922 93306 471978
rect 93374 471922 93430 471978
rect 93498 471922 93554 471978
rect 93622 471922 93678 471978
rect 93250 454294 93306 454350
rect 93374 454294 93430 454350
rect 93498 454294 93554 454350
rect 93622 454294 93678 454350
rect 93250 454170 93306 454226
rect 93374 454170 93430 454226
rect 93498 454170 93554 454226
rect 93622 454170 93678 454226
rect 93250 454046 93306 454102
rect 93374 454046 93430 454102
rect 93498 454046 93554 454102
rect 93622 454046 93678 454102
rect 93250 453922 93306 453978
rect 93374 453922 93430 453978
rect 93498 453922 93554 453978
rect 93622 453922 93678 453978
rect 93250 436294 93306 436350
rect 93374 436294 93430 436350
rect 93498 436294 93554 436350
rect 93622 436294 93678 436350
rect 93250 436170 93306 436226
rect 93374 436170 93430 436226
rect 93498 436170 93554 436226
rect 93622 436170 93678 436226
rect 93250 436046 93306 436102
rect 93374 436046 93430 436102
rect 93498 436046 93554 436102
rect 93622 436046 93678 436102
rect 93250 435922 93306 435978
rect 93374 435922 93430 435978
rect 93498 435922 93554 435978
rect 93622 435922 93678 435978
rect 93250 418294 93306 418350
rect 93374 418294 93430 418350
rect 93498 418294 93554 418350
rect 93622 418294 93678 418350
rect 93250 418170 93306 418226
rect 93374 418170 93430 418226
rect 93498 418170 93554 418226
rect 93622 418170 93678 418226
rect 93250 418046 93306 418102
rect 93374 418046 93430 418102
rect 93498 418046 93554 418102
rect 93622 418046 93678 418102
rect 93250 417922 93306 417978
rect 93374 417922 93430 417978
rect 93498 417922 93554 417978
rect 93622 417922 93678 417978
rect 93250 400294 93306 400350
rect 93374 400294 93430 400350
rect 93498 400294 93554 400350
rect 93622 400294 93678 400350
rect 93250 400170 93306 400226
rect 93374 400170 93430 400226
rect 93498 400170 93554 400226
rect 93622 400170 93678 400226
rect 93250 400046 93306 400102
rect 93374 400046 93430 400102
rect 93498 400046 93554 400102
rect 93622 400046 93678 400102
rect 93250 399922 93306 399978
rect 93374 399922 93430 399978
rect 93498 399922 93554 399978
rect 93622 399922 93678 399978
rect 93250 382294 93306 382350
rect 93374 382294 93430 382350
rect 93498 382294 93554 382350
rect 93622 382294 93678 382350
rect 93250 382170 93306 382226
rect 93374 382170 93430 382226
rect 93498 382170 93554 382226
rect 93622 382170 93678 382226
rect 93250 382046 93306 382102
rect 93374 382046 93430 382102
rect 93498 382046 93554 382102
rect 93622 382046 93678 382102
rect 93250 381922 93306 381978
rect 93374 381922 93430 381978
rect 93498 381922 93554 381978
rect 93622 381922 93678 381978
rect 93250 364294 93306 364350
rect 93374 364294 93430 364350
rect 93498 364294 93554 364350
rect 93622 364294 93678 364350
rect 93250 364170 93306 364226
rect 93374 364170 93430 364226
rect 93498 364170 93554 364226
rect 93622 364170 93678 364226
rect 93250 364046 93306 364102
rect 93374 364046 93430 364102
rect 93498 364046 93554 364102
rect 93622 364046 93678 364102
rect 93250 363922 93306 363978
rect 93374 363922 93430 363978
rect 93498 363922 93554 363978
rect 93622 363922 93678 363978
rect 93250 346294 93306 346350
rect 93374 346294 93430 346350
rect 93498 346294 93554 346350
rect 93622 346294 93678 346350
rect 93250 346170 93306 346226
rect 93374 346170 93430 346226
rect 93498 346170 93554 346226
rect 93622 346170 93678 346226
rect 93250 346046 93306 346102
rect 93374 346046 93430 346102
rect 93498 346046 93554 346102
rect 93622 346046 93678 346102
rect 93250 345922 93306 345978
rect 93374 345922 93430 345978
rect 93498 345922 93554 345978
rect 93622 345922 93678 345978
rect 93250 328294 93306 328350
rect 93374 328294 93430 328350
rect 93498 328294 93554 328350
rect 93622 328294 93678 328350
rect 93250 328170 93306 328226
rect 93374 328170 93430 328226
rect 93498 328170 93554 328226
rect 93622 328170 93678 328226
rect 93250 328046 93306 328102
rect 93374 328046 93430 328102
rect 93498 328046 93554 328102
rect 93622 328046 93678 328102
rect 93250 327922 93306 327978
rect 93374 327922 93430 327978
rect 93498 327922 93554 327978
rect 93622 327922 93678 327978
rect 93250 310294 93306 310350
rect 93374 310294 93430 310350
rect 93498 310294 93554 310350
rect 93622 310294 93678 310350
rect 93250 310170 93306 310226
rect 93374 310170 93430 310226
rect 93498 310170 93554 310226
rect 93622 310170 93678 310226
rect 93250 310046 93306 310102
rect 93374 310046 93430 310102
rect 93498 310046 93554 310102
rect 93622 310046 93678 310102
rect 93250 309922 93306 309978
rect 93374 309922 93430 309978
rect 93498 309922 93554 309978
rect 93622 309922 93678 309978
rect 93250 292294 93306 292350
rect 93374 292294 93430 292350
rect 93498 292294 93554 292350
rect 93622 292294 93678 292350
rect 93250 292170 93306 292226
rect 93374 292170 93430 292226
rect 93498 292170 93554 292226
rect 93622 292170 93678 292226
rect 93250 292046 93306 292102
rect 93374 292046 93430 292102
rect 93498 292046 93554 292102
rect 93622 292046 93678 292102
rect 93250 291922 93306 291978
rect 93374 291922 93430 291978
rect 93498 291922 93554 291978
rect 93622 291922 93678 291978
rect 93250 274294 93306 274350
rect 93374 274294 93430 274350
rect 93498 274294 93554 274350
rect 93622 274294 93678 274350
rect 93250 274170 93306 274226
rect 93374 274170 93430 274226
rect 93498 274170 93554 274226
rect 93622 274170 93678 274226
rect 93250 274046 93306 274102
rect 93374 274046 93430 274102
rect 93498 274046 93554 274102
rect 93622 274046 93678 274102
rect 93250 273922 93306 273978
rect 93374 273922 93430 273978
rect 93498 273922 93554 273978
rect 93622 273922 93678 273978
rect 93250 256294 93306 256350
rect 93374 256294 93430 256350
rect 93498 256294 93554 256350
rect 93622 256294 93678 256350
rect 93250 256170 93306 256226
rect 93374 256170 93430 256226
rect 93498 256170 93554 256226
rect 93622 256170 93678 256226
rect 93250 256046 93306 256102
rect 93374 256046 93430 256102
rect 93498 256046 93554 256102
rect 93622 256046 93678 256102
rect 93250 255922 93306 255978
rect 93374 255922 93430 255978
rect 93498 255922 93554 255978
rect 93622 255922 93678 255978
rect 93250 238294 93306 238350
rect 93374 238294 93430 238350
rect 93498 238294 93554 238350
rect 93622 238294 93678 238350
rect 93250 238170 93306 238226
rect 93374 238170 93430 238226
rect 93498 238170 93554 238226
rect 93622 238170 93678 238226
rect 93250 238046 93306 238102
rect 93374 238046 93430 238102
rect 93498 238046 93554 238102
rect 93622 238046 93678 238102
rect 93250 237922 93306 237978
rect 93374 237922 93430 237978
rect 93498 237922 93554 237978
rect 93622 237922 93678 237978
rect 78970 226294 79026 226350
rect 79094 226294 79150 226350
rect 79218 226294 79274 226350
rect 79342 226294 79398 226350
rect 78970 226170 79026 226226
rect 79094 226170 79150 226226
rect 79218 226170 79274 226226
rect 79342 226170 79398 226226
rect 78970 226046 79026 226102
rect 79094 226046 79150 226102
rect 79218 226046 79274 226102
rect 79342 226046 79398 226102
rect 78970 225922 79026 225978
rect 79094 225922 79150 225978
rect 79218 225922 79274 225978
rect 79342 225922 79398 225978
rect 79878 226294 79934 226350
rect 80002 226294 80058 226350
rect 79878 226170 79934 226226
rect 80002 226170 80058 226226
rect 79878 226046 79934 226102
rect 80002 226046 80058 226102
rect 79878 225922 79934 225978
rect 80002 225922 80058 225978
rect 96970 598116 97026 598172
rect 97094 598116 97150 598172
rect 97218 598116 97274 598172
rect 97342 598116 97398 598172
rect 96970 597992 97026 598048
rect 97094 597992 97150 598048
rect 97218 597992 97274 598048
rect 97342 597992 97398 598048
rect 96970 597868 97026 597924
rect 97094 597868 97150 597924
rect 97218 597868 97274 597924
rect 97342 597868 97398 597924
rect 96970 597744 97026 597800
rect 97094 597744 97150 597800
rect 97218 597744 97274 597800
rect 97342 597744 97398 597800
rect 96970 586294 97026 586350
rect 97094 586294 97150 586350
rect 97218 586294 97274 586350
rect 97342 586294 97398 586350
rect 96970 586170 97026 586226
rect 97094 586170 97150 586226
rect 97218 586170 97274 586226
rect 97342 586170 97398 586226
rect 96970 586046 97026 586102
rect 97094 586046 97150 586102
rect 97218 586046 97274 586102
rect 97342 586046 97398 586102
rect 96970 585922 97026 585978
rect 97094 585922 97150 585978
rect 97218 585922 97274 585978
rect 97342 585922 97398 585978
rect 96970 568294 97026 568350
rect 97094 568294 97150 568350
rect 97218 568294 97274 568350
rect 97342 568294 97398 568350
rect 96970 568170 97026 568226
rect 97094 568170 97150 568226
rect 97218 568170 97274 568226
rect 97342 568170 97398 568226
rect 96970 568046 97026 568102
rect 97094 568046 97150 568102
rect 97218 568046 97274 568102
rect 97342 568046 97398 568102
rect 96970 567922 97026 567978
rect 97094 567922 97150 567978
rect 97218 567922 97274 567978
rect 97342 567922 97398 567978
rect 96970 550294 97026 550350
rect 97094 550294 97150 550350
rect 97218 550294 97274 550350
rect 97342 550294 97398 550350
rect 96970 550170 97026 550226
rect 97094 550170 97150 550226
rect 97218 550170 97274 550226
rect 97342 550170 97398 550226
rect 96970 550046 97026 550102
rect 97094 550046 97150 550102
rect 97218 550046 97274 550102
rect 97342 550046 97398 550102
rect 96970 549922 97026 549978
rect 97094 549922 97150 549978
rect 97218 549922 97274 549978
rect 97342 549922 97398 549978
rect 96970 532294 97026 532350
rect 97094 532294 97150 532350
rect 97218 532294 97274 532350
rect 97342 532294 97398 532350
rect 96970 532170 97026 532226
rect 97094 532170 97150 532226
rect 97218 532170 97274 532226
rect 97342 532170 97398 532226
rect 96970 532046 97026 532102
rect 97094 532046 97150 532102
rect 97218 532046 97274 532102
rect 97342 532046 97398 532102
rect 96970 531922 97026 531978
rect 97094 531922 97150 531978
rect 97218 531922 97274 531978
rect 97342 531922 97398 531978
rect 96970 514294 97026 514350
rect 97094 514294 97150 514350
rect 97218 514294 97274 514350
rect 97342 514294 97398 514350
rect 96970 514170 97026 514226
rect 97094 514170 97150 514226
rect 97218 514170 97274 514226
rect 97342 514170 97398 514226
rect 96970 514046 97026 514102
rect 97094 514046 97150 514102
rect 97218 514046 97274 514102
rect 97342 514046 97398 514102
rect 96970 513922 97026 513978
rect 97094 513922 97150 513978
rect 97218 513922 97274 513978
rect 97342 513922 97398 513978
rect 96970 496294 97026 496350
rect 97094 496294 97150 496350
rect 97218 496294 97274 496350
rect 97342 496294 97398 496350
rect 96970 496170 97026 496226
rect 97094 496170 97150 496226
rect 97218 496170 97274 496226
rect 97342 496170 97398 496226
rect 96970 496046 97026 496102
rect 97094 496046 97150 496102
rect 97218 496046 97274 496102
rect 97342 496046 97398 496102
rect 96970 495922 97026 495978
rect 97094 495922 97150 495978
rect 97218 495922 97274 495978
rect 97342 495922 97398 495978
rect 96970 478294 97026 478350
rect 97094 478294 97150 478350
rect 97218 478294 97274 478350
rect 97342 478294 97398 478350
rect 96970 478170 97026 478226
rect 97094 478170 97150 478226
rect 97218 478170 97274 478226
rect 97342 478170 97398 478226
rect 96970 478046 97026 478102
rect 97094 478046 97150 478102
rect 97218 478046 97274 478102
rect 97342 478046 97398 478102
rect 96970 477922 97026 477978
rect 97094 477922 97150 477978
rect 97218 477922 97274 477978
rect 97342 477922 97398 477978
rect 96970 460294 97026 460350
rect 97094 460294 97150 460350
rect 97218 460294 97274 460350
rect 97342 460294 97398 460350
rect 96970 460170 97026 460226
rect 97094 460170 97150 460226
rect 97218 460170 97274 460226
rect 97342 460170 97398 460226
rect 96970 460046 97026 460102
rect 97094 460046 97150 460102
rect 97218 460046 97274 460102
rect 97342 460046 97398 460102
rect 96970 459922 97026 459978
rect 97094 459922 97150 459978
rect 97218 459922 97274 459978
rect 97342 459922 97398 459978
rect 96970 442294 97026 442350
rect 97094 442294 97150 442350
rect 97218 442294 97274 442350
rect 97342 442294 97398 442350
rect 96970 442170 97026 442226
rect 97094 442170 97150 442226
rect 97218 442170 97274 442226
rect 97342 442170 97398 442226
rect 96970 442046 97026 442102
rect 97094 442046 97150 442102
rect 97218 442046 97274 442102
rect 97342 442046 97398 442102
rect 96970 441922 97026 441978
rect 97094 441922 97150 441978
rect 97218 441922 97274 441978
rect 97342 441922 97398 441978
rect 96970 424294 97026 424350
rect 97094 424294 97150 424350
rect 97218 424294 97274 424350
rect 97342 424294 97398 424350
rect 96970 424170 97026 424226
rect 97094 424170 97150 424226
rect 97218 424170 97274 424226
rect 97342 424170 97398 424226
rect 96970 424046 97026 424102
rect 97094 424046 97150 424102
rect 97218 424046 97274 424102
rect 97342 424046 97398 424102
rect 96970 423922 97026 423978
rect 97094 423922 97150 423978
rect 97218 423922 97274 423978
rect 97342 423922 97398 423978
rect 96970 406294 97026 406350
rect 97094 406294 97150 406350
rect 97218 406294 97274 406350
rect 97342 406294 97398 406350
rect 96970 406170 97026 406226
rect 97094 406170 97150 406226
rect 97218 406170 97274 406226
rect 97342 406170 97398 406226
rect 96970 406046 97026 406102
rect 97094 406046 97150 406102
rect 97218 406046 97274 406102
rect 97342 406046 97398 406102
rect 96970 405922 97026 405978
rect 97094 405922 97150 405978
rect 97218 405922 97274 405978
rect 97342 405922 97398 405978
rect 96970 388294 97026 388350
rect 97094 388294 97150 388350
rect 97218 388294 97274 388350
rect 97342 388294 97398 388350
rect 96970 388170 97026 388226
rect 97094 388170 97150 388226
rect 97218 388170 97274 388226
rect 97342 388170 97398 388226
rect 96970 388046 97026 388102
rect 97094 388046 97150 388102
rect 97218 388046 97274 388102
rect 97342 388046 97398 388102
rect 96970 387922 97026 387978
rect 97094 387922 97150 387978
rect 97218 387922 97274 387978
rect 97342 387922 97398 387978
rect 96970 370294 97026 370350
rect 97094 370294 97150 370350
rect 97218 370294 97274 370350
rect 97342 370294 97398 370350
rect 96970 370170 97026 370226
rect 97094 370170 97150 370226
rect 97218 370170 97274 370226
rect 97342 370170 97398 370226
rect 96970 370046 97026 370102
rect 97094 370046 97150 370102
rect 97218 370046 97274 370102
rect 97342 370046 97398 370102
rect 96970 369922 97026 369978
rect 97094 369922 97150 369978
rect 97218 369922 97274 369978
rect 97342 369922 97398 369978
rect 96970 352294 97026 352350
rect 97094 352294 97150 352350
rect 97218 352294 97274 352350
rect 97342 352294 97398 352350
rect 96970 352170 97026 352226
rect 97094 352170 97150 352226
rect 97218 352170 97274 352226
rect 97342 352170 97398 352226
rect 96970 352046 97026 352102
rect 97094 352046 97150 352102
rect 97218 352046 97274 352102
rect 97342 352046 97398 352102
rect 96970 351922 97026 351978
rect 97094 351922 97150 351978
rect 97218 351922 97274 351978
rect 97342 351922 97398 351978
rect 96970 334294 97026 334350
rect 97094 334294 97150 334350
rect 97218 334294 97274 334350
rect 97342 334294 97398 334350
rect 96970 334170 97026 334226
rect 97094 334170 97150 334226
rect 97218 334170 97274 334226
rect 97342 334170 97398 334226
rect 96970 334046 97026 334102
rect 97094 334046 97150 334102
rect 97218 334046 97274 334102
rect 97342 334046 97398 334102
rect 96970 333922 97026 333978
rect 97094 333922 97150 333978
rect 97218 333922 97274 333978
rect 97342 333922 97398 333978
rect 96970 316294 97026 316350
rect 97094 316294 97150 316350
rect 97218 316294 97274 316350
rect 97342 316294 97398 316350
rect 96970 316170 97026 316226
rect 97094 316170 97150 316226
rect 97218 316170 97274 316226
rect 97342 316170 97398 316226
rect 96970 316046 97026 316102
rect 97094 316046 97150 316102
rect 97218 316046 97274 316102
rect 97342 316046 97398 316102
rect 96970 315922 97026 315978
rect 97094 315922 97150 315978
rect 97218 315922 97274 315978
rect 97342 315922 97398 315978
rect 96970 298294 97026 298350
rect 97094 298294 97150 298350
rect 97218 298294 97274 298350
rect 97342 298294 97398 298350
rect 96970 298170 97026 298226
rect 97094 298170 97150 298226
rect 97218 298170 97274 298226
rect 97342 298170 97398 298226
rect 96970 298046 97026 298102
rect 97094 298046 97150 298102
rect 97218 298046 97274 298102
rect 97342 298046 97398 298102
rect 96970 297922 97026 297978
rect 97094 297922 97150 297978
rect 97218 297922 97274 297978
rect 97342 297922 97398 297978
rect 96970 280294 97026 280350
rect 97094 280294 97150 280350
rect 97218 280294 97274 280350
rect 97342 280294 97398 280350
rect 96970 280170 97026 280226
rect 97094 280170 97150 280226
rect 97218 280170 97274 280226
rect 97342 280170 97398 280226
rect 96970 280046 97026 280102
rect 97094 280046 97150 280102
rect 97218 280046 97274 280102
rect 97342 280046 97398 280102
rect 96970 279922 97026 279978
rect 97094 279922 97150 279978
rect 97218 279922 97274 279978
rect 97342 279922 97398 279978
rect 96970 262294 97026 262350
rect 97094 262294 97150 262350
rect 97218 262294 97274 262350
rect 97342 262294 97398 262350
rect 96970 262170 97026 262226
rect 97094 262170 97150 262226
rect 97218 262170 97274 262226
rect 97342 262170 97398 262226
rect 96970 262046 97026 262102
rect 97094 262046 97150 262102
rect 97218 262046 97274 262102
rect 97342 262046 97398 262102
rect 96970 261922 97026 261978
rect 97094 261922 97150 261978
rect 97218 261922 97274 261978
rect 97342 261922 97398 261978
rect 96970 244294 97026 244350
rect 97094 244294 97150 244350
rect 97218 244294 97274 244350
rect 97342 244294 97398 244350
rect 96970 244170 97026 244226
rect 97094 244170 97150 244226
rect 97218 244170 97274 244226
rect 97342 244170 97398 244226
rect 96970 244046 97026 244102
rect 97094 244046 97150 244102
rect 97218 244046 97274 244102
rect 97342 244046 97398 244102
rect 96970 243922 97026 243978
rect 97094 243922 97150 243978
rect 97218 243922 97274 243978
rect 97342 243922 97398 243978
rect 111250 597156 111306 597212
rect 111374 597156 111430 597212
rect 111498 597156 111554 597212
rect 111622 597156 111678 597212
rect 111250 597032 111306 597088
rect 111374 597032 111430 597088
rect 111498 597032 111554 597088
rect 111622 597032 111678 597088
rect 111250 596908 111306 596964
rect 111374 596908 111430 596964
rect 111498 596908 111554 596964
rect 111622 596908 111678 596964
rect 111250 596784 111306 596840
rect 111374 596784 111430 596840
rect 111498 596784 111554 596840
rect 111622 596784 111678 596840
rect 111250 580294 111306 580350
rect 111374 580294 111430 580350
rect 111498 580294 111554 580350
rect 111622 580294 111678 580350
rect 111250 580170 111306 580226
rect 111374 580170 111430 580226
rect 111498 580170 111554 580226
rect 111622 580170 111678 580226
rect 111250 580046 111306 580102
rect 111374 580046 111430 580102
rect 111498 580046 111554 580102
rect 111622 580046 111678 580102
rect 111250 579922 111306 579978
rect 111374 579922 111430 579978
rect 111498 579922 111554 579978
rect 111622 579922 111678 579978
rect 111250 562294 111306 562350
rect 111374 562294 111430 562350
rect 111498 562294 111554 562350
rect 111622 562294 111678 562350
rect 111250 562170 111306 562226
rect 111374 562170 111430 562226
rect 111498 562170 111554 562226
rect 111622 562170 111678 562226
rect 111250 562046 111306 562102
rect 111374 562046 111430 562102
rect 111498 562046 111554 562102
rect 111622 562046 111678 562102
rect 111250 561922 111306 561978
rect 111374 561922 111430 561978
rect 111498 561922 111554 561978
rect 111622 561922 111678 561978
rect 111250 544294 111306 544350
rect 111374 544294 111430 544350
rect 111498 544294 111554 544350
rect 111622 544294 111678 544350
rect 111250 544170 111306 544226
rect 111374 544170 111430 544226
rect 111498 544170 111554 544226
rect 111622 544170 111678 544226
rect 111250 544046 111306 544102
rect 111374 544046 111430 544102
rect 111498 544046 111554 544102
rect 111622 544046 111678 544102
rect 111250 543922 111306 543978
rect 111374 543922 111430 543978
rect 111498 543922 111554 543978
rect 111622 543922 111678 543978
rect 111250 526294 111306 526350
rect 111374 526294 111430 526350
rect 111498 526294 111554 526350
rect 111622 526294 111678 526350
rect 111250 526170 111306 526226
rect 111374 526170 111430 526226
rect 111498 526170 111554 526226
rect 111622 526170 111678 526226
rect 111250 526046 111306 526102
rect 111374 526046 111430 526102
rect 111498 526046 111554 526102
rect 111622 526046 111678 526102
rect 111250 525922 111306 525978
rect 111374 525922 111430 525978
rect 111498 525922 111554 525978
rect 111622 525922 111678 525978
rect 111250 508294 111306 508350
rect 111374 508294 111430 508350
rect 111498 508294 111554 508350
rect 111622 508294 111678 508350
rect 111250 508170 111306 508226
rect 111374 508170 111430 508226
rect 111498 508170 111554 508226
rect 111622 508170 111678 508226
rect 111250 508046 111306 508102
rect 111374 508046 111430 508102
rect 111498 508046 111554 508102
rect 111622 508046 111678 508102
rect 111250 507922 111306 507978
rect 111374 507922 111430 507978
rect 111498 507922 111554 507978
rect 111622 507922 111678 507978
rect 111250 490294 111306 490350
rect 111374 490294 111430 490350
rect 111498 490294 111554 490350
rect 111622 490294 111678 490350
rect 111250 490170 111306 490226
rect 111374 490170 111430 490226
rect 111498 490170 111554 490226
rect 111622 490170 111678 490226
rect 111250 490046 111306 490102
rect 111374 490046 111430 490102
rect 111498 490046 111554 490102
rect 111622 490046 111678 490102
rect 111250 489922 111306 489978
rect 111374 489922 111430 489978
rect 111498 489922 111554 489978
rect 111622 489922 111678 489978
rect 111250 472294 111306 472350
rect 111374 472294 111430 472350
rect 111498 472294 111554 472350
rect 111622 472294 111678 472350
rect 111250 472170 111306 472226
rect 111374 472170 111430 472226
rect 111498 472170 111554 472226
rect 111622 472170 111678 472226
rect 111250 472046 111306 472102
rect 111374 472046 111430 472102
rect 111498 472046 111554 472102
rect 111622 472046 111678 472102
rect 111250 471922 111306 471978
rect 111374 471922 111430 471978
rect 111498 471922 111554 471978
rect 111622 471922 111678 471978
rect 111250 454294 111306 454350
rect 111374 454294 111430 454350
rect 111498 454294 111554 454350
rect 111622 454294 111678 454350
rect 111250 454170 111306 454226
rect 111374 454170 111430 454226
rect 111498 454170 111554 454226
rect 111622 454170 111678 454226
rect 111250 454046 111306 454102
rect 111374 454046 111430 454102
rect 111498 454046 111554 454102
rect 111622 454046 111678 454102
rect 111250 453922 111306 453978
rect 111374 453922 111430 453978
rect 111498 453922 111554 453978
rect 111622 453922 111678 453978
rect 111250 436294 111306 436350
rect 111374 436294 111430 436350
rect 111498 436294 111554 436350
rect 111622 436294 111678 436350
rect 111250 436170 111306 436226
rect 111374 436170 111430 436226
rect 111498 436170 111554 436226
rect 111622 436170 111678 436226
rect 111250 436046 111306 436102
rect 111374 436046 111430 436102
rect 111498 436046 111554 436102
rect 111622 436046 111678 436102
rect 111250 435922 111306 435978
rect 111374 435922 111430 435978
rect 111498 435922 111554 435978
rect 111622 435922 111678 435978
rect 111250 418294 111306 418350
rect 111374 418294 111430 418350
rect 111498 418294 111554 418350
rect 111622 418294 111678 418350
rect 111250 418170 111306 418226
rect 111374 418170 111430 418226
rect 111498 418170 111554 418226
rect 111622 418170 111678 418226
rect 111250 418046 111306 418102
rect 111374 418046 111430 418102
rect 111498 418046 111554 418102
rect 111622 418046 111678 418102
rect 111250 417922 111306 417978
rect 111374 417922 111430 417978
rect 111498 417922 111554 417978
rect 111622 417922 111678 417978
rect 111250 400294 111306 400350
rect 111374 400294 111430 400350
rect 111498 400294 111554 400350
rect 111622 400294 111678 400350
rect 111250 400170 111306 400226
rect 111374 400170 111430 400226
rect 111498 400170 111554 400226
rect 111622 400170 111678 400226
rect 111250 400046 111306 400102
rect 111374 400046 111430 400102
rect 111498 400046 111554 400102
rect 111622 400046 111678 400102
rect 111250 399922 111306 399978
rect 111374 399922 111430 399978
rect 111498 399922 111554 399978
rect 111622 399922 111678 399978
rect 111250 382294 111306 382350
rect 111374 382294 111430 382350
rect 111498 382294 111554 382350
rect 111622 382294 111678 382350
rect 111250 382170 111306 382226
rect 111374 382170 111430 382226
rect 111498 382170 111554 382226
rect 111622 382170 111678 382226
rect 111250 382046 111306 382102
rect 111374 382046 111430 382102
rect 111498 382046 111554 382102
rect 111622 382046 111678 382102
rect 111250 381922 111306 381978
rect 111374 381922 111430 381978
rect 111498 381922 111554 381978
rect 111622 381922 111678 381978
rect 111250 364294 111306 364350
rect 111374 364294 111430 364350
rect 111498 364294 111554 364350
rect 111622 364294 111678 364350
rect 111250 364170 111306 364226
rect 111374 364170 111430 364226
rect 111498 364170 111554 364226
rect 111622 364170 111678 364226
rect 111250 364046 111306 364102
rect 111374 364046 111430 364102
rect 111498 364046 111554 364102
rect 111622 364046 111678 364102
rect 111250 363922 111306 363978
rect 111374 363922 111430 363978
rect 111498 363922 111554 363978
rect 111622 363922 111678 363978
rect 111250 346294 111306 346350
rect 111374 346294 111430 346350
rect 111498 346294 111554 346350
rect 111622 346294 111678 346350
rect 111250 346170 111306 346226
rect 111374 346170 111430 346226
rect 111498 346170 111554 346226
rect 111622 346170 111678 346226
rect 111250 346046 111306 346102
rect 111374 346046 111430 346102
rect 111498 346046 111554 346102
rect 111622 346046 111678 346102
rect 111250 345922 111306 345978
rect 111374 345922 111430 345978
rect 111498 345922 111554 345978
rect 111622 345922 111678 345978
rect 111250 328294 111306 328350
rect 111374 328294 111430 328350
rect 111498 328294 111554 328350
rect 111622 328294 111678 328350
rect 111250 328170 111306 328226
rect 111374 328170 111430 328226
rect 111498 328170 111554 328226
rect 111622 328170 111678 328226
rect 111250 328046 111306 328102
rect 111374 328046 111430 328102
rect 111498 328046 111554 328102
rect 111622 328046 111678 328102
rect 111250 327922 111306 327978
rect 111374 327922 111430 327978
rect 111498 327922 111554 327978
rect 111622 327922 111678 327978
rect 111250 310294 111306 310350
rect 111374 310294 111430 310350
rect 111498 310294 111554 310350
rect 111622 310294 111678 310350
rect 111250 310170 111306 310226
rect 111374 310170 111430 310226
rect 111498 310170 111554 310226
rect 111622 310170 111678 310226
rect 111250 310046 111306 310102
rect 111374 310046 111430 310102
rect 111498 310046 111554 310102
rect 111622 310046 111678 310102
rect 111250 309922 111306 309978
rect 111374 309922 111430 309978
rect 111498 309922 111554 309978
rect 111622 309922 111678 309978
rect 111250 292294 111306 292350
rect 111374 292294 111430 292350
rect 111498 292294 111554 292350
rect 111622 292294 111678 292350
rect 111250 292170 111306 292226
rect 111374 292170 111430 292226
rect 111498 292170 111554 292226
rect 111622 292170 111678 292226
rect 111250 292046 111306 292102
rect 111374 292046 111430 292102
rect 111498 292046 111554 292102
rect 111622 292046 111678 292102
rect 111250 291922 111306 291978
rect 111374 291922 111430 291978
rect 111498 291922 111554 291978
rect 111622 291922 111678 291978
rect 111250 274294 111306 274350
rect 111374 274294 111430 274350
rect 111498 274294 111554 274350
rect 111622 274294 111678 274350
rect 111250 274170 111306 274226
rect 111374 274170 111430 274226
rect 111498 274170 111554 274226
rect 111622 274170 111678 274226
rect 111250 274046 111306 274102
rect 111374 274046 111430 274102
rect 111498 274046 111554 274102
rect 111622 274046 111678 274102
rect 111250 273922 111306 273978
rect 111374 273922 111430 273978
rect 111498 273922 111554 273978
rect 111622 273922 111678 273978
rect 111250 256294 111306 256350
rect 111374 256294 111430 256350
rect 111498 256294 111554 256350
rect 111622 256294 111678 256350
rect 111250 256170 111306 256226
rect 111374 256170 111430 256226
rect 111498 256170 111554 256226
rect 111622 256170 111678 256226
rect 111250 256046 111306 256102
rect 111374 256046 111430 256102
rect 111498 256046 111554 256102
rect 111622 256046 111678 256102
rect 111250 255922 111306 255978
rect 111374 255922 111430 255978
rect 111498 255922 111554 255978
rect 111622 255922 111678 255978
rect 129250 597156 129306 597212
rect 129374 597156 129430 597212
rect 129498 597156 129554 597212
rect 129622 597156 129678 597212
rect 129250 597032 129306 597088
rect 129374 597032 129430 597088
rect 129498 597032 129554 597088
rect 129622 597032 129678 597088
rect 129250 596908 129306 596964
rect 129374 596908 129430 596964
rect 129498 596908 129554 596964
rect 129622 596908 129678 596964
rect 129250 596784 129306 596840
rect 129374 596784 129430 596840
rect 129498 596784 129554 596840
rect 129622 596784 129678 596840
rect 129250 580294 129306 580350
rect 129374 580294 129430 580350
rect 129498 580294 129554 580350
rect 129622 580294 129678 580350
rect 129250 580170 129306 580226
rect 129374 580170 129430 580226
rect 129498 580170 129554 580226
rect 129622 580170 129678 580226
rect 129250 580046 129306 580102
rect 129374 580046 129430 580102
rect 129498 580046 129554 580102
rect 129622 580046 129678 580102
rect 129250 579922 129306 579978
rect 129374 579922 129430 579978
rect 129498 579922 129554 579978
rect 129622 579922 129678 579978
rect 129250 562294 129306 562350
rect 129374 562294 129430 562350
rect 129498 562294 129554 562350
rect 129622 562294 129678 562350
rect 129250 562170 129306 562226
rect 129374 562170 129430 562226
rect 129498 562170 129554 562226
rect 129622 562170 129678 562226
rect 129250 562046 129306 562102
rect 129374 562046 129430 562102
rect 129498 562046 129554 562102
rect 129622 562046 129678 562102
rect 129250 561922 129306 561978
rect 129374 561922 129430 561978
rect 129498 561922 129554 561978
rect 129622 561922 129678 561978
rect 129250 544294 129306 544350
rect 129374 544294 129430 544350
rect 129498 544294 129554 544350
rect 129622 544294 129678 544350
rect 129250 544170 129306 544226
rect 129374 544170 129430 544226
rect 129498 544170 129554 544226
rect 129622 544170 129678 544226
rect 129250 544046 129306 544102
rect 129374 544046 129430 544102
rect 129498 544046 129554 544102
rect 129622 544046 129678 544102
rect 129250 543922 129306 543978
rect 129374 543922 129430 543978
rect 129498 543922 129554 543978
rect 129622 543922 129678 543978
rect 129250 526294 129306 526350
rect 129374 526294 129430 526350
rect 129498 526294 129554 526350
rect 129622 526294 129678 526350
rect 129250 526170 129306 526226
rect 129374 526170 129430 526226
rect 129498 526170 129554 526226
rect 129622 526170 129678 526226
rect 129250 526046 129306 526102
rect 129374 526046 129430 526102
rect 129498 526046 129554 526102
rect 129622 526046 129678 526102
rect 129250 525922 129306 525978
rect 129374 525922 129430 525978
rect 129498 525922 129554 525978
rect 129622 525922 129678 525978
rect 129250 508294 129306 508350
rect 129374 508294 129430 508350
rect 129498 508294 129554 508350
rect 129622 508294 129678 508350
rect 129250 508170 129306 508226
rect 129374 508170 129430 508226
rect 129498 508170 129554 508226
rect 129622 508170 129678 508226
rect 129250 508046 129306 508102
rect 129374 508046 129430 508102
rect 129498 508046 129554 508102
rect 129622 508046 129678 508102
rect 129250 507922 129306 507978
rect 129374 507922 129430 507978
rect 129498 507922 129554 507978
rect 129622 507922 129678 507978
rect 129250 490294 129306 490350
rect 129374 490294 129430 490350
rect 129498 490294 129554 490350
rect 129622 490294 129678 490350
rect 129250 490170 129306 490226
rect 129374 490170 129430 490226
rect 129498 490170 129554 490226
rect 129622 490170 129678 490226
rect 129250 490046 129306 490102
rect 129374 490046 129430 490102
rect 129498 490046 129554 490102
rect 129622 490046 129678 490102
rect 129250 489922 129306 489978
rect 129374 489922 129430 489978
rect 129498 489922 129554 489978
rect 129622 489922 129678 489978
rect 129250 472294 129306 472350
rect 129374 472294 129430 472350
rect 129498 472294 129554 472350
rect 129622 472294 129678 472350
rect 129250 472170 129306 472226
rect 129374 472170 129430 472226
rect 129498 472170 129554 472226
rect 129622 472170 129678 472226
rect 129250 472046 129306 472102
rect 129374 472046 129430 472102
rect 129498 472046 129554 472102
rect 129622 472046 129678 472102
rect 129250 471922 129306 471978
rect 129374 471922 129430 471978
rect 129498 471922 129554 471978
rect 129622 471922 129678 471978
rect 129250 454294 129306 454350
rect 129374 454294 129430 454350
rect 129498 454294 129554 454350
rect 129622 454294 129678 454350
rect 129250 454170 129306 454226
rect 129374 454170 129430 454226
rect 129498 454170 129554 454226
rect 129622 454170 129678 454226
rect 129250 454046 129306 454102
rect 129374 454046 129430 454102
rect 129498 454046 129554 454102
rect 129622 454046 129678 454102
rect 129250 453922 129306 453978
rect 129374 453922 129430 453978
rect 129498 453922 129554 453978
rect 129622 453922 129678 453978
rect 129250 436294 129306 436350
rect 129374 436294 129430 436350
rect 129498 436294 129554 436350
rect 129622 436294 129678 436350
rect 129250 436170 129306 436226
rect 129374 436170 129430 436226
rect 129498 436170 129554 436226
rect 129622 436170 129678 436226
rect 129250 436046 129306 436102
rect 129374 436046 129430 436102
rect 129498 436046 129554 436102
rect 129622 436046 129678 436102
rect 129250 435922 129306 435978
rect 129374 435922 129430 435978
rect 129498 435922 129554 435978
rect 129622 435922 129678 435978
rect 129250 418294 129306 418350
rect 129374 418294 129430 418350
rect 129498 418294 129554 418350
rect 129622 418294 129678 418350
rect 129250 418170 129306 418226
rect 129374 418170 129430 418226
rect 129498 418170 129554 418226
rect 129622 418170 129678 418226
rect 129250 418046 129306 418102
rect 129374 418046 129430 418102
rect 129498 418046 129554 418102
rect 129622 418046 129678 418102
rect 129250 417922 129306 417978
rect 129374 417922 129430 417978
rect 129498 417922 129554 417978
rect 129622 417922 129678 417978
rect 129250 400294 129306 400350
rect 129374 400294 129430 400350
rect 129498 400294 129554 400350
rect 129622 400294 129678 400350
rect 129250 400170 129306 400226
rect 129374 400170 129430 400226
rect 129498 400170 129554 400226
rect 129622 400170 129678 400226
rect 129250 400046 129306 400102
rect 129374 400046 129430 400102
rect 129498 400046 129554 400102
rect 129622 400046 129678 400102
rect 129250 399922 129306 399978
rect 129374 399922 129430 399978
rect 129498 399922 129554 399978
rect 129622 399922 129678 399978
rect 129250 382294 129306 382350
rect 129374 382294 129430 382350
rect 129498 382294 129554 382350
rect 129622 382294 129678 382350
rect 129250 382170 129306 382226
rect 129374 382170 129430 382226
rect 129498 382170 129554 382226
rect 129622 382170 129678 382226
rect 129250 382046 129306 382102
rect 129374 382046 129430 382102
rect 129498 382046 129554 382102
rect 129622 382046 129678 382102
rect 129250 381922 129306 381978
rect 129374 381922 129430 381978
rect 129498 381922 129554 381978
rect 129622 381922 129678 381978
rect 129250 364294 129306 364350
rect 129374 364294 129430 364350
rect 129498 364294 129554 364350
rect 129622 364294 129678 364350
rect 129250 364170 129306 364226
rect 129374 364170 129430 364226
rect 129498 364170 129554 364226
rect 129622 364170 129678 364226
rect 129250 364046 129306 364102
rect 129374 364046 129430 364102
rect 129498 364046 129554 364102
rect 129622 364046 129678 364102
rect 129250 363922 129306 363978
rect 129374 363922 129430 363978
rect 129498 363922 129554 363978
rect 129622 363922 129678 363978
rect 129250 346294 129306 346350
rect 129374 346294 129430 346350
rect 129498 346294 129554 346350
rect 129622 346294 129678 346350
rect 129250 346170 129306 346226
rect 129374 346170 129430 346226
rect 129498 346170 129554 346226
rect 129622 346170 129678 346226
rect 129250 346046 129306 346102
rect 129374 346046 129430 346102
rect 129498 346046 129554 346102
rect 129622 346046 129678 346102
rect 129250 345922 129306 345978
rect 129374 345922 129430 345978
rect 129498 345922 129554 345978
rect 129622 345922 129678 345978
rect 129250 328294 129306 328350
rect 129374 328294 129430 328350
rect 129498 328294 129554 328350
rect 129622 328294 129678 328350
rect 129250 328170 129306 328226
rect 129374 328170 129430 328226
rect 129498 328170 129554 328226
rect 129622 328170 129678 328226
rect 129250 328046 129306 328102
rect 129374 328046 129430 328102
rect 129498 328046 129554 328102
rect 129622 328046 129678 328102
rect 129250 327922 129306 327978
rect 129374 327922 129430 327978
rect 129498 327922 129554 327978
rect 129622 327922 129678 327978
rect 129250 310294 129306 310350
rect 129374 310294 129430 310350
rect 129498 310294 129554 310350
rect 129622 310294 129678 310350
rect 129250 310170 129306 310226
rect 129374 310170 129430 310226
rect 129498 310170 129554 310226
rect 129622 310170 129678 310226
rect 129250 310046 129306 310102
rect 129374 310046 129430 310102
rect 129498 310046 129554 310102
rect 129622 310046 129678 310102
rect 129250 309922 129306 309978
rect 129374 309922 129430 309978
rect 129498 309922 129554 309978
rect 129622 309922 129678 309978
rect 129250 292294 129306 292350
rect 129374 292294 129430 292350
rect 129498 292294 129554 292350
rect 129622 292294 129678 292350
rect 129250 292170 129306 292226
rect 129374 292170 129430 292226
rect 129498 292170 129554 292226
rect 129622 292170 129678 292226
rect 129250 292046 129306 292102
rect 129374 292046 129430 292102
rect 129498 292046 129554 292102
rect 129622 292046 129678 292102
rect 129250 291922 129306 291978
rect 129374 291922 129430 291978
rect 129498 291922 129554 291978
rect 129622 291922 129678 291978
rect 129250 274294 129306 274350
rect 129374 274294 129430 274350
rect 129498 274294 129554 274350
rect 129622 274294 129678 274350
rect 129250 274170 129306 274226
rect 129374 274170 129430 274226
rect 129498 274170 129554 274226
rect 129622 274170 129678 274226
rect 129250 274046 129306 274102
rect 129374 274046 129430 274102
rect 129498 274046 129554 274102
rect 129622 274046 129678 274102
rect 129250 273922 129306 273978
rect 129374 273922 129430 273978
rect 129498 273922 129554 273978
rect 129622 273922 129678 273978
rect 129250 256294 129306 256350
rect 129374 256294 129430 256350
rect 129498 256294 129554 256350
rect 129622 256294 129678 256350
rect 129250 256170 129306 256226
rect 129374 256170 129430 256226
rect 129498 256170 129554 256226
rect 129622 256170 129678 256226
rect 129250 256046 129306 256102
rect 129374 256046 129430 256102
rect 129498 256046 129554 256102
rect 129622 256046 129678 256102
rect 129250 255922 129306 255978
rect 129374 255922 129430 255978
rect 129498 255922 129554 255978
rect 129622 255922 129678 255978
rect 111250 238294 111306 238350
rect 111374 238294 111430 238350
rect 111498 238294 111554 238350
rect 111622 238294 111678 238350
rect 111250 238170 111306 238226
rect 111374 238170 111430 238226
rect 111498 238170 111554 238226
rect 111622 238170 111678 238226
rect 111250 238046 111306 238102
rect 111374 238046 111430 238102
rect 111498 238046 111554 238102
rect 111622 238046 111678 238102
rect 111250 237922 111306 237978
rect 111374 237922 111430 237978
rect 111498 237922 111554 237978
rect 111622 237922 111678 237978
rect 96970 226294 97026 226350
rect 97094 226294 97150 226350
rect 97218 226294 97274 226350
rect 97342 226294 97398 226350
rect 96970 226170 97026 226226
rect 97094 226170 97150 226226
rect 97218 226170 97274 226226
rect 97342 226170 97398 226226
rect 96970 226046 97026 226102
rect 97094 226046 97150 226102
rect 97218 226046 97274 226102
rect 97342 226046 97398 226102
rect 96970 225922 97026 225978
rect 97094 225922 97150 225978
rect 97218 225922 97274 225978
rect 97342 225922 97398 225978
rect 93250 220294 93306 220350
rect 93374 220294 93430 220350
rect 93498 220294 93554 220350
rect 93622 220294 93678 220350
rect 93250 220170 93306 220226
rect 93374 220170 93430 220226
rect 93498 220170 93554 220226
rect 93622 220170 93678 220226
rect 93250 220046 93306 220102
rect 93374 220046 93430 220102
rect 93498 220046 93554 220102
rect 93622 220046 93678 220102
rect 93250 219922 93306 219978
rect 93374 219922 93430 219978
rect 93498 219922 93554 219978
rect 93622 219922 93678 219978
rect 95238 220294 95294 220350
rect 95362 220294 95418 220350
rect 95238 220170 95294 220226
rect 95362 220170 95418 220226
rect 95238 220046 95294 220102
rect 95362 220046 95418 220102
rect 95238 219922 95294 219978
rect 95362 219922 95418 219978
rect 110598 226294 110654 226350
rect 110722 226294 110778 226350
rect 110598 226170 110654 226226
rect 110722 226170 110778 226226
rect 110598 226046 110654 226102
rect 110722 226046 110778 226102
rect 110598 225922 110654 225978
rect 110722 225922 110778 225978
rect 111250 220294 111306 220350
rect 111374 220294 111430 220350
rect 111498 220294 111554 220350
rect 111622 220294 111678 220350
rect 111250 220170 111306 220226
rect 111374 220170 111430 220226
rect 111498 220170 111554 220226
rect 111622 220170 111678 220226
rect 111250 220046 111306 220102
rect 111374 220046 111430 220102
rect 111498 220046 111554 220102
rect 111622 220046 111678 220102
rect 111250 219922 111306 219978
rect 111374 219922 111430 219978
rect 111498 219922 111554 219978
rect 111622 219922 111678 219978
rect 114970 226294 115026 226350
rect 115094 226294 115150 226350
rect 115218 226294 115274 226350
rect 115342 226294 115398 226350
rect 114970 226170 115026 226226
rect 115094 226170 115150 226226
rect 115218 226170 115274 226226
rect 115342 226170 115398 226226
rect 114970 226046 115026 226102
rect 115094 226046 115150 226102
rect 115218 226046 115274 226102
rect 115342 226046 115398 226102
rect 114970 225922 115026 225978
rect 115094 225922 115150 225978
rect 115218 225922 115274 225978
rect 115342 225922 115398 225978
rect 129250 238294 129306 238350
rect 129374 238294 129430 238350
rect 129498 238294 129554 238350
rect 129622 238294 129678 238350
rect 129250 238170 129306 238226
rect 129374 238170 129430 238226
rect 129498 238170 129554 238226
rect 129622 238170 129678 238226
rect 129250 238046 129306 238102
rect 129374 238046 129430 238102
rect 129498 238046 129554 238102
rect 129622 238046 129678 238102
rect 129250 237922 129306 237978
rect 129374 237922 129430 237978
rect 129498 237922 129554 237978
rect 129622 237922 129678 237978
rect 125958 220294 126014 220350
rect 126082 220294 126138 220350
rect 125958 220170 126014 220226
rect 126082 220170 126138 220226
rect 125958 220046 126014 220102
rect 126082 220046 126138 220102
rect 125958 219922 126014 219978
rect 126082 219922 126138 219978
rect 129250 220294 129306 220350
rect 129374 220294 129430 220350
rect 129498 220294 129554 220350
rect 129622 220294 129678 220350
rect 129250 220170 129306 220226
rect 129374 220170 129430 220226
rect 129498 220170 129554 220226
rect 129622 220170 129678 220226
rect 129250 220046 129306 220102
rect 129374 220046 129430 220102
rect 129498 220046 129554 220102
rect 129622 220046 129678 220102
rect 129250 219922 129306 219978
rect 129374 219922 129430 219978
rect 129498 219922 129554 219978
rect 129622 219922 129678 219978
rect 132970 598116 133026 598172
rect 133094 598116 133150 598172
rect 133218 598116 133274 598172
rect 133342 598116 133398 598172
rect 132970 597992 133026 598048
rect 133094 597992 133150 598048
rect 133218 597992 133274 598048
rect 133342 597992 133398 598048
rect 132970 597868 133026 597924
rect 133094 597868 133150 597924
rect 133218 597868 133274 597924
rect 133342 597868 133398 597924
rect 132970 597744 133026 597800
rect 133094 597744 133150 597800
rect 133218 597744 133274 597800
rect 133342 597744 133398 597800
rect 132970 586294 133026 586350
rect 133094 586294 133150 586350
rect 133218 586294 133274 586350
rect 133342 586294 133398 586350
rect 132970 586170 133026 586226
rect 133094 586170 133150 586226
rect 133218 586170 133274 586226
rect 133342 586170 133398 586226
rect 132970 586046 133026 586102
rect 133094 586046 133150 586102
rect 133218 586046 133274 586102
rect 133342 586046 133398 586102
rect 132970 585922 133026 585978
rect 133094 585922 133150 585978
rect 133218 585922 133274 585978
rect 133342 585922 133398 585978
rect 132970 568294 133026 568350
rect 133094 568294 133150 568350
rect 133218 568294 133274 568350
rect 133342 568294 133398 568350
rect 132970 568170 133026 568226
rect 133094 568170 133150 568226
rect 133218 568170 133274 568226
rect 133342 568170 133398 568226
rect 132970 568046 133026 568102
rect 133094 568046 133150 568102
rect 133218 568046 133274 568102
rect 133342 568046 133398 568102
rect 132970 567922 133026 567978
rect 133094 567922 133150 567978
rect 133218 567922 133274 567978
rect 133342 567922 133398 567978
rect 132970 550294 133026 550350
rect 133094 550294 133150 550350
rect 133218 550294 133274 550350
rect 133342 550294 133398 550350
rect 132970 550170 133026 550226
rect 133094 550170 133150 550226
rect 133218 550170 133274 550226
rect 133342 550170 133398 550226
rect 132970 550046 133026 550102
rect 133094 550046 133150 550102
rect 133218 550046 133274 550102
rect 133342 550046 133398 550102
rect 132970 549922 133026 549978
rect 133094 549922 133150 549978
rect 133218 549922 133274 549978
rect 133342 549922 133398 549978
rect 132970 532294 133026 532350
rect 133094 532294 133150 532350
rect 133218 532294 133274 532350
rect 133342 532294 133398 532350
rect 132970 532170 133026 532226
rect 133094 532170 133150 532226
rect 133218 532170 133274 532226
rect 133342 532170 133398 532226
rect 132970 532046 133026 532102
rect 133094 532046 133150 532102
rect 133218 532046 133274 532102
rect 133342 532046 133398 532102
rect 132970 531922 133026 531978
rect 133094 531922 133150 531978
rect 133218 531922 133274 531978
rect 133342 531922 133398 531978
rect 132970 514294 133026 514350
rect 133094 514294 133150 514350
rect 133218 514294 133274 514350
rect 133342 514294 133398 514350
rect 132970 514170 133026 514226
rect 133094 514170 133150 514226
rect 133218 514170 133274 514226
rect 133342 514170 133398 514226
rect 132970 514046 133026 514102
rect 133094 514046 133150 514102
rect 133218 514046 133274 514102
rect 133342 514046 133398 514102
rect 132970 513922 133026 513978
rect 133094 513922 133150 513978
rect 133218 513922 133274 513978
rect 133342 513922 133398 513978
rect 132970 496294 133026 496350
rect 133094 496294 133150 496350
rect 133218 496294 133274 496350
rect 133342 496294 133398 496350
rect 132970 496170 133026 496226
rect 133094 496170 133150 496226
rect 133218 496170 133274 496226
rect 133342 496170 133398 496226
rect 132970 496046 133026 496102
rect 133094 496046 133150 496102
rect 133218 496046 133274 496102
rect 133342 496046 133398 496102
rect 132970 495922 133026 495978
rect 133094 495922 133150 495978
rect 133218 495922 133274 495978
rect 133342 495922 133398 495978
rect 132970 478294 133026 478350
rect 133094 478294 133150 478350
rect 133218 478294 133274 478350
rect 133342 478294 133398 478350
rect 132970 478170 133026 478226
rect 133094 478170 133150 478226
rect 133218 478170 133274 478226
rect 133342 478170 133398 478226
rect 132970 478046 133026 478102
rect 133094 478046 133150 478102
rect 133218 478046 133274 478102
rect 133342 478046 133398 478102
rect 132970 477922 133026 477978
rect 133094 477922 133150 477978
rect 133218 477922 133274 477978
rect 133342 477922 133398 477978
rect 132970 460294 133026 460350
rect 133094 460294 133150 460350
rect 133218 460294 133274 460350
rect 133342 460294 133398 460350
rect 132970 460170 133026 460226
rect 133094 460170 133150 460226
rect 133218 460170 133274 460226
rect 133342 460170 133398 460226
rect 132970 460046 133026 460102
rect 133094 460046 133150 460102
rect 133218 460046 133274 460102
rect 133342 460046 133398 460102
rect 132970 459922 133026 459978
rect 133094 459922 133150 459978
rect 133218 459922 133274 459978
rect 133342 459922 133398 459978
rect 132970 442294 133026 442350
rect 133094 442294 133150 442350
rect 133218 442294 133274 442350
rect 133342 442294 133398 442350
rect 132970 442170 133026 442226
rect 133094 442170 133150 442226
rect 133218 442170 133274 442226
rect 133342 442170 133398 442226
rect 132970 442046 133026 442102
rect 133094 442046 133150 442102
rect 133218 442046 133274 442102
rect 133342 442046 133398 442102
rect 132970 441922 133026 441978
rect 133094 441922 133150 441978
rect 133218 441922 133274 441978
rect 133342 441922 133398 441978
rect 132970 424294 133026 424350
rect 133094 424294 133150 424350
rect 133218 424294 133274 424350
rect 133342 424294 133398 424350
rect 132970 424170 133026 424226
rect 133094 424170 133150 424226
rect 133218 424170 133274 424226
rect 133342 424170 133398 424226
rect 132970 424046 133026 424102
rect 133094 424046 133150 424102
rect 133218 424046 133274 424102
rect 133342 424046 133398 424102
rect 132970 423922 133026 423978
rect 133094 423922 133150 423978
rect 133218 423922 133274 423978
rect 133342 423922 133398 423978
rect 132970 406294 133026 406350
rect 133094 406294 133150 406350
rect 133218 406294 133274 406350
rect 133342 406294 133398 406350
rect 132970 406170 133026 406226
rect 133094 406170 133150 406226
rect 133218 406170 133274 406226
rect 133342 406170 133398 406226
rect 132970 406046 133026 406102
rect 133094 406046 133150 406102
rect 133218 406046 133274 406102
rect 133342 406046 133398 406102
rect 132970 405922 133026 405978
rect 133094 405922 133150 405978
rect 133218 405922 133274 405978
rect 133342 405922 133398 405978
rect 132970 388294 133026 388350
rect 133094 388294 133150 388350
rect 133218 388294 133274 388350
rect 133342 388294 133398 388350
rect 132970 388170 133026 388226
rect 133094 388170 133150 388226
rect 133218 388170 133274 388226
rect 133342 388170 133398 388226
rect 132970 388046 133026 388102
rect 133094 388046 133150 388102
rect 133218 388046 133274 388102
rect 133342 388046 133398 388102
rect 132970 387922 133026 387978
rect 133094 387922 133150 387978
rect 133218 387922 133274 387978
rect 133342 387922 133398 387978
rect 132970 370294 133026 370350
rect 133094 370294 133150 370350
rect 133218 370294 133274 370350
rect 133342 370294 133398 370350
rect 132970 370170 133026 370226
rect 133094 370170 133150 370226
rect 133218 370170 133274 370226
rect 133342 370170 133398 370226
rect 132970 370046 133026 370102
rect 133094 370046 133150 370102
rect 133218 370046 133274 370102
rect 133342 370046 133398 370102
rect 132970 369922 133026 369978
rect 133094 369922 133150 369978
rect 133218 369922 133274 369978
rect 133342 369922 133398 369978
rect 132970 352294 133026 352350
rect 133094 352294 133150 352350
rect 133218 352294 133274 352350
rect 133342 352294 133398 352350
rect 132970 352170 133026 352226
rect 133094 352170 133150 352226
rect 133218 352170 133274 352226
rect 133342 352170 133398 352226
rect 132970 352046 133026 352102
rect 133094 352046 133150 352102
rect 133218 352046 133274 352102
rect 133342 352046 133398 352102
rect 132970 351922 133026 351978
rect 133094 351922 133150 351978
rect 133218 351922 133274 351978
rect 133342 351922 133398 351978
rect 132970 334294 133026 334350
rect 133094 334294 133150 334350
rect 133218 334294 133274 334350
rect 133342 334294 133398 334350
rect 132970 334170 133026 334226
rect 133094 334170 133150 334226
rect 133218 334170 133274 334226
rect 133342 334170 133398 334226
rect 132970 334046 133026 334102
rect 133094 334046 133150 334102
rect 133218 334046 133274 334102
rect 133342 334046 133398 334102
rect 132970 333922 133026 333978
rect 133094 333922 133150 333978
rect 133218 333922 133274 333978
rect 133342 333922 133398 333978
rect 132970 316294 133026 316350
rect 133094 316294 133150 316350
rect 133218 316294 133274 316350
rect 133342 316294 133398 316350
rect 132970 316170 133026 316226
rect 133094 316170 133150 316226
rect 133218 316170 133274 316226
rect 133342 316170 133398 316226
rect 132970 316046 133026 316102
rect 133094 316046 133150 316102
rect 133218 316046 133274 316102
rect 133342 316046 133398 316102
rect 132970 315922 133026 315978
rect 133094 315922 133150 315978
rect 133218 315922 133274 315978
rect 133342 315922 133398 315978
rect 132970 298294 133026 298350
rect 133094 298294 133150 298350
rect 133218 298294 133274 298350
rect 133342 298294 133398 298350
rect 132970 298170 133026 298226
rect 133094 298170 133150 298226
rect 133218 298170 133274 298226
rect 133342 298170 133398 298226
rect 132970 298046 133026 298102
rect 133094 298046 133150 298102
rect 133218 298046 133274 298102
rect 133342 298046 133398 298102
rect 132970 297922 133026 297978
rect 133094 297922 133150 297978
rect 133218 297922 133274 297978
rect 133342 297922 133398 297978
rect 132970 280294 133026 280350
rect 133094 280294 133150 280350
rect 133218 280294 133274 280350
rect 133342 280294 133398 280350
rect 132970 280170 133026 280226
rect 133094 280170 133150 280226
rect 133218 280170 133274 280226
rect 133342 280170 133398 280226
rect 132970 280046 133026 280102
rect 133094 280046 133150 280102
rect 133218 280046 133274 280102
rect 133342 280046 133398 280102
rect 132970 279922 133026 279978
rect 133094 279922 133150 279978
rect 133218 279922 133274 279978
rect 133342 279922 133398 279978
rect 132970 262294 133026 262350
rect 133094 262294 133150 262350
rect 133218 262294 133274 262350
rect 133342 262294 133398 262350
rect 132970 262170 133026 262226
rect 133094 262170 133150 262226
rect 133218 262170 133274 262226
rect 133342 262170 133398 262226
rect 132970 262046 133026 262102
rect 133094 262046 133150 262102
rect 133218 262046 133274 262102
rect 133342 262046 133398 262102
rect 132970 261922 133026 261978
rect 133094 261922 133150 261978
rect 133218 261922 133274 261978
rect 133342 261922 133398 261978
rect 132970 244294 133026 244350
rect 133094 244294 133150 244350
rect 133218 244294 133274 244350
rect 133342 244294 133398 244350
rect 132970 244170 133026 244226
rect 133094 244170 133150 244226
rect 133218 244170 133274 244226
rect 133342 244170 133398 244226
rect 132970 244046 133026 244102
rect 133094 244046 133150 244102
rect 133218 244046 133274 244102
rect 133342 244046 133398 244102
rect 132970 243922 133026 243978
rect 133094 243922 133150 243978
rect 133218 243922 133274 243978
rect 133342 243922 133398 243978
rect 147250 597156 147306 597212
rect 147374 597156 147430 597212
rect 147498 597156 147554 597212
rect 147622 597156 147678 597212
rect 147250 597032 147306 597088
rect 147374 597032 147430 597088
rect 147498 597032 147554 597088
rect 147622 597032 147678 597088
rect 147250 596908 147306 596964
rect 147374 596908 147430 596964
rect 147498 596908 147554 596964
rect 147622 596908 147678 596964
rect 147250 596784 147306 596840
rect 147374 596784 147430 596840
rect 147498 596784 147554 596840
rect 147622 596784 147678 596840
rect 147250 580294 147306 580350
rect 147374 580294 147430 580350
rect 147498 580294 147554 580350
rect 147622 580294 147678 580350
rect 147250 580170 147306 580226
rect 147374 580170 147430 580226
rect 147498 580170 147554 580226
rect 147622 580170 147678 580226
rect 147250 580046 147306 580102
rect 147374 580046 147430 580102
rect 147498 580046 147554 580102
rect 147622 580046 147678 580102
rect 147250 579922 147306 579978
rect 147374 579922 147430 579978
rect 147498 579922 147554 579978
rect 147622 579922 147678 579978
rect 147250 562294 147306 562350
rect 147374 562294 147430 562350
rect 147498 562294 147554 562350
rect 147622 562294 147678 562350
rect 147250 562170 147306 562226
rect 147374 562170 147430 562226
rect 147498 562170 147554 562226
rect 147622 562170 147678 562226
rect 147250 562046 147306 562102
rect 147374 562046 147430 562102
rect 147498 562046 147554 562102
rect 147622 562046 147678 562102
rect 147250 561922 147306 561978
rect 147374 561922 147430 561978
rect 147498 561922 147554 561978
rect 147622 561922 147678 561978
rect 147250 544294 147306 544350
rect 147374 544294 147430 544350
rect 147498 544294 147554 544350
rect 147622 544294 147678 544350
rect 147250 544170 147306 544226
rect 147374 544170 147430 544226
rect 147498 544170 147554 544226
rect 147622 544170 147678 544226
rect 147250 544046 147306 544102
rect 147374 544046 147430 544102
rect 147498 544046 147554 544102
rect 147622 544046 147678 544102
rect 147250 543922 147306 543978
rect 147374 543922 147430 543978
rect 147498 543922 147554 543978
rect 147622 543922 147678 543978
rect 147250 526294 147306 526350
rect 147374 526294 147430 526350
rect 147498 526294 147554 526350
rect 147622 526294 147678 526350
rect 147250 526170 147306 526226
rect 147374 526170 147430 526226
rect 147498 526170 147554 526226
rect 147622 526170 147678 526226
rect 147250 526046 147306 526102
rect 147374 526046 147430 526102
rect 147498 526046 147554 526102
rect 147622 526046 147678 526102
rect 147250 525922 147306 525978
rect 147374 525922 147430 525978
rect 147498 525922 147554 525978
rect 147622 525922 147678 525978
rect 147250 508294 147306 508350
rect 147374 508294 147430 508350
rect 147498 508294 147554 508350
rect 147622 508294 147678 508350
rect 147250 508170 147306 508226
rect 147374 508170 147430 508226
rect 147498 508170 147554 508226
rect 147622 508170 147678 508226
rect 147250 508046 147306 508102
rect 147374 508046 147430 508102
rect 147498 508046 147554 508102
rect 147622 508046 147678 508102
rect 147250 507922 147306 507978
rect 147374 507922 147430 507978
rect 147498 507922 147554 507978
rect 147622 507922 147678 507978
rect 147250 490294 147306 490350
rect 147374 490294 147430 490350
rect 147498 490294 147554 490350
rect 147622 490294 147678 490350
rect 147250 490170 147306 490226
rect 147374 490170 147430 490226
rect 147498 490170 147554 490226
rect 147622 490170 147678 490226
rect 147250 490046 147306 490102
rect 147374 490046 147430 490102
rect 147498 490046 147554 490102
rect 147622 490046 147678 490102
rect 147250 489922 147306 489978
rect 147374 489922 147430 489978
rect 147498 489922 147554 489978
rect 147622 489922 147678 489978
rect 147250 472294 147306 472350
rect 147374 472294 147430 472350
rect 147498 472294 147554 472350
rect 147622 472294 147678 472350
rect 147250 472170 147306 472226
rect 147374 472170 147430 472226
rect 147498 472170 147554 472226
rect 147622 472170 147678 472226
rect 147250 472046 147306 472102
rect 147374 472046 147430 472102
rect 147498 472046 147554 472102
rect 147622 472046 147678 472102
rect 147250 471922 147306 471978
rect 147374 471922 147430 471978
rect 147498 471922 147554 471978
rect 147622 471922 147678 471978
rect 147250 454294 147306 454350
rect 147374 454294 147430 454350
rect 147498 454294 147554 454350
rect 147622 454294 147678 454350
rect 147250 454170 147306 454226
rect 147374 454170 147430 454226
rect 147498 454170 147554 454226
rect 147622 454170 147678 454226
rect 147250 454046 147306 454102
rect 147374 454046 147430 454102
rect 147498 454046 147554 454102
rect 147622 454046 147678 454102
rect 147250 453922 147306 453978
rect 147374 453922 147430 453978
rect 147498 453922 147554 453978
rect 147622 453922 147678 453978
rect 147250 436294 147306 436350
rect 147374 436294 147430 436350
rect 147498 436294 147554 436350
rect 147622 436294 147678 436350
rect 147250 436170 147306 436226
rect 147374 436170 147430 436226
rect 147498 436170 147554 436226
rect 147622 436170 147678 436226
rect 147250 436046 147306 436102
rect 147374 436046 147430 436102
rect 147498 436046 147554 436102
rect 147622 436046 147678 436102
rect 147250 435922 147306 435978
rect 147374 435922 147430 435978
rect 147498 435922 147554 435978
rect 147622 435922 147678 435978
rect 147250 418294 147306 418350
rect 147374 418294 147430 418350
rect 147498 418294 147554 418350
rect 147622 418294 147678 418350
rect 147250 418170 147306 418226
rect 147374 418170 147430 418226
rect 147498 418170 147554 418226
rect 147622 418170 147678 418226
rect 147250 418046 147306 418102
rect 147374 418046 147430 418102
rect 147498 418046 147554 418102
rect 147622 418046 147678 418102
rect 147250 417922 147306 417978
rect 147374 417922 147430 417978
rect 147498 417922 147554 417978
rect 147622 417922 147678 417978
rect 147250 400294 147306 400350
rect 147374 400294 147430 400350
rect 147498 400294 147554 400350
rect 147622 400294 147678 400350
rect 147250 400170 147306 400226
rect 147374 400170 147430 400226
rect 147498 400170 147554 400226
rect 147622 400170 147678 400226
rect 147250 400046 147306 400102
rect 147374 400046 147430 400102
rect 147498 400046 147554 400102
rect 147622 400046 147678 400102
rect 147250 399922 147306 399978
rect 147374 399922 147430 399978
rect 147498 399922 147554 399978
rect 147622 399922 147678 399978
rect 147250 382294 147306 382350
rect 147374 382294 147430 382350
rect 147498 382294 147554 382350
rect 147622 382294 147678 382350
rect 147250 382170 147306 382226
rect 147374 382170 147430 382226
rect 147498 382170 147554 382226
rect 147622 382170 147678 382226
rect 147250 382046 147306 382102
rect 147374 382046 147430 382102
rect 147498 382046 147554 382102
rect 147622 382046 147678 382102
rect 147250 381922 147306 381978
rect 147374 381922 147430 381978
rect 147498 381922 147554 381978
rect 147622 381922 147678 381978
rect 147250 364294 147306 364350
rect 147374 364294 147430 364350
rect 147498 364294 147554 364350
rect 147622 364294 147678 364350
rect 147250 364170 147306 364226
rect 147374 364170 147430 364226
rect 147498 364170 147554 364226
rect 147622 364170 147678 364226
rect 147250 364046 147306 364102
rect 147374 364046 147430 364102
rect 147498 364046 147554 364102
rect 147622 364046 147678 364102
rect 147250 363922 147306 363978
rect 147374 363922 147430 363978
rect 147498 363922 147554 363978
rect 147622 363922 147678 363978
rect 147250 346294 147306 346350
rect 147374 346294 147430 346350
rect 147498 346294 147554 346350
rect 147622 346294 147678 346350
rect 147250 346170 147306 346226
rect 147374 346170 147430 346226
rect 147498 346170 147554 346226
rect 147622 346170 147678 346226
rect 147250 346046 147306 346102
rect 147374 346046 147430 346102
rect 147498 346046 147554 346102
rect 147622 346046 147678 346102
rect 147250 345922 147306 345978
rect 147374 345922 147430 345978
rect 147498 345922 147554 345978
rect 147622 345922 147678 345978
rect 147250 328294 147306 328350
rect 147374 328294 147430 328350
rect 147498 328294 147554 328350
rect 147622 328294 147678 328350
rect 147250 328170 147306 328226
rect 147374 328170 147430 328226
rect 147498 328170 147554 328226
rect 147622 328170 147678 328226
rect 147250 328046 147306 328102
rect 147374 328046 147430 328102
rect 147498 328046 147554 328102
rect 147622 328046 147678 328102
rect 147250 327922 147306 327978
rect 147374 327922 147430 327978
rect 147498 327922 147554 327978
rect 147622 327922 147678 327978
rect 147250 310294 147306 310350
rect 147374 310294 147430 310350
rect 147498 310294 147554 310350
rect 147622 310294 147678 310350
rect 147250 310170 147306 310226
rect 147374 310170 147430 310226
rect 147498 310170 147554 310226
rect 147622 310170 147678 310226
rect 147250 310046 147306 310102
rect 147374 310046 147430 310102
rect 147498 310046 147554 310102
rect 147622 310046 147678 310102
rect 147250 309922 147306 309978
rect 147374 309922 147430 309978
rect 147498 309922 147554 309978
rect 147622 309922 147678 309978
rect 147250 292294 147306 292350
rect 147374 292294 147430 292350
rect 147498 292294 147554 292350
rect 147622 292294 147678 292350
rect 147250 292170 147306 292226
rect 147374 292170 147430 292226
rect 147498 292170 147554 292226
rect 147622 292170 147678 292226
rect 147250 292046 147306 292102
rect 147374 292046 147430 292102
rect 147498 292046 147554 292102
rect 147622 292046 147678 292102
rect 147250 291922 147306 291978
rect 147374 291922 147430 291978
rect 147498 291922 147554 291978
rect 147622 291922 147678 291978
rect 147250 274294 147306 274350
rect 147374 274294 147430 274350
rect 147498 274294 147554 274350
rect 147622 274294 147678 274350
rect 147250 274170 147306 274226
rect 147374 274170 147430 274226
rect 147498 274170 147554 274226
rect 147622 274170 147678 274226
rect 147250 274046 147306 274102
rect 147374 274046 147430 274102
rect 147498 274046 147554 274102
rect 147622 274046 147678 274102
rect 147250 273922 147306 273978
rect 147374 273922 147430 273978
rect 147498 273922 147554 273978
rect 147622 273922 147678 273978
rect 147250 256294 147306 256350
rect 147374 256294 147430 256350
rect 147498 256294 147554 256350
rect 147622 256294 147678 256350
rect 147250 256170 147306 256226
rect 147374 256170 147430 256226
rect 147498 256170 147554 256226
rect 147622 256170 147678 256226
rect 147250 256046 147306 256102
rect 147374 256046 147430 256102
rect 147498 256046 147554 256102
rect 147622 256046 147678 256102
rect 147250 255922 147306 255978
rect 147374 255922 147430 255978
rect 147498 255922 147554 255978
rect 147622 255922 147678 255978
rect 147250 238294 147306 238350
rect 147374 238294 147430 238350
rect 147498 238294 147554 238350
rect 147622 238294 147678 238350
rect 147250 238170 147306 238226
rect 147374 238170 147430 238226
rect 147498 238170 147554 238226
rect 147622 238170 147678 238226
rect 147250 238046 147306 238102
rect 147374 238046 147430 238102
rect 147498 238046 147554 238102
rect 147622 238046 147678 238102
rect 147250 237922 147306 237978
rect 147374 237922 147430 237978
rect 147498 237922 147554 237978
rect 147622 237922 147678 237978
rect 132970 226294 133026 226350
rect 133094 226294 133150 226350
rect 133218 226294 133274 226350
rect 133342 226294 133398 226350
rect 132970 226170 133026 226226
rect 133094 226170 133150 226226
rect 133218 226170 133274 226226
rect 133342 226170 133398 226226
rect 132970 226046 133026 226102
rect 133094 226046 133150 226102
rect 133218 226046 133274 226102
rect 133342 226046 133398 226102
rect 132970 225922 133026 225978
rect 133094 225922 133150 225978
rect 133218 225922 133274 225978
rect 133342 225922 133398 225978
rect 141318 226294 141374 226350
rect 141442 226294 141498 226350
rect 141318 226170 141374 226226
rect 141442 226170 141498 226226
rect 141318 226046 141374 226102
rect 141442 226046 141498 226102
rect 141318 225922 141374 225978
rect 141442 225922 141498 225978
rect 147250 220294 147306 220350
rect 147374 220294 147430 220350
rect 147498 220294 147554 220350
rect 147622 220294 147678 220350
rect 147250 220170 147306 220226
rect 147374 220170 147430 220226
rect 147498 220170 147554 220226
rect 147622 220170 147678 220226
rect 147250 220046 147306 220102
rect 147374 220046 147430 220102
rect 147498 220046 147554 220102
rect 147622 220046 147678 220102
rect 147250 219922 147306 219978
rect 147374 219922 147430 219978
rect 147498 219922 147554 219978
rect 147622 219922 147678 219978
rect 150970 598116 151026 598172
rect 151094 598116 151150 598172
rect 151218 598116 151274 598172
rect 151342 598116 151398 598172
rect 150970 597992 151026 598048
rect 151094 597992 151150 598048
rect 151218 597992 151274 598048
rect 151342 597992 151398 598048
rect 150970 597868 151026 597924
rect 151094 597868 151150 597924
rect 151218 597868 151274 597924
rect 151342 597868 151398 597924
rect 150970 597744 151026 597800
rect 151094 597744 151150 597800
rect 151218 597744 151274 597800
rect 151342 597744 151398 597800
rect 150970 586294 151026 586350
rect 151094 586294 151150 586350
rect 151218 586294 151274 586350
rect 151342 586294 151398 586350
rect 150970 586170 151026 586226
rect 151094 586170 151150 586226
rect 151218 586170 151274 586226
rect 151342 586170 151398 586226
rect 150970 586046 151026 586102
rect 151094 586046 151150 586102
rect 151218 586046 151274 586102
rect 151342 586046 151398 586102
rect 150970 585922 151026 585978
rect 151094 585922 151150 585978
rect 151218 585922 151274 585978
rect 151342 585922 151398 585978
rect 150970 568294 151026 568350
rect 151094 568294 151150 568350
rect 151218 568294 151274 568350
rect 151342 568294 151398 568350
rect 150970 568170 151026 568226
rect 151094 568170 151150 568226
rect 151218 568170 151274 568226
rect 151342 568170 151398 568226
rect 150970 568046 151026 568102
rect 151094 568046 151150 568102
rect 151218 568046 151274 568102
rect 151342 568046 151398 568102
rect 150970 567922 151026 567978
rect 151094 567922 151150 567978
rect 151218 567922 151274 567978
rect 151342 567922 151398 567978
rect 150970 550294 151026 550350
rect 151094 550294 151150 550350
rect 151218 550294 151274 550350
rect 151342 550294 151398 550350
rect 150970 550170 151026 550226
rect 151094 550170 151150 550226
rect 151218 550170 151274 550226
rect 151342 550170 151398 550226
rect 150970 550046 151026 550102
rect 151094 550046 151150 550102
rect 151218 550046 151274 550102
rect 151342 550046 151398 550102
rect 150970 549922 151026 549978
rect 151094 549922 151150 549978
rect 151218 549922 151274 549978
rect 151342 549922 151398 549978
rect 150970 532294 151026 532350
rect 151094 532294 151150 532350
rect 151218 532294 151274 532350
rect 151342 532294 151398 532350
rect 150970 532170 151026 532226
rect 151094 532170 151150 532226
rect 151218 532170 151274 532226
rect 151342 532170 151398 532226
rect 150970 532046 151026 532102
rect 151094 532046 151150 532102
rect 151218 532046 151274 532102
rect 151342 532046 151398 532102
rect 150970 531922 151026 531978
rect 151094 531922 151150 531978
rect 151218 531922 151274 531978
rect 151342 531922 151398 531978
rect 150970 514294 151026 514350
rect 151094 514294 151150 514350
rect 151218 514294 151274 514350
rect 151342 514294 151398 514350
rect 150970 514170 151026 514226
rect 151094 514170 151150 514226
rect 151218 514170 151274 514226
rect 151342 514170 151398 514226
rect 150970 514046 151026 514102
rect 151094 514046 151150 514102
rect 151218 514046 151274 514102
rect 151342 514046 151398 514102
rect 150970 513922 151026 513978
rect 151094 513922 151150 513978
rect 151218 513922 151274 513978
rect 151342 513922 151398 513978
rect 150970 496294 151026 496350
rect 151094 496294 151150 496350
rect 151218 496294 151274 496350
rect 151342 496294 151398 496350
rect 150970 496170 151026 496226
rect 151094 496170 151150 496226
rect 151218 496170 151274 496226
rect 151342 496170 151398 496226
rect 150970 496046 151026 496102
rect 151094 496046 151150 496102
rect 151218 496046 151274 496102
rect 151342 496046 151398 496102
rect 150970 495922 151026 495978
rect 151094 495922 151150 495978
rect 151218 495922 151274 495978
rect 151342 495922 151398 495978
rect 150970 478294 151026 478350
rect 151094 478294 151150 478350
rect 151218 478294 151274 478350
rect 151342 478294 151398 478350
rect 150970 478170 151026 478226
rect 151094 478170 151150 478226
rect 151218 478170 151274 478226
rect 151342 478170 151398 478226
rect 150970 478046 151026 478102
rect 151094 478046 151150 478102
rect 151218 478046 151274 478102
rect 151342 478046 151398 478102
rect 150970 477922 151026 477978
rect 151094 477922 151150 477978
rect 151218 477922 151274 477978
rect 151342 477922 151398 477978
rect 150970 460294 151026 460350
rect 151094 460294 151150 460350
rect 151218 460294 151274 460350
rect 151342 460294 151398 460350
rect 150970 460170 151026 460226
rect 151094 460170 151150 460226
rect 151218 460170 151274 460226
rect 151342 460170 151398 460226
rect 150970 460046 151026 460102
rect 151094 460046 151150 460102
rect 151218 460046 151274 460102
rect 151342 460046 151398 460102
rect 150970 459922 151026 459978
rect 151094 459922 151150 459978
rect 151218 459922 151274 459978
rect 151342 459922 151398 459978
rect 150970 442294 151026 442350
rect 151094 442294 151150 442350
rect 151218 442294 151274 442350
rect 151342 442294 151398 442350
rect 150970 442170 151026 442226
rect 151094 442170 151150 442226
rect 151218 442170 151274 442226
rect 151342 442170 151398 442226
rect 150970 442046 151026 442102
rect 151094 442046 151150 442102
rect 151218 442046 151274 442102
rect 151342 442046 151398 442102
rect 150970 441922 151026 441978
rect 151094 441922 151150 441978
rect 151218 441922 151274 441978
rect 151342 441922 151398 441978
rect 150970 424294 151026 424350
rect 151094 424294 151150 424350
rect 151218 424294 151274 424350
rect 151342 424294 151398 424350
rect 150970 424170 151026 424226
rect 151094 424170 151150 424226
rect 151218 424170 151274 424226
rect 151342 424170 151398 424226
rect 150970 424046 151026 424102
rect 151094 424046 151150 424102
rect 151218 424046 151274 424102
rect 151342 424046 151398 424102
rect 150970 423922 151026 423978
rect 151094 423922 151150 423978
rect 151218 423922 151274 423978
rect 151342 423922 151398 423978
rect 150970 406294 151026 406350
rect 151094 406294 151150 406350
rect 151218 406294 151274 406350
rect 151342 406294 151398 406350
rect 150970 406170 151026 406226
rect 151094 406170 151150 406226
rect 151218 406170 151274 406226
rect 151342 406170 151398 406226
rect 150970 406046 151026 406102
rect 151094 406046 151150 406102
rect 151218 406046 151274 406102
rect 151342 406046 151398 406102
rect 150970 405922 151026 405978
rect 151094 405922 151150 405978
rect 151218 405922 151274 405978
rect 151342 405922 151398 405978
rect 150970 388294 151026 388350
rect 151094 388294 151150 388350
rect 151218 388294 151274 388350
rect 151342 388294 151398 388350
rect 150970 388170 151026 388226
rect 151094 388170 151150 388226
rect 151218 388170 151274 388226
rect 151342 388170 151398 388226
rect 150970 388046 151026 388102
rect 151094 388046 151150 388102
rect 151218 388046 151274 388102
rect 151342 388046 151398 388102
rect 150970 387922 151026 387978
rect 151094 387922 151150 387978
rect 151218 387922 151274 387978
rect 151342 387922 151398 387978
rect 150970 370294 151026 370350
rect 151094 370294 151150 370350
rect 151218 370294 151274 370350
rect 151342 370294 151398 370350
rect 150970 370170 151026 370226
rect 151094 370170 151150 370226
rect 151218 370170 151274 370226
rect 151342 370170 151398 370226
rect 150970 370046 151026 370102
rect 151094 370046 151150 370102
rect 151218 370046 151274 370102
rect 151342 370046 151398 370102
rect 150970 369922 151026 369978
rect 151094 369922 151150 369978
rect 151218 369922 151274 369978
rect 151342 369922 151398 369978
rect 150970 352294 151026 352350
rect 151094 352294 151150 352350
rect 151218 352294 151274 352350
rect 151342 352294 151398 352350
rect 150970 352170 151026 352226
rect 151094 352170 151150 352226
rect 151218 352170 151274 352226
rect 151342 352170 151398 352226
rect 150970 352046 151026 352102
rect 151094 352046 151150 352102
rect 151218 352046 151274 352102
rect 151342 352046 151398 352102
rect 150970 351922 151026 351978
rect 151094 351922 151150 351978
rect 151218 351922 151274 351978
rect 151342 351922 151398 351978
rect 150970 334294 151026 334350
rect 151094 334294 151150 334350
rect 151218 334294 151274 334350
rect 151342 334294 151398 334350
rect 150970 334170 151026 334226
rect 151094 334170 151150 334226
rect 151218 334170 151274 334226
rect 151342 334170 151398 334226
rect 150970 334046 151026 334102
rect 151094 334046 151150 334102
rect 151218 334046 151274 334102
rect 151342 334046 151398 334102
rect 150970 333922 151026 333978
rect 151094 333922 151150 333978
rect 151218 333922 151274 333978
rect 151342 333922 151398 333978
rect 150970 316294 151026 316350
rect 151094 316294 151150 316350
rect 151218 316294 151274 316350
rect 151342 316294 151398 316350
rect 150970 316170 151026 316226
rect 151094 316170 151150 316226
rect 151218 316170 151274 316226
rect 151342 316170 151398 316226
rect 150970 316046 151026 316102
rect 151094 316046 151150 316102
rect 151218 316046 151274 316102
rect 151342 316046 151398 316102
rect 150970 315922 151026 315978
rect 151094 315922 151150 315978
rect 151218 315922 151274 315978
rect 151342 315922 151398 315978
rect 150970 298294 151026 298350
rect 151094 298294 151150 298350
rect 151218 298294 151274 298350
rect 151342 298294 151398 298350
rect 150970 298170 151026 298226
rect 151094 298170 151150 298226
rect 151218 298170 151274 298226
rect 151342 298170 151398 298226
rect 150970 298046 151026 298102
rect 151094 298046 151150 298102
rect 151218 298046 151274 298102
rect 151342 298046 151398 298102
rect 150970 297922 151026 297978
rect 151094 297922 151150 297978
rect 151218 297922 151274 297978
rect 151342 297922 151398 297978
rect 150970 280294 151026 280350
rect 151094 280294 151150 280350
rect 151218 280294 151274 280350
rect 151342 280294 151398 280350
rect 150970 280170 151026 280226
rect 151094 280170 151150 280226
rect 151218 280170 151274 280226
rect 151342 280170 151398 280226
rect 150970 280046 151026 280102
rect 151094 280046 151150 280102
rect 151218 280046 151274 280102
rect 151342 280046 151398 280102
rect 150970 279922 151026 279978
rect 151094 279922 151150 279978
rect 151218 279922 151274 279978
rect 151342 279922 151398 279978
rect 150970 262294 151026 262350
rect 151094 262294 151150 262350
rect 151218 262294 151274 262350
rect 151342 262294 151398 262350
rect 150970 262170 151026 262226
rect 151094 262170 151150 262226
rect 151218 262170 151274 262226
rect 151342 262170 151398 262226
rect 150970 262046 151026 262102
rect 151094 262046 151150 262102
rect 151218 262046 151274 262102
rect 151342 262046 151398 262102
rect 150970 261922 151026 261978
rect 151094 261922 151150 261978
rect 151218 261922 151274 261978
rect 151342 261922 151398 261978
rect 150970 244294 151026 244350
rect 151094 244294 151150 244350
rect 151218 244294 151274 244350
rect 151342 244294 151398 244350
rect 150970 244170 151026 244226
rect 151094 244170 151150 244226
rect 151218 244170 151274 244226
rect 151342 244170 151398 244226
rect 150970 244046 151026 244102
rect 151094 244046 151150 244102
rect 151218 244046 151274 244102
rect 151342 244046 151398 244102
rect 150970 243922 151026 243978
rect 151094 243922 151150 243978
rect 151218 243922 151274 243978
rect 151342 243922 151398 243978
rect 168970 598116 169026 598172
rect 169094 598116 169150 598172
rect 169218 598116 169274 598172
rect 169342 598116 169398 598172
rect 168970 597992 169026 598048
rect 169094 597992 169150 598048
rect 169218 597992 169274 598048
rect 169342 597992 169398 598048
rect 168970 597868 169026 597924
rect 169094 597868 169150 597924
rect 169218 597868 169274 597924
rect 169342 597868 169398 597924
rect 168970 597744 169026 597800
rect 169094 597744 169150 597800
rect 169218 597744 169274 597800
rect 169342 597744 169398 597800
rect 168970 586294 169026 586350
rect 169094 586294 169150 586350
rect 169218 586294 169274 586350
rect 169342 586294 169398 586350
rect 168970 586170 169026 586226
rect 169094 586170 169150 586226
rect 169218 586170 169274 586226
rect 169342 586170 169398 586226
rect 168970 586046 169026 586102
rect 169094 586046 169150 586102
rect 169218 586046 169274 586102
rect 169342 586046 169398 586102
rect 168970 585922 169026 585978
rect 169094 585922 169150 585978
rect 169218 585922 169274 585978
rect 169342 585922 169398 585978
rect 168970 568294 169026 568350
rect 169094 568294 169150 568350
rect 169218 568294 169274 568350
rect 169342 568294 169398 568350
rect 168970 568170 169026 568226
rect 169094 568170 169150 568226
rect 169218 568170 169274 568226
rect 169342 568170 169398 568226
rect 168970 568046 169026 568102
rect 169094 568046 169150 568102
rect 169218 568046 169274 568102
rect 169342 568046 169398 568102
rect 168970 567922 169026 567978
rect 169094 567922 169150 567978
rect 169218 567922 169274 567978
rect 169342 567922 169398 567978
rect 168970 550294 169026 550350
rect 169094 550294 169150 550350
rect 169218 550294 169274 550350
rect 169342 550294 169398 550350
rect 168970 550170 169026 550226
rect 169094 550170 169150 550226
rect 169218 550170 169274 550226
rect 169342 550170 169398 550226
rect 168970 550046 169026 550102
rect 169094 550046 169150 550102
rect 169218 550046 169274 550102
rect 169342 550046 169398 550102
rect 168970 549922 169026 549978
rect 169094 549922 169150 549978
rect 169218 549922 169274 549978
rect 169342 549922 169398 549978
rect 168970 532294 169026 532350
rect 169094 532294 169150 532350
rect 169218 532294 169274 532350
rect 169342 532294 169398 532350
rect 168970 532170 169026 532226
rect 169094 532170 169150 532226
rect 169218 532170 169274 532226
rect 169342 532170 169398 532226
rect 168970 532046 169026 532102
rect 169094 532046 169150 532102
rect 169218 532046 169274 532102
rect 169342 532046 169398 532102
rect 168970 531922 169026 531978
rect 169094 531922 169150 531978
rect 169218 531922 169274 531978
rect 169342 531922 169398 531978
rect 168970 514294 169026 514350
rect 169094 514294 169150 514350
rect 169218 514294 169274 514350
rect 169342 514294 169398 514350
rect 168970 514170 169026 514226
rect 169094 514170 169150 514226
rect 169218 514170 169274 514226
rect 169342 514170 169398 514226
rect 168970 514046 169026 514102
rect 169094 514046 169150 514102
rect 169218 514046 169274 514102
rect 169342 514046 169398 514102
rect 168970 513922 169026 513978
rect 169094 513922 169150 513978
rect 169218 513922 169274 513978
rect 169342 513922 169398 513978
rect 168970 496294 169026 496350
rect 169094 496294 169150 496350
rect 169218 496294 169274 496350
rect 169342 496294 169398 496350
rect 168970 496170 169026 496226
rect 169094 496170 169150 496226
rect 169218 496170 169274 496226
rect 169342 496170 169398 496226
rect 168970 496046 169026 496102
rect 169094 496046 169150 496102
rect 169218 496046 169274 496102
rect 169342 496046 169398 496102
rect 168970 495922 169026 495978
rect 169094 495922 169150 495978
rect 169218 495922 169274 495978
rect 169342 495922 169398 495978
rect 168970 478294 169026 478350
rect 169094 478294 169150 478350
rect 169218 478294 169274 478350
rect 169342 478294 169398 478350
rect 168970 478170 169026 478226
rect 169094 478170 169150 478226
rect 169218 478170 169274 478226
rect 169342 478170 169398 478226
rect 168970 478046 169026 478102
rect 169094 478046 169150 478102
rect 169218 478046 169274 478102
rect 169342 478046 169398 478102
rect 168970 477922 169026 477978
rect 169094 477922 169150 477978
rect 169218 477922 169274 477978
rect 169342 477922 169398 477978
rect 168970 460294 169026 460350
rect 169094 460294 169150 460350
rect 169218 460294 169274 460350
rect 169342 460294 169398 460350
rect 168970 460170 169026 460226
rect 169094 460170 169150 460226
rect 169218 460170 169274 460226
rect 169342 460170 169398 460226
rect 168970 460046 169026 460102
rect 169094 460046 169150 460102
rect 169218 460046 169274 460102
rect 169342 460046 169398 460102
rect 168970 459922 169026 459978
rect 169094 459922 169150 459978
rect 169218 459922 169274 459978
rect 169342 459922 169398 459978
rect 168970 442294 169026 442350
rect 169094 442294 169150 442350
rect 169218 442294 169274 442350
rect 169342 442294 169398 442350
rect 168970 442170 169026 442226
rect 169094 442170 169150 442226
rect 169218 442170 169274 442226
rect 169342 442170 169398 442226
rect 168970 442046 169026 442102
rect 169094 442046 169150 442102
rect 169218 442046 169274 442102
rect 169342 442046 169398 442102
rect 168970 441922 169026 441978
rect 169094 441922 169150 441978
rect 169218 441922 169274 441978
rect 169342 441922 169398 441978
rect 168970 424294 169026 424350
rect 169094 424294 169150 424350
rect 169218 424294 169274 424350
rect 169342 424294 169398 424350
rect 168970 424170 169026 424226
rect 169094 424170 169150 424226
rect 169218 424170 169274 424226
rect 169342 424170 169398 424226
rect 168970 424046 169026 424102
rect 169094 424046 169150 424102
rect 169218 424046 169274 424102
rect 169342 424046 169398 424102
rect 168970 423922 169026 423978
rect 169094 423922 169150 423978
rect 169218 423922 169274 423978
rect 169342 423922 169398 423978
rect 168970 406294 169026 406350
rect 169094 406294 169150 406350
rect 169218 406294 169274 406350
rect 169342 406294 169398 406350
rect 168970 406170 169026 406226
rect 169094 406170 169150 406226
rect 169218 406170 169274 406226
rect 169342 406170 169398 406226
rect 168970 406046 169026 406102
rect 169094 406046 169150 406102
rect 169218 406046 169274 406102
rect 169342 406046 169398 406102
rect 168970 405922 169026 405978
rect 169094 405922 169150 405978
rect 169218 405922 169274 405978
rect 169342 405922 169398 405978
rect 168970 388294 169026 388350
rect 169094 388294 169150 388350
rect 169218 388294 169274 388350
rect 169342 388294 169398 388350
rect 168970 388170 169026 388226
rect 169094 388170 169150 388226
rect 169218 388170 169274 388226
rect 169342 388170 169398 388226
rect 168970 388046 169026 388102
rect 169094 388046 169150 388102
rect 169218 388046 169274 388102
rect 169342 388046 169398 388102
rect 168970 387922 169026 387978
rect 169094 387922 169150 387978
rect 169218 387922 169274 387978
rect 169342 387922 169398 387978
rect 168970 370294 169026 370350
rect 169094 370294 169150 370350
rect 169218 370294 169274 370350
rect 169342 370294 169398 370350
rect 168970 370170 169026 370226
rect 169094 370170 169150 370226
rect 169218 370170 169274 370226
rect 169342 370170 169398 370226
rect 168970 370046 169026 370102
rect 169094 370046 169150 370102
rect 169218 370046 169274 370102
rect 169342 370046 169398 370102
rect 168970 369922 169026 369978
rect 169094 369922 169150 369978
rect 169218 369922 169274 369978
rect 169342 369922 169398 369978
rect 168970 352294 169026 352350
rect 169094 352294 169150 352350
rect 169218 352294 169274 352350
rect 169342 352294 169398 352350
rect 168970 352170 169026 352226
rect 169094 352170 169150 352226
rect 169218 352170 169274 352226
rect 169342 352170 169398 352226
rect 168970 352046 169026 352102
rect 169094 352046 169150 352102
rect 169218 352046 169274 352102
rect 169342 352046 169398 352102
rect 168970 351922 169026 351978
rect 169094 351922 169150 351978
rect 169218 351922 169274 351978
rect 169342 351922 169398 351978
rect 168970 334294 169026 334350
rect 169094 334294 169150 334350
rect 169218 334294 169274 334350
rect 169342 334294 169398 334350
rect 168970 334170 169026 334226
rect 169094 334170 169150 334226
rect 169218 334170 169274 334226
rect 169342 334170 169398 334226
rect 168970 334046 169026 334102
rect 169094 334046 169150 334102
rect 169218 334046 169274 334102
rect 169342 334046 169398 334102
rect 168970 333922 169026 333978
rect 169094 333922 169150 333978
rect 169218 333922 169274 333978
rect 169342 333922 169398 333978
rect 168970 316294 169026 316350
rect 169094 316294 169150 316350
rect 169218 316294 169274 316350
rect 169342 316294 169398 316350
rect 168970 316170 169026 316226
rect 169094 316170 169150 316226
rect 169218 316170 169274 316226
rect 169342 316170 169398 316226
rect 168970 316046 169026 316102
rect 169094 316046 169150 316102
rect 169218 316046 169274 316102
rect 169342 316046 169398 316102
rect 168970 315922 169026 315978
rect 169094 315922 169150 315978
rect 169218 315922 169274 315978
rect 169342 315922 169398 315978
rect 168970 298294 169026 298350
rect 169094 298294 169150 298350
rect 169218 298294 169274 298350
rect 169342 298294 169398 298350
rect 168970 298170 169026 298226
rect 169094 298170 169150 298226
rect 169218 298170 169274 298226
rect 169342 298170 169398 298226
rect 168970 298046 169026 298102
rect 169094 298046 169150 298102
rect 169218 298046 169274 298102
rect 169342 298046 169398 298102
rect 168970 297922 169026 297978
rect 169094 297922 169150 297978
rect 169218 297922 169274 297978
rect 169342 297922 169398 297978
rect 168970 280294 169026 280350
rect 169094 280294 169150 280350
rect 169218 280294 169274 280350
rect 169342 280294 169398 280350
rect 168970 280170 169026 280226
rect 169094 280170 169150 280226
rect 169218 280170 169274 280226
rect 169342 280170 169398 280226
rect 168970 280046 169026 280102
rect 169094 280046 169150 280102
rect 169218 280046 169274 280102
rect 169342 280046 169398 280102
rect 168970 279922 169026 279978
rect 169094 279922 169150 279978
rect 169218 279922 169274 279978
rect 169342 279922 169398 279978
rect 168970 262294 169026 262350
rect 169094 262294 169150 262350
rect 169218 262294 169274 262350
rect 169342 262294 169398 262350
rect 168970 262170 169026 262226
rect 169094 262170 169150 262226
rect 169218 262170 169274 262226
rect 169342 262170 169398 262226
rect 168970 262046 169026 262102
rect 169094 262046 169150 262102
rect 169218 262046 169274 262102
rect 169342 262046 169398 262102
rect 168970 261922 169026 261978
rect 169094 261922 169150 261978
rect 169218 261922 169274 261978
rect 169342 261922 169398 261978
rect 168970 244294 169026 244350
rect 169094 244294 169150 244350
rect 169218 244294 169274 244350
rect 169342 244294 169398 244350
rect 168970 244170 169026 244226
rect 169094 244170 169150 244226
rect 169218 244170 169274 244226
rect 169342 244170 169398 244226
rect 168970 244046 169026 244102
rect 169094 244046 169150 244102
rect 169218 244046 169274 244102
rect 169342 244046 169398 244102
rect 168970 243922 169026 243978
rect 169094 243922 169150 243978
rect 169218 243922 169274 243978
rect 169342 243922 169398 243978
rect 150970 226294 151026 226350
rect 151094 226294 151150 226350
rect 151218 226294 151274 226350
rect 151342 226294 151398 226350
rect 150970 226170 151026 226226
rect 151094 226170 151150 226226
rect 151218 226170 151274 226226
rect 151342 226170 151398 226226
rect 150970 226046 151026 226102
rect 151094 226046 151150 226102
rect 151218 226046 151274 226102
rect 151342 226046 151398 226102
rect 150970 225922 151026 225978
rect 151094 225922 151150 225978
rect 151218 225922 151274 225978
rect 151342 225922 151398 225978
rect 165250 238294 165306 238350
rect 165374 238294 165430 238350
rect 165498 238294 165554 238350
rect 165622 238294 165678 238350
rect 165250 238170 165306 238226
rect 165374 238170 165430 238226
rect 165498 238170 165554 238226
rect 165622 238170 165678 238226
rect 165250 238046 165306 238102
rect 165374 238046 165430 238102
rect 165498 238046 165554 238102
rect 165622 238046 165678 238102
rect 165250 237922 165306 237978
rect 165374 237922 165430 237978
rect 165498 237922 165554 237978
rect 165622 237922 165678 237978
rect 156678 220294 156734 220350
rect 156802 220294 156858 220350
rect 156678 220170 156734 220226
rect 156802 220170 156858 220226
rect 156678 220046 156734 220102
rect 156802 220046 156858 220102
rect 156678 219922 156734 219978
rect 156802 219922 156858 219978
rect 165250 220294 165306 220350
rect 165374 220294 165430 220350
rect 165498 220294 165554 220350
rect 165622 220294 165678 220350
rect 165250 220170 165306 220226
rect 165374 220170 165430 220226
rect 165498 220170 165554 220226
rect 165622 220170 165678 220226
rect 165250 220046 165306 220102
rect 165374 220046 165430 220102
rect 165498 220046 165554 220102
rect 165622 220046 165678 220102
rect 165250 219922 165306 219978
rect 165374 219922 165430 219978
rect 165498 219922 165554 219978
rect 165622 219922 165678 219978
rect 183250 597156 183306 597212
rect 183374 597156 183430 597212
rect 183498 597156 183554 597212
rect 183622 597156 183678 597212
rect 183250 597032 183306 597088
rect 183374 597032 183430 597088
rect 183498 597032 183554 597088
rect 183622 597032 183678 597088
rect 183250 596908 183306 596964
rect 183374 596908 183430 596964
rect 183498 596908 183554 596964
rect 183622 596908 183678 596964
rect 183250 596784 183306 596840
rect 183374 596784 183430 596840
rect 183498 596784 183554 596840
rect 183622 596784 183678 596840
rect 183250 580294 183306 580350
rect 183374 580294 183430 580350
rect 183498 580294 183554 580350
rect 183622 580294 183678 580350
rect 183250 580170 183306 580226
rect 183374 580170 183430 580226
rect 183498 580170 183554 580226
rect 183622 580170 183678 580226
rect 183250 580046 183306 580102
rect 183374 580046 183430 580102
rect 183498 580046 183554 580102
rect 183622 580046 183678 580102
rect 183250 579922 183306 579978
rect 183374 579922 183430 579978
rect 183498 579922 183554 579978
rect 183622 579922 183678 579978
rect 183250 562294 183306 562350
rect 183374 562294 183430 562350
rect 183498 562294 183554 562350
rect 183622 562294 183678 562350
rect 183250 562170 183306 562226
rect 183374 562170 183430 562226
rect 183498 562170 183554 562226
rect 183622 562170 183678 562226
rect 183250 562046 183306 562102
rect 183374 562046 183430 562102
rect 183498 562046 183554 562102
rect 183622 562046 183678 562102
rect 183250 561922 183306 561978
rect 183374 561922 183430 561978
rect 183498 561922 183554 561978
rect 183622 561922 183678 561978
rect 183250 544294 183306 544350
rect 183374 544294 183430 544350
rect 183498 544294 183554 544350
rect 183622 544294 183678 544350
rect 183250 544170 183306 544226
rect 183374 544170 183430 544226
rect 183498 544170 183554 544226
rect 183622 544170 183678 544226
rect 183250 544046 183306 544102
rect 183374 544046 183430 544102
rect 183498 544046 183554 544102
rect 183622 544046 183678 544102
rect 183250 543922 183306 543978
rect 183374 543922 183430 543978
rect 183498 543922 183554 543978
rect 183622 543922 183678 543978
rect 183250 526294 183306 526350
rect 183374 526294 183430 526350
rect 183498 526294 183554 526350
rect 183622 526294 183678 526350
rect 183250 526170 183306 526226
rect 183374 526170 183430 526226
rect 183498 526170 183554 526226
rect 183622 526170 183678 526226
rect 183250 526046 183306 526102
rect 183374 526046 183430 526102
rect 183498 526046 183554 526102
rect 183622 526046 183678 526102
rect 183250 525922 183306 525978
rect 183374 525922 183430 525978
rect 183498 525922 183554 525978
rect 183622 525922 183678 525978
rect 183250 508294 183306 508350
rect 183374 508294 183430 508350
rect 183498 508294 183554 508350
rect 183622 508294 183678 508350
rect 183250 508170 183306 508226
rect 183374 508170 183430 508226
rect 183498 508170 183554 508226
rect 183622 508170 183678 508226
rect 183250 508046 183306 508102
rect 183374 508046 183430 508102
rect 183498 508046 183554 508102
rect 183622 508046 183678 508102
rect 183250 507922 183306 507978
rect 183374 507922 183430 507978
rect 183498 507922 183554 507978
rect 183622 507922 183678 507978
rect 183250 490294 183306 490350
rect 183374 490294 183430 490350
rect 183498 490294 183554 490350
rect 183622 490294 183678 490350
rect 183250 490170 183306 490226
rect 183374 490170 183430 490226
rect 183498 490170 183554 490226
rect 183622 490170 183678 490226
rect 183250 490046 183306 490102
rect 183374 490046 183430 490102
rect 183498 490046 183554 490102
rect 183622 490046 183678 490102
rect 183250 489922 183306 489978
rect 183374 489922 183430 489978
rect 183498 489922 183554 489978
rect 183622 489922 183678 489978
rect 183250 472294 183306 472350
rect 183374 472294 183430 472350
rect 183498 472294 183554 472350
rect 183622 472294 183678 472350
rect 183250 472170 183306 472226
rect 183374 472170 183430 472226
rect 183498 472170 183554 472226
rect 183622 472170 183678 472226
rect 183250 472046 183306 472102
rect 183374 472046 183430 472102
rect 183498 472046 183554 472102
rect 183622 472046 183678 472102
rect 183250 471922 183306 471978
rect 183374 471922 183430 471978
rect 183498 471922 183554 471978
rect 183622 471922 183678 471978
rect 183250 454294 183306 454350
rect 183374 454294 183430 454350
rect 183498 454294 183554 454350
rect 183622 454294 183678 454350
rect 183250 454170 183306 454226
rect 183374 454170 183430 454226
rect 183498 454170 183554 454226
rect 183622 454170 183678 454226
rect 183250 454046 183306 454102
rect 183374 454046 183430 454102
rect 183498 454046 183554 454102
rect 183622 454046 183678 454102
rect 183250 453922 183306 453978
rect 183374 453922 183430 453978
rect 183498 453922 183554 453978
rect 183622 453922 183678 453978
rect 183250 436294 183306 436350
rect 183374 436294 183430 436350
rect 183498 436294 183554 436350
rect 183622 436294 183678 436350
rect 183250 436170 183306 436226
rect 183374 436170 183430 436226
rect 183498 436170 183554 436226
rect 183622 436170 183678 436226
rect 183250 436046 183306 436102
rect 183374 436046 183430 436102
rect 183498 436046 183554 436102
rect 183622 436046 183678 436102
rect 183250 435922 183306 435978
rect 183374 435922 183430 435978
rect 183498 435922 183554 435978
rect 183622 435922 183678 435978
rect 183250 418294 183306 418350
rect 183374 418294 183430 418350
rect 183498 418294 183554 418350
rect 183622 418294 183678 418350
rect 183250 418170 183306 418226
rect 183374 418170 183430 418226
rect 183498 418170 183554 418226
rect 183622 418170 183678 418226
rect 183250 418046 183306 418102
rect 183374 418046 183430 418102
rect 183498 418046 183554 418102
rect 183622 418046 183678 418102
rect 183250 417922 183306 417978
rect 183374 417922 183430 417978
rect 183498 417922 183554 417978
rect 183622 417922 183678 417978
rect 183250 400294 183306 400350
rect 183374 400294 183430 400350
rect 183498 400294 183554 400350
rect 183622 400294 183678 400350
rect 183250 400170 183306 400226
rect 183374 400170 183430 400226
rect 183498 400170 183554 400226
rect 183622 400170 183678 400226
rect 183250 400046 183306 400102
rect 183374 400046 183430 400102
rect 183498 400046 183554 400102
rect 183622 400046 183678 400102
rect 183250 399922 183306 399978
rect 183374 399922 183430 399978
rect 183498 399922 183554 399978
rect 183622 399922 183678 399978
rect 183250 382294 183306 382350
rect 183374 382294 183430 382350
rect 183498 382294 183554 382350
rect 183622 382294 183678 382350
rect 183250 382170 183306 382226
rect 183374 382170 183430 382226
rect 183498 382170 183554 382226
rect 183622 382170 183678 382226
rect 183250 382046 183306 382102
rect 183374 382046 183430 382102
rect 183498 382046 183554 382102
rect 183622 382046 183678 382102
rect 183250 381922 183306 381978
rect 183374 381922 183430 381978
rect 183498 381922 183554 381978
rect 183622 381922 183678 381978
rect 183250 364294 183306 364350
rect 183374 364294 183430 364350
rect 183498 364294 183554 364350
rect 183622 364294 183678 364350
rect 183250 364170 183306 364226
rect 183374 364170 183430 364226
rect 183498 364170 183554 364226
rect 183622 364170 183678 364226
rect 183250 364046 183306 364102
rect 183374 364046 183430 364102
rect 183498 364046 183554 364102
rect 183622 364046 183678 364102
rect 183250 363922 183306 363978
rect 183374 363922 183430 363978
rect 183498 363922 183554 363978
rect 183622 363922 183678 363978
rect 183250 346294 183306 346350
rect 183374 346294 183430 346350
rect 183498 346294 183554 346350
rect 183622 346294 183678 346350
rect 183250 346170 183306 346226
rect 183374 346170 183430 346226
rect 183498 346170 183554 346226
rect 183622 346170 183678 346226
rect 183250 346046 183306 346102
rect 183374 346046 183430 346102
rect 183498 346046 183554 346102
rect 183622 346046 183678 346102
rect 183250 345922 183306 345978
rect 183374 345922 183430 345978
rect 183498 345922 183554 345978
rect 183622 345922 183678 345978
rect 183250 328294 183306 328350
rect 183374 328294 183430 328350
rect 183498 328294 183554 328350
rect 183622 328294 183678 328350
rect 183250 328170 183306 328226
rect 183374 328170 183430 328226
rect 183498 328170 183554 328226
rect 183622 328170 183678 328226
rect 183250 328046 183306 328102
rect 183374 328046 183430 328102
rect 183498 328046 183554 328102
rect 183622 328046 183678 328102
rect 183250 327922 183306 327978
rect 183374 327922 183430 327978
rect 183498 327922 183554 327978
rect 183622 327922 183678 327978
rect 183250 310294 183306 310350
rect 183374 310294 183430 310350
rect 183498 310294 183554 310350
rect 183622 310294 183678 310350
rect 183250 310170 183306 310226
rect 183374 310170 183430 310226
rect 183498 310170 183554 310226
rect 183622 310170 183678 310226
rect 183250 310046 183306 310102
rect 183374 310046 183430 310102
rect 183498 310046 183554 310102
rect 183622 310046 183678 310102
rect 183250 309922 183306 309978
rect 183374 309922 183430 309978
rect 183498 309922 183554 309978
rect 183622 309922 183678 309978
rect 183250 292294 183306 292350
rect 183374 292294 183430 292350
rect 183498 292294 183554 292350
rect 183622 292294 183678 292350
rect 183250 292170 183306 292226
rect 183374 292170 183430 292226
rect 183498 292170 183554 292226
rect 183622 292170 183678 292226
rect 183250 292046 183306 292102
rect 183374 292046 183430 292102
rect 183498 292046 183554 292102
rect 183622 292046 183678 292102
rect 183250 291922 183306 291978
rect 183374 291922 183430 291978
rect 183498 291922 183554 291978
rect 183622 291922 183678 291978
rect 183250 274294 183306 274350
rect 183374 274294 183430 274350
rect 183498 274294 183554 274350
rect 183622 274294 183678 274350
rect 183250 274170 183306 274226
rect 183374 274170 183430 274226
rect 183498 274170 183554 274226
rect 183622 274170 183678 274226
rect 183250 274046 183306 274102
rect 183374 274046 183430 274102
rect 183498 274046 183554 274102
rect 183622 274046 183678 274102
rect 183250 273922 183306 273978
rect 183374 273922 183430 273978
rect 183498 273922 183554 273978
rect 183622 273922 183678 273978
rect 183250 256294 183306 256350
rect 183374 256294 183430 256350
rect 183498 256294 183554 256350
rect 183622 256294 183678 256350
rect 183250 256170 183306 256226
rect 183374 256170 183430 256226
rect 183498 256170 183554 256226
rect 183622 256170 183678 256226
rect 183250 256046 183306 256102
rect 183374 256046 183430 256102
rect 183498 256046 183554 256102
rect 183622 256046 183678 256102
rect 183250 255922 183306 255978
rect 183374 255922 183430 255978
rect 183498 255922 183554 255978
rect 183622 255922 183678 255978
rect 183250 238294 183306 238350
rect 183374 238294 183430 238350
rect 183498 238294 183554 238350
rect 183622 238294 183678 238350
rect 183250 238170 183306 238226
rect 183374 238170 183430 238226
rect 183498 238170 183554 238226
rect 183622 238170 183678 238226
rect 183250 238046 183306 238102
rect 183374 238046 183430 238102
rect 183498 238046 183554 238102
rect 183622 238046 183678 238102
rect 183250 237922 183306 237978
rect 183374 237922 183430 237978
rect 183498 237922 183554 237978
rect 183622 237922 183678 237978
rect 168970 226294 169026 226350
rect 169094 226294 169150 226350
rect 169218 226294 169274 226350
rect 169342 226294 169398 226350
rect 168970 226170 169026 226226
rect 169094 226170 169150 226226
rect 169218 226170 169274 226226
rect 169342 226170 169398 226226
rect 168970 226046 169026 226102
rect 169094 226046 169150 226102
rect 169218 226046 169274 226102
rect 169342 226046 169398 226102
rect 168970 225922 169026 225978
rect 169094 225922 169150 225978
rect 169218 225922 169274 225978
rect 169342 225922 169398 225978
rect 172038 226294 172094 226350
rect 172162 226294 172218 226350
rect 172038 226170 172094 226226
rect 172162 226170 172218 226226
rect 172038 226046 172094 226102
rect 172162 226046 172218 226102
rect 172038 225922 172094 225978
rect 172162 225922 172218 225978
rect 186970 598116 187026 598172
rect 187094 598116 187150 598172
rect 187218 598116 187274 598172
rect 187342 598116 187398 598172
rect 186970 597992 187026 598048
rect 187094 597992 187150 598048
rect 187218 597992 187274 598048
rect 187342 597992 187398 598048
rect 186970 597868 187026 597924
rect 187094 597868 187150 597924
rect 187218 597868 187274 597924
rect 187342 597868 187398 597924
rect 186970 597744 187026 597800
rect 187094 597744 187150 597800
rect 187218 597744 187274 597800
rect 187342 597744 187398 597800
rect 186970 586294 187026 586350
rect 187094 586294 187150 586350
rect 187218 586294 187274 586350
rect 187342 586294 187398 586350
rect 186970 586170 187026 586226
rect 187094 586170 187150 586226
rect 187218 586170 187274 586226
rect 187342 586170 187398 586226
rect 186970 586046 187026 586102
rect 187094 586046 187150 586102
rect 187218 586046 187274 586102
rect 187342 586046 187398 586102
rect 186970 585922 187026 585978
rect 187094 585922 187150 585978
rect 187218 585922 187274 585978
rect 187342 585922 187398 585978
rect 186970 568294 187026 568350
rect 187094 568294 187150 568350
rect 187218 568294 187274 568350
rect 187342 568294 187398 568350
rect 186970 568170 187026 568226
rect 187094 568170 187150 568226
rect 187218 568170 187274 568226
rect 187342 568170 187398 568226
rect 186970 568046 187026 568102
rect 187094 568046 187150 568102
rect 187218 568046 187274 568102
rect 187342 568046 187398 568102
rect 186970 567922 187026 567978
rect 187094 567922 187150 567978
rect 187218 567922 187274 567978
rect 187342 567922 187398 567978
rect 186970 550294 187026 550350
rect 187094 550294 187150 550350
rect 187218 550294 187274 550350
rect 187342 550294 187398 550350
rect 186970 550170 187026 550226
rect 187094 550170 187150 550226
rect 187218 550170 187274 550226
rect 187342 550170 187398 550226
rect 186970 550046 187026 550102
rect 187094 550046 187150 550102
rect 187218 550046 187274 550102
rect 187342 550046 187398 550102
rect 186970 549922 187026 549978
rect 187094 549922 187150 549978
rect 187218 549922 187274 549978
rect 187342 549922 187398 549978
rect 186970 532294 187026 532350
rect 187094 532294 187150 532350
rect 187218 532294 187274 532350
rect 187342 532294 187398 532350
rect 186970 532170 187026 532226
rect 187094 532170 187150 532226
rect 187218 532170 187274 532226
rect 187342 532170 187398 532226
rect 186970 532046 187026 532102
rect 187094 532046 187150 532102
rect 187218 532046 187274 532102
rect 187342 532046 187398 532102
rect 186970 531922 187026 531978
rect 187094 531922 187150 531978
rect 187218 531922 187274 531978
rect 187342 531922 187398 531978
rect 186970 514294 187026 514350
rect 187094 514294 187150 514350
rect 187218 514294 187274 514350
rect 187342 514294 187398 514350
rect 186970 514170 187026 514226
rect 187094 514170 187150 514226
rect 187218 514170 187274 514226
rect 187342 514170 187398 514226
rect 186970 514046 187026 514102
rect 187094 514046 187150 514102
rect 187218 514046 187274 514102
rect 187342 514046 187398 514102
rect 186970 513922 187026 513978
rect 187094 513922 187150 513978
rect 187218 513922 187274 513978
rect 187342 513922 187398 513978
rect 186970 496294 187026 496350
rect 187094 496294 187150 496350
rect 187218 496294 187274 496350
rect 187342 496294 187398 496350
rect 186970 496170 187026 496226
rect 187094 496170 187150 496226
rect 187218 496170 187274 496226
rect 187342 496170 187398 496226
rect 186970 496046 187026 496102
rect 187094 496046 187150 496102
rect 187218 496046 187274 496102
rect 187342 496046 187398 496102
rect 186970 495922 187026 495978
rect 187094 495922 187150 495978
rect 187218 495922 187274 495978
rect 187342 495922 187398 495978
rect 186970 478294 187026 478350
rect 187094 478294 187150 478350
rect 187218 478294 187274 478350
rect 187342 478294 187398 478350
rect 186970 478170 187026 478226
rect 187094 478170 187150 478226
rect 187218 478170 187274 478226
rect 187342 478170 187398 478226
rect 186970 478046 187026 478102
rect 187094 478046 187150 478102
rect 187218 478046 187274 478102
rect 187342 478046 187398 478102
rect 186970 477922 187026 477978
rect 187094 477922 187150 477978
rect 187218 477922 187274 477978
rect 187342 477922 187398 477978
rect 186970 460294 187026 460350
rect 187094 460294 187150 460350
rect 187218 460294 187274 460350
rect 187342 460294 187398 460350
rect 186970 460170 187026 460226
rect 187094 460170 187150 460226
rect 187218 460170 187274 460226
rect 187342 460170 187398 460226
rect 186970 460046 187026 460102
rect 187094 460046 187150 460102
rect 187218 460046 187274 460102
rect 187342 460046 187398 460102
rect 186970 459922 187026 459978
rect 187094 459922 187150 459978
rect 187218 459922 187274 459978
rect 187342 459922 187398 459978
rect 186970 442294 187026 442350
rect 187094 442294 187150 442350
rect 187218 442294 187274 442350
rect 187342 442294 187398 442350
rect 186970 442170 187026 442226
rect 187094 442170 187150 442226
rect 187218 442170 187274 442226
rect 187342 442170 187398 442226
rect 186970 442046 187026 442102
rect 187094 442046 187150 442102
rect 187218 442046 187274 442102
rect 187342 442046 187398 442102
rect 186970 441922 187026 441978
rect 187094 441922 187150 441978
rect 187218 441922 187274 441978
rect 187342 441922 187398 441978
rect 186970 424294 187026 424350
rect 187094 424294 187150 424350
rect 187218 424294 187274 424350
rect 187342 424294 187398 424350
rect 186970 424170 187026 424226
rect 187094 424170 187150 424226
rect 187218 424170 187274 424226
rect 187342 424170 187398 424226
rect 186970 424046 187026 424102
rect 187094 424046 187150 424102
rect 187218 424046 187274 424102
rect 187342 424046 187398 424102
rect 186970 423922 187026 423978
rect 187094 423922 187150 423978
rect 187218 423922 187274 423978
rect 187342 423922 187398 423978
rect 186970 406294 187026 406350
rect 187094 406294 187150 406350
rect 187218 406294 187274 406350
rect 187342 406294 187398 406350
rect 186970 406170 187026 406226
rect 187094 406170 187150 406226
rect 187218 406170 187274 406226
rect 187342 406170 187398 406226
rect 186970 406046 187026 406102
rect 187094 406046 187150 406102
rect 187218 406046 187274 406102
rect 187342 406046 187398 406102
rect 186970 405922 187026 405978
rect 187094 405922 187150 405978
rect 187218 405922 187274 405978
rect 187342 405922 187398 405978
rect 186970 388294 187026 388350
rect 187094 388294 187150 388350
rect 187218 388294 187274 388350
rect 187342 388294 187398 388350
rect 186970 388170 187026 388226
rect 187094 388170 187150 388226
rect 187218 388170 187274 388226
rect 187342 388170 187398 388226
rect 186970 388046 187026 388102
rect 187094 388046 187150 388102
rect 187218 388046 187274 388102
rect 187342 388046 187398 388102
rect 186970 387922 187026 387978
rect 187094 387922 187150 387978
rect 187218 387922 187274 387978
rect 187342 387922 187398 387978
rect 186970 370294 187026 370350
rect 187094 370294 187150 370350
rect 187218 370294 187274 370350
rect 187342 370294 187398 370350
rect 186970 370170 187026 370226
rect 187094 370170 187150 370226
rect 187218 370170 187274 370226
rect 187342 370170 187398 370226
rect 186970 370046 187026 370102
rect 187094 370046 187150 370102
rect 187218 370046 187274 370102
rect 187342 370046 187398 370102
rect 186970 369922 187026 369978
rect 187094 369922 187150 369978
rect 187218 369922 187274 369978
rect 187342 369922 187398 369978
rect 186970 352294 187026 352350
rect 187094 352294 187150 352350
rect 187218 352294 187274 352350
rect 187342 352294 187398 352350
rect 186970 352170 187026 352226
rect 187094 352170 187150 352226
rect 187218 352170 187274 352226
rect 187342 352170 187398 352226
rect 186970 352046 187026 352102
rect 187094 352046 187150 352102
rect 187218 352046 187274 352102
rect 187342 352046 187398 352102
rect 186970 351922 187026 351978
rect 187094 351922 187150 351978
rect 187218 351922 187274 351978
rect 187342 351922 187398 351978
rect 186970 334294 187026 334350
rect 187094 334294 187150 334350
rect 187218 334294 187274 334350
rect 187342 334294 187398 334350
rect 186970 334170 187026 334226
rect 187094 334170 187150 334226
rect 187218 334170 187274 334226
rect 187342 334170 187398 334226
rect 186970 334046 187026 334102
rect 187094 334046 187150 334102
rect 187218 334046 187274 334102
rect 187342 334046 187398 334102
rect 186970 333922 187026 333978
rect 187094 333922 187150 333978
rect 187218 333922 187274 333978
rect 187342 333922 187398 333978
rect 186970 316294 187026 316350
rect 187094 316294 187150 316350
rect 187218 316294 187274 316350
rect 187342 316294 187398 316350
rect 186970 316170 187026 316226
rect 187094 316170 187150 316226
rect 187218 316170 187274 316226
rect 187342 316170 187398 316226
rect 186970 316046 187026 316102
rect 187094 316046 187150 316102
rect 187218 316046 187274 316102
rect 187342 316046 187398 316102
rect 186970 315922 187026 315978
rect 187094 315922 187150 315978
rect 187218 315922 187274 315978
rect 187342 315922 187398 315978
rect 186970 298294 187026 298350
rect 187094 298294 187150 298350
rect 187218 298294 187274 298350
rect 187342 298294 187398 298350
rect 186970 298170 187026 298226
rect 187094 298170 187150 298226
rect 187218 298170 187274 298226
rect 187342 298170 187398 298226
rect 186970 298046 187026 298102
rect 187094 298046 187150 298102
rect 187218 298046 187274 298102
rect 187342 298046 187398 298102
rect 186970 297922 187026 297978
rect 187094 297922 187150 297978
rect 187218 297922 187274 297978
rect 187342 297922 187398 297978
rect 186970 280294 187026 280350
rect 187094 280294 187150 280350
rect 187218 280294 187274 280350
rect 187342 280294 187398 280350
rect 186970 280170 187026 280226
rect 187094 280170 187150 280226
rect 187218 280170 187274 280226
rect 187342 280170 187398 280226
rect 186970 280046 187026 280102
rect 187094 280046 187150 280102
rect 187218 280046 187274 280102
rect 187342 280046 187398 280102
rect 186970 279922 187026 279978
rect 187094 279922 187150 279978
rect 187218 279922 187274 279978
rect 187342 279922 187398 279978
rect 186970 262294 187026 262350
rect 187094 262294 187150 262350
rect 187218 262294 187274 262350
rect 187342 262294 187398 262350
rect 186970 262170 187026 262226
rect 187094 262170 187150 262226
rect 187218 262170 187274 262226
rect 187342 262170 187398 262226
rect 186970 262046 187026 262102
rect 187094 262046 187150 262102
rect 187218 262046 187274 262102
rect 187342 262046 187398 262102
rect 186970 261922 187026 261978
rect 187094 261922 187150 261978
rect 187218 261922 187274 261978
rect 187342 261922 187398 261978
rect 186970 244294 187026 244350
rect 187094 244294 187150 244350
rect 187218 244294 187274 244350
rect 187342 244294 187398 244350
rect 186970 244170 187026 244226
rect 187094 244170 187150 244226
rect 187218 244170 187274 244226
rect 187342 244170 187398 244226
rect 186970 244046 187026 244102
rect 187094 244046 187150 244102
rect 187218 244046 187274 244102
rect 187342 244046 187398 244102
rect 186970 243922 187026 243978
rect 187094 243922 187150 243978
rect 187218 243922 187274 243978
rect 187342 243922 187398 243978
rect 201250 597156 201306 597212
rect 201374 597156 201430 597212
rect 201498 597156 201554 597212
rect 201622 597156 201678 597212
rect 201250 597032 201306 597088
rect 201374 597032 201430 597088
rect 201498 597032 201554 597088
rect 201622 597032 201678 597088
rect 201250 596908 201306 596964
rect 201374 596908 201430 596964
rect 201498 596908 201554 596964
rect 201622 596908 201678 596964
rect 201250 596784 201306 596840
rect 201374 596784 201430 596840
rect 201498 596784 201554 596840
rect 201622 596784 201678 596840
rect 201250 580294 201306 580350
rect 201374 580294 201430 580350
rect 201498 580294 201554 580350
rect 201622 580294 201678 580350
rect 201250 580170 201306 580226
rect 201374 580170 201430 580226
rect 201498 580170 201554 580226
rect 201622 580170 201678 580226
rect 201250 580046 201306 580102
rect 201374 580046 201430 580102
rect 201498 580046 201554 580102
rect 201622 580046 201678 580102
rect 201250 579922 201306 579978
rect 201374 579922 201430 579978
rect 201498 579922 201554 579978
rect 201622 579922 201678 579978
rect 201250 562294 201306 562350
rect 201374 562294 201430 562350
rect 201498 562294 201554 562350
rect 201622 562294 201678 562350
rect 201250 562170 201306 562226
rect 201374 562170 201430 562226
rect 201498 562170 201554 562226
rect 201622 562170 201678 562226
rect 201250 562046 201306 562102
rect 201374 562046 201430 562102
rect 201498 562046 201554 562102
rect 201622 562046 201678 562102
rect 201250 561922 201306 561978
rect 201374 561922 201430 561978
rect 201498 561922 201554 561978
rect 201622 561922 201678 561978
rect 201250 544294 201306 544350
rect 201374 544294 201430 544350
rect 201498 544294 201554 544350
rect 201622 544294 201678 544350
rect 201250 544170 201306 544226
rect 201374 544170 201430 544226
rect 201498 544170 201554 544226
rect 201622 544170 201678 544226
rect 201250 544046 201306 544102
rect 201374 544046 201430 544102
rect 201498 544046 201554 544102
rect 201622 544046 201678 544102
rect 201250 543922 201306 543978
rect 201374 543922 201430 543978
rect 201498 543922 201554 543978
rect 201622 543922 201678 543978
rect 201250 526294 201306 526350
rect 201374 526294 201430 526350
rect 201498 526294 201554 526350
rect 201622 526294 201678 526350
rect 201250 526170 201306 526226
rect 201374 526170 201430 526226
rect 201498 526170 201554 526226
rect 201622 526170 201678 526226
rect 201250 526046 201306 526102
rect 201374 526046 201430 526102
rect 201498 526046 201554 526102
rect 201622 526046 201678 526102
rect 201250 525922 201306 525978
rect 201374 525922 201430 525978
rect 201498 525922 201554 525978
rect 201622 525922 201678 525978
rect 201250 508294 201306 508350
rect 201374 508294 201430 508350
rect 201498 508294 201554 508350
rect 201622 508294 201678 508350
rect 201250 508170 201306 508226
rect 201374 508170 201430 508226
rect 201498 508170 201554 508226
rect 201622 508170 201678 508226
rect 201250 508046 201306 508102
rect 201374 508046 201430 508102
rect 201498 508046 201554 508102
rect 201622 508046 201678 508102
rect 201250 507922 201306 507978
rect 201374 507922 201430 507978
rect 201498 507922 201554 507978
rect 201622 507922 201678 507978
rect 201250 490294 201306 490350
rect 201374 490294 201430 490350
rect 201498 490294 201554 490350
rect 201622 490294 201678 490350
rect 201250 490170 201306 490226
rect 201374 490170 201430 490226
rect 201498 490170 201554 490226
rect 201622 490170 201678 490226
rect 201250 490046 201306 490102
rect 201374 490046 201430 490102
rect 201498 490046 201554 490102
rect 201622 490046 201678 490102
rect 201250 489922 201306 489978
rect 201374 489922 201430 489978
rect 201498 489922 201554 489978
rect 201622 489922 201678 489978
rect 201250 472294 201306 472350
rect 201374 472294 201430 472350
rect 201498 472294 201554 472350
rect 201622 472294 201678 472350
rect 201250 472170 201306 472226
rect 201374 472170 201430 472226
rect 201498 472170 201554 472226
rect 201622 472170 201678 472226
rect 201250 472046 201306 472102
rect 201374 472046 201430 472102
rect 201498 472046 201554 472102
rect 201622 472046 201678 472102
rect 201250 471922 201306 471978
rect 201374 471922 201430 471978
rect 201498 471922 201554 471978
rect 201622 471922 201678 471978
rect 201250 454294 201306 454350
rect 201374 454294 201430 454350
rect 201498 454294 201554 454350
rect 201622 454294 201678 454350
rect 201250 454170 201306 454226
rect 201374 454170 201430 454226
rect 201498 454170 201554 454226
rect 201622 454170 201678 454226
rect 201250 454046 201306 454102
rect 201374 454046 201430 454102
rect 201498 454046 201554 454102
rect 201622 454046 201678 454102
rect 201250 453922 201306 453978
rect 201374 453922 201430 453978
rect 201498 453922 201554 453978
rect 201622 453922 201678 453978
rect 201250 436294 201306 436350
rect 201374 436294 201430 436350
rect 201498 436294 201554 436350
rect 201622 436294 201678 436350
rect 201250 436170 201306 436226
rect 201374 436170 201430 436226
rect 201498 436170 201554 436226
rect 201622 436170 201678 436226
rect 201250 436046 201306 436102
rect 201374 436046 201430 436102
rect 201498 436046 201554 436102
rect 201622 436046 201678 436102
rect 201250 435922 201306 435978
rect 201374 435922 201430 435978
rect 201498 435922 201554 435978
rect 201622 435922 201678 435978
rect 201250 418294 201306 418350
rect 201374 418294 201430 418350
rect 201498 418294 201554 418350
rect 201622 418294 201678 418350
rect 201250 418170 201306 418226
rect 201374 418170 201430 418226
rect 201498 418170 201554 418226
rect 201622 418170 201678 418226
rect 201250 418046 201306 418102
rect 201374 418046 201430 418102
rect 201498 418046 201554 418102
rect 201622 418046 201678 418102
rect 201250 417922 201306 417978
rect 201374 417922 201430 417978
rect 201498 417922 201554 417978
rect 201622 417922 201678 417978
rect 201250 400294 201306 400350
rect 201374 400294 201430 400350
rect 201498 400294 201554 400350
rect 201622 400294 201678 400350
rect 201250 400170 201306 400226
rect 201374 400170 201430 400226
rect 201498 400170 201554 400226
rect 201622 400170 201678 400226
rect 201250 400046 201306 400102
rect 201374 400046 201430 400102
rect 201498 400046 201554 400102
rect 201622 400046 201678 400102
rect 201250 399922 201306 399978
rect 201374 399922 201430 399978
rect 201498 399922 201554 399978
rect 201622 399922 201678 399978
rect 201250 382294 201306 382350
rect 201374 382294 201430 382350
rect 201498 382294 201554 382350
rect 201622 382294 201678 382350
rect 201250 382170 201306 382226
rect 201374 382170 201430 382226
rect 201498 382170 201554 382226
rect 201622 382170 201678 382226
rect 201250 382046 201306 382102
rect 201374 382046 201430 382102
rect 201498 382046 201554 382102
rect 201622 382046 201678 382102
rect 201250 381922 201306 381978
rect 201374 381922 201430 381978
rect 201498 381922 201554 381978
rect 201622 381922 201678 381978
rect 201250 364294 201306 364350
rect 201374 364294 201430 364350
rect 201498 364294 201554 364350
rect 201622 364294 201678 364350
rect 201250 364170 201306 364226
rect 201374 364170 201430 364226
rect 201498 364170 201554 364226
rect 201622 364170 201678 364226
rect 201250 364046 201306 364102
rect 201374 364046 201430 364102
rect 201498 364046 201554 364102
rect 201622 364046 201678 364102
rect 201250 363922 201306 363978
rect 201374 363922 201430 363978
rect 201498 363922 201554 363978
rect 201622 363922 201678 363978
rect 201250 346294 201306 346350
rect 201374 346294 201430 346350
rect 201498 346294 201554 346350
rect 201622 346294 201678 346350
rect 201250 346170 201306 346226
rect 201374 346170 201430 346226
rect 201498 346170 201554 346226
rect 201622 346170 201678 346226
rect 201250 346046 201306 346102
rect 201374 346046 201430 346102
rect 201498 346046 201554 346102
rect 201622 346046 201678 346102
rect 201250 345922 201306 345978
rect 201374 345922 201430 345978
rect 201498 345922 201554 345978
rect 201622 345922 201678 345978
rect 201250 328294 201306 328350
rect 201374 328294 201430 328350
rect 201498 328294 201554 328350
rect 201622 328294 201678 328350
rect 201250 328170 201306 328226
rect 201374 328170 201430 328226
rect 201498 328170 201554 328226
rect 201622 328170 201678 328226
rect 201250 328046 201306 328102
rect 201374 328046 201430 328102
rect 201498 328046 201554 328102
rect 201622 328046 201678 328102
rect 201250 327922 201306 327978
rect 201374 327922 201430 327978
rect 201498 327922 201554 327978
rect 201622 327922 201678 327978
rect 201250 310294 201306 310350
rect 201374 310294 201430 310350
rect 201498 310294 201554 310350
rect 201622 310294 201678 310350
rect 201250 310170 201306 310226
rect 201374 310170 201430 310226
rect 201498 310170 201554 310226
rect 201622 310170 201678 310226
rect 201250 310046 201306 310102
rect 201374 310046 201430 310102
rect 201498 310046 201554 310102
rect 201622 310046 201678 310102
rect 201250 309922 201306 309978
rect 201374 309922 201430 309978
rect 201498 309922 201554 309978
rect 201622 309922 201678 309978
rect 201250 292294 201306 292350
rect 201374 292294 201430 292350
rect 201498 292294 201554 292350
rect 201622 292294 201678 292350
rect 201250 292170 201306 292226
rect 201374 292170 201430 292226
rect 201498 292170 201554 292226
rect 201622 292170 201678 292226
rect 201250 292046 201306 292102
rect 201374 292046 201430 292102
rect 201498 292046 201554 292102
rect 201622 292046 201678 292102
rect 201250 291922 201306 291978
rect 201374 291922 201430 291978
rect 201498 291922 201554 291978
rect 201622 291922 201678 291978
rect 201250 274294 201306 274350
rect 201374 274294 201430 274350
rect 201498 274294 201554 274350
rect 201622 274294 201678 274350
rect 201250 274170 201306 274226
rect 201374 274170 201430 274226
rect 201498 274170 201554 274226
rect 201622 274170 201678 274226
rect 201250 274046 201306 274102
rect 201374 274046 201430 274102
rect 201498 274046 201554 274102
rect 201622 274046 201678 274102
rect 201250 273922 201306 273978
rect 201374 273922 201430 273978
rect 201498 273922 201554 273978
rect 201622 273922 201678 273978
rect 201250 256294 201306 256350
rect 201374 256294 201430 256350
rect 201498 256294 201554 256350
rect 201622 256294 201678 256350
rect 201250 256170 201306 256226
rect 201374 256170 201430 256226
rect 201498 256170 201554 256226
rect 201622 256170 201678 256226
rect 201250 256046 201306 256102
rect 201374 256046 201430 256102
rect 201498 256046 201554 256102
rect 201622 256046 201678 256102
rect 201250 255922 201306 255978
rect 201374 255922 201430 255978
rect 201498 255922 201554 255978
rect 201622 255922 201678 255978
rect 219250 597156 219306 597212
rect 219374 597156 219430 597212
rect 219498 597156 219554 597212
rect 219622 597156 219678 597212
rect 219250 597032 219306 597088
rect 219374 597032 219430 597088
rect 219498 597032 219554 597088
rect 219622 597032 219678 597088
rect 219250 596908 219306 596964
rect 219374 596908 219430 596964
rect 219498 596908 219554 596964
rect 219622 596908 219678 596964
rect 219250 596784 219306 596840
rect 219374 596784 219430 596840
rect 219498 596784 219554 596840
rect 219622 596784 219678 596840
rect 219250 580294 219306 580350
rect 219374 580294 219430 580350
rect 219498 580294 219554 580350
rect 219622 580294 219678 580350
rect 219250 580170 219306 580226
rect 219374 580170 219430 580226
rect 219498 580170 219554 580226
rect 219622 580170 219678 580226
rect 219250 580046 219306 580102
rect 219374 580046 219430 580102
rect 219498 580046 219554 580102
rect 219622 580046 219678 580102
rect 219250 579922 219306 579978
rect 219374 579922 219430 579978
rect 219498 579922 219554 579978
rect 219622 579922 219678 579978
rect 219250 562294 219306 562350
rect 219374 562294 219430 562350
rect 219498 562294 219554 562350
rect 219622 562294 219678 562350
rect 219250 562170 219306 562226
rect 219374 562170 219430 562226
rect 219498 562170 219554 562226
rect 219622 562170 219678 562226
rect 219250 562046 219306 562102
rect 219374 562046 219430 562102
rect 219498 562046 219554 562102
rect 219622 562046 219678 562102
rect 219250 561922 219306 561978
rect 219374 561922 219430 561978
rect 219498 561922 219554 561978
rect 219622 561922 219678 561978
rect 219250 544294 219306 544350
rect 219374 544294 219430 544350
rect 219498 544294 219554 544350
rect 219622 544294 219678 544350
rect 219250 544170 219306 544226
rect 219374 544170 219430 544226
rect 219498 544170 219554 544226
rect 219622 544170 219678 544226
rect 219250 544046 219306 544102
rect 219374 544046 219430 544102
rect 219498 544046 219554 544102
rect 219622 544046 219678 544102
rect 219250 543922 219306 543978
rect 219374 543922 219430 543978
rect 219498 543922 219554 543978
rect 219622 543922 219678 543978
rect 219250 526294 219306 526350
rect 219374 526294 219430 526350
rect 219498 526294 219554 526350
rect 219622 526294 219678 526350
rect 219250 526170 219306 526226
rect 219374 526170 219430 526226
rect 219498 526170 219554 526226
rect 219622 526170 219678 526226
rect 219250 526046 219306 526102
rect 219374 526046 219430 526102
rect 219498 526046 219554 526102
rect 219622 526046 219678 526102
rect 219250 525922 219306 525978
rect 219374 525922 219430 525978
rect 219498 525922 219554 525978
rect 219622 525922 219678 525978
rect 219250 508294 219306 508350
rect 219374 508294 219430 508350
rect 219498 508294 219554 508350
rect 219622 508294 219678 508350
rect 219250 508170 219306 508226
rect 219374 508170 219430 508226
rect 219498 508170 219554 508226
rect 219622 508170 219678 508226
rect 219250 508046 219306 508102
rect 219374 508046 219430 508102
rect 219498 508046 219554 508102
rect 219622 508046 219678 508102
rect 219250 507922 219306 507978
rect 219374 507922 219430 507978
rect 219498 507922 219554 507978
rect 219622 507922 219678 507978
rect 219250 490294 219306 490350
rect 219374 490294 219430 490350
rect 219498 490294 219554 490350
rect 219622 490294 219678 490350
rect 219250 490170 219306 490226
rect 219374 490170 219430 490226
rect 219498 490170 219554 490226
rect 219622 490170 219678 490226
rect 219250 490046 219306 490102
rect 219374 490046 219430 490102
rect 219498 490046 219554 490102
rect 219622 490046 219678 490102
rect 219250 489922 219306 489978
rect 219374 489922 219430 489978
rect 219498 489922 219554 489978
rect 219622 489922 219678 489978
rect 219250 472294 219306 472350
rect 219374 472294 219430 472350
rect 219498 472294 219554 472350
rect 219622 472294 219678 472350
rect 219250 472170 219306 472226
rect 219374 472170 219430 472226
rect 219498 472170 219554 472226
rect 219622 472170 219678 472226
rect 219250 472046 219306 472102
rect 219374 472046 219430 472102
rect 219498 472046 219554 472102
rect 219622 472046 219678 472102
rect 219250 471922 219306 471978
rect 219374 471922 219430 471978
rect 219498 471922 219554 471978
rect 219622 471922 219678 471978
rect 219250 454294 219306 454350
rect 219374 454294 219430 454350
rect 219498 454294 219554 454350
rect 219622 454294 219678 454350
rect 219250 454170 219306 454226
rect 219374 454170 219430 454226
rect 219498 454170 219554 454226
rect 219622 454170 219678 454226
rect 219250 454046 219306 454102
rect 219374 454046 219430 454102
rect 219498 454046 219554 454102
rect 219622 454046 219678 454102
rect 219250 453922 219306 453978
rect 219374 453922 219430 453978
rect 219498 453922 219554 453978
rect 219622 453922 219678 453978
rect 219250 436294 219306 436350
rect 219374 436294 219430 436350
rect 219498 436294 219554 436350
rect 219622 436294 219678 436350
rect 219250 436170 219306 436226
rect 219374 436170 219430 436226
rect 219498 436170 219554 436226
rect 219622 436170 219678 436226
rect 219250 436046 219306 436102
rect 219374 436046 219430 436102
rect 219498 436046 219554 436102
rect 219622 436046 219678 436102
rect 219250 435922 219306 435978
rect 219374 435922 219430 435978
rect 219498 435922 219554 435978
rect 219622 435922 219678 435978
rect 219250 418294 219306 418350
rect 219374 418294 219430 418350
rect 219498 418294 219554 418350
rect 219622 418294 219678 418350
rect 219250 418170 219306 418226
rect 219374 418170 219430 418226
rect 219498 418170 219554 418226
rect 219622 418170 219678 418226
rect 219250 418046 219306 418102
rect 219374 418046 219430 418102
rect 219498 418046 219554 418102
rect 219622 418046 219678 418102
rect 219250 417922 219306 417978
rect 219374 417922 219430 417978
rect 219498 417922 219554 417978
rect 219622 417922 219678 417978
rect 219250 400294 219306 400350
rect 219374 400294 219430 400350
rect 219498 400294 219554 400350
rect 219622 400294 219678 400350
rect 219250 400170 219306 400226
rect 219374 400170 219430 400226
rect 219498 400170 219554 400226
rect 219622 400170 219678 400226
rect 219250 400046 219306 400102
rect 219374 400046 219430 400102
rect 219498 400046 219554 400102
rect 219622 400046 219678 400102
rect 219250 399922 219306 399978
rect 219374 399922 219430 399978
rect 219498 399922 219554 399978
rect 219622 399922 219678 399978
rect 219250 382294 219306 382350
rect 219374 382294 219430 382350
rect 219498 382294 219554 382350
rect 219622 382294 219678 382350
rect 219250 382170 219306 382226
rect 219374 382170 219430 382226
rect 219498 382170 219554 382226
rect 219622 382170 219678 382226
rect 219250 382046 219306 382102
rect 219374 382046 219430 382102
rect 219498 382046 219554 382102
rect 219622 382046 219678 382102
rect 219250 381922 219306 381978
rect 219374 381922 219430 381978
rect 219498 381922 219554 381978
rect 219622 381922 219678 381978
rect 219250 364294 219306 364350
rect 219374 364294 219430 364350
rect 219498 364294 219554 364350
rect 219622 364294 219678 364350
rect 219250 364170 219306 364226
rect 219374 364170 219430 364226
rect 219498 364170 219554 364226
rect 219622 364170 219678 364226
rect 219250 364046 219306 364102
rect 219374 364046 219430 364102
rect 219498 364046 219554 364102
rect 219622 364046 219678 364102
rect 219250 363922 219306 363978
rect 219374 363922 219430 363978
rect 219498 363922 219554 363978
rect 219622 363922 219678 363978
rect 219250 346294 219306 346350
rect 219374 346294 219430 346350
rect 219498 346294 219554 346350
rect 219622 346294 219678 346350
rect 219250 346170 219306 346226
rect 219374 346170 219430 346226
rect 219498 346170 219554 346226
rect 219622 346170 219678 346226
rect 219250 346046 219306 346102
rect 219374 346046 219430 346102
rect 219498 346046 219554 346102
rect 219622 346046 219678 346102
rect 219250 345922 219306 345978
rect 219374 345922 219430 345978
rect 219498 345922 219554 345978
rect 219622 345922 219678 345978
rect 219250 328294 219306 328350
rect 219374 328294 219430 328350
rect 219498 328294 219554 328350
rect 219622 328294 219678 328350
rect 219250 328170 219306 328226
rect 219374 328170 219430 328226
rect 219498 328170 219554 328226
rect 219622 328170 219678 328226
rect 219250 328046 219306 328102
rect 219374 328046 219430 328102
rect 219498 328046 219554 328102
rect 219622 328046 219678 328102
rect 219250 327922 219306 327978
rect 219374 327922 219430 327978
rect 219498 327922 219554 327978
rect 219622 327922 219678 327978
rect 219250 310294 219306 310350
rect 219374 310294 219430 310350
rect 219498 310294 219554 310350
rect 219622 310294 219678 310350
rect 219250 310170 219306 310226
rect 219374 310170 219430 310226
rect 219498 310170 219554 310226
rect 219622 310170 219678 310226
rect 219250 310046 219306 310102
rect 219374 310046 219430 310102
rect 219498 310046 219554 310102
rect 219622 310046 219678 310102
rect 219250 309922 219306 309978
rect 219374 309922 219430 309978
rect 219498 309922 219554 309978
rect 219622 309922 219678 309978
rect 219250 292294 219306 292350
rect 219374 292294 219430 292350
rect 219498 292294 219554 292350
rect 219622 292294 219678 292350
rect 219250 292170 219306 292226
rect 219374 292170 219430 292226
rect 219498 292170 219554 292226
rect 219622 292170 219678 292226
rect 219250 292046 219306 292102
rect 219374 292046 219430 292102
rect 219498 292046 219554 292102
rect 219622 292046 219678 292102
rect 219250 291922 219306 291978
rect 219374 291922 219430 291978
rect 219498 291922 219554 291978
rect 219622 291922 219678 291978
rect 219250 274294 219306 274350
rect 219374 274294 219430 274350
rect 219498 274294 219554 274350
rect 219622 274294 219678 274350
rect 219250 274170 219306 274226
rect 219374 274170 219430 274226
rect 219498 274170 219554 274226
rect 219622 274170 219678 274226
rect 219250 274046 219306 274102
rect 219374 274046 219430 274102
rect 219498 274046 219554 274102
rect 219622 274046 219678 274102
rect 219250 273922 219306 273978
rect 219374 273922 219430 273978
rect 219498 273922 219554 273978
rect 219622 273922 219678 273978
rect 219250 256294 219306 256350
rect 219374 256294 219430 256350
rect 219498 256294 219554 256350
rect 219622 256294 219678 256350
rect 219250 256170 219306 256226
rect 219374 256170 219430 256226
rect 219498 256170 219554 256226
rect 219622 256170 219678 256226
rect 219250 256046 219306 256102
rect 219374 256046 219430 256102
rect 219498 256046 219554 256102
rect 219622 256046 219678 256102
rect 219250 255922 219306 255978
rect 219374 255922 219430 255978
rect 219498 255922 219554 255978
rect 219622 255922 219678 255978
rect 201250 238294 201306 238350
rect 201374 238294 201430 238350
rect 201498 238294 201554 238350
rect 201622 238294 201678 238350
rect 201250 238170 201306 238226
rect 201374 238170 201430 238226
rect 201498 238170 201554 238226
rect 201622 238170 201678 238226
rect 201250 238046 201306 238102
rect 201374 238046 201430 238102
rect 201498 238046 201554 238102
rect 201622 238046 201678 238102
rect 201250 237922 201306 237978
rect 201374 237922 201430 237978
rect 201498 237922 201554 237978
rect 201622 237922 201678 237978
rect 183250 220294 183306 220350
rect 183374 220294 183430 220350
rect 183498 220294 183554 220350
rect 183622 220294 183678 220350
rect 183250 220170 183306 220226
rect 183374 220170 183430 220226
rect 183498 220170 183554 220226
rect 183622 220170 183678 220226
rect 183250 220046 183306 220102
rect 183374 220046 183430 220102
rect 183498 220046 183554 220102
rect 183622 220046 183678 220102
rect 183250 219922 183306 219978
rect 183374 219922 183430 219978
rect 183498 219922 183554 219978
rect 183622 219922 183678 219978
rect 187398 220294 187454 220350
rect 187522 220294 187578 220350
rect 187398 220170 187454 220226
rect 187522 220170 187578 220226
rect 187398 220046 187454 220102
rect 187522 220046 187578 220102
rect 187398 219922 187454 219978
rect 187522 219922 187578 219978
rect 202758 226294 202814 226350
rect 202882 226294 202938 226350
rect 202758 226170 202814 226226
rect 202882 226170 202938 226226
rect 202758 226046 202814 226102
rect 202882 226046 202938 226102
rect 202758 225922 202814 225978
rect 202882 225922 202938 225978
rect 204970 226294 205026 226350
rect 205094 226294 205150 226350
rect 205218 226294 205274 226350
rect 205342 226294 205398 226350
rect 204970 226170 205026 226226
rect 205094 226170 205150 226226
rect 205218 226170 205274 226226
rect 205342 226170 205398 226226
rect 204970 226046 205026 226102
rect 205094 226046 205150 226102
rect 205218 226046 205274 226102
rect 205342 226046 205398 226102
rect 204970 225922 205026 225978
rect 205094 225922 205150 225978
rect 205218 225922 205274 225978
rect 205342 225922 205398 225978
rect 201250 220294 201306 220350
rect 201374 220294 201430 220350
rect 201498 220294 201554 220350
rect 201622 220294 201678 220350
rect 201250 220170 201306 220226
rect 201374 220170 201430 220226
rect 201498 220170 201554 220226
rect 201622 220170 201678 220226
rect 201250 220046 201306 220102
rect 201374 220046 201430 220102
rect 201498 220046 201554 220102
rect 201622 220046 201678 220102
rect 201250 219922 201306 219978
rect 201374 219922 201430 219978
rect 201498 219922 201554 219978
rect 201622 219922 201678 219978
rect 219250 238294 219306 238350
rect 219374 238294 219430 238350
rect 219498 238294 219554 238350
rect 219622 238294 219678 238350
rect 219250 238170 219306 238226
rect 219374 238170 219430 238226
rect 219498 238170 219554 238226
rect 219622 238170 219678 238226
rect 219250 238046 219306 238102
rect 219374 238046 219430 238102
rect 219498 238046 219554 238102
rect 219622 238046 219678 238102
rect 219250 237922 219306 237978
rect 219374 237922 219430 237978
rect 219498 237922 219554 237978
rect 219622 237922 219678 237978
rect 218118 220294 218174 220350
rect 218242 220294 218298 220350
rect 218118 220170 218174 220226
rect 218242 220170 218298 220226
rect 218118 220046 218174 220102
rect 218242 220046 218298 220102
rect 218118 219922 218174 219978
rect 218242 219922 218298 219978
rect 219250 220294 219306 220350
rect 219374 220294 219430 220350
rect 219498 220294 219554 220350
rect 219622 220294 219678 220350
rect 219250 220170 219306 220226
rect 219374 220170 219430 220226
rect 219498 220170 219554 220226
rect 219622 220170 219678 220226
rect 219250 220046 219306 220102
rect 219374 220046 219430 220102
rect 219498 220046 219554 220102
rect 219622 220046 219678 220102
rect 219250 219922 219306 219978
rect 219374 219922 219430 219978
rect 219498 219922 219554 219978
rect 219622 219922 219678 219978
rect 222970 598116 223026 598172
rect 223094 598116 223150 598172
rect 223218 598116 223274 598172
rect 223342 598116 223398 598172
rect 222970 597992 223026 598048
rect 223094 597992 223150 598048
rect 223218 597992 223274 598048
rect 223342 597992 223398 598048
rect 222970 597868 223026 597924
rect 223094 597868 223150 597924
rect 223218 597868 223274 597924
rect 223342 597868 223398 597924
rect 222970 597744 223026 597800
rect 223094 597744 223150 597800
rect 223218 597744 223274 597800
rect 223342 597744 223398 597800
rect 222970 586294 223026 586350
rect 223094 586294 223150 586350
rect 223218 586294 223274 586350
rect 223342 586294 223398 586350
rect 222970 586170 223026 586226
rect 223094 586170 223150 586226
rect 223218 586170 223274 586226
rect 223342 586170 223398 586226
rect 222970 586046 223026 586102
rect 223094 586046 223150 586102
rect 223218 586046 223274 586102
rect 223342 586046 223398 586102
rect 222970 585922 223026 585978
rect 223094 585922 223150 585978
rect 223218 585922 223274 585978
rect 223342 585922 223398 585978
rect 222970 568294 223026 568350
rect 223094 568294 223150 568350
rect 223218 568294 223274 568350
rect 223342 568294 223398 568350
rect 222970 568170 223026 568226
rect 223094 568170 223150 568226
rect 223218 568170 223274 568226
rect 223342 568170 223398 568226
rect 222970 568046 223026 568102
rect 223094 568046 223150 568102
rect 223218 568046 223274 568102
rect 223342 568046 223398 568102
rect 222970 567922 223026 567978
rect 223094 567922 223150 567978
rect 223218 567922 223274 567978
rect 223342 567922 223398 567978
rect 222970 550294 223026 550350
rect 223094 550294 223150 550350
rect 223218 550294 223274 550350
rect 223342 550294 223398 550350
rect 222970 550170 223026 550226
rect 223094 550170 223150 550226
rect 223218 550170 223274 550226
rect 223342 550170 223398 550226
rect 222970 550046 223026 550102
rect 223094 550046 223150 550102
rect 223218 550046 223274 550102
rect 223342 550046 223398 550102
rect 222970 549922 223026 549978
rect 223094 549922 223150 549978
rect 223218 549922 223274 549978
rect 223342 549922 223398 549978
rect 222970 532294 223026 532350
rect 223094 532294 223150 532350
rect 223218 532294 223274 532350
rect 223342 532294 223398 532350
rect 222970 532170 223026 532226
rect 223094 532170 223150 532226
rect 223218 532170 223274 532226
rect 223342 532170 223398 532226
rect 222970 532046 223026 532102
rect 223094 532046 223150 532102
rect 223218 532046 223274 532102
rect 223342 532046 223398 532102
rect 222970 531922 223026 531978
rect 223094 531922 223150 531978
rect 223218 531922 223274 531978
rect 223342 531922 223398 531978
rect 222970 514294 223026 514350
rect 223094 514294 223150 514350
rect 223218 514294 223274 514350
rect 223342 514294 223398 514350
rect 222970 514170 223026 514226
rect 223094 514170 223150 514226
rect 223218 514170 223274 514226
rect 223342 514170 223398 514226
rect 222970 514046 223026 514102
rect 223094 514046 223150 514102
rect 223218 514046 223274 514102
rect 223342 514046 223398 514102
rect 222970 513922 223026 513978
rect 223094 513922 223150 513978
rect 223218 513922 223274 513978
rect 223342 513922 223398 513978
rect 222970 496294 223026 496350
rect 223094 496294 223150 496350
rect 223218 496294 223274 496350
rect 223342 496294 223398 496350
rect 222970 496170 223026 496226
rect 223094 496170 223150 496226
rect 223218 496170 223274 496226
rect 223342 496170 223398 496226
rect 222970 496046 223026 496102
rect 223094 496046 223150 496102
rect 223218 496046 223274 496102
rect 223342 496046 223398 496102
rect 222970 495922 223026 495978
rect 223094 495922 223150 495978
rect 223218 495922 223274 495978
rect 223342 495922 223398 495978
rect 222970 478294 223026 478350
rect 223094 478294 223150 478350
rect 223218 478294 223274 478350
rect 223342 478294 223398 478350
rect 222970 478170 223026 478226
rect 223094 478170 223150 478226
rect 223218 478170 223274 478226
rect 223342 478170 223398 478226
rect 222970 478046 223026 478102
rect 223094 478046 223150 478102
rect 223218 478046 223274 478102
rect 223342 478046 223398 478102
rect 222970 477922 223026 477978
rect 223094 477922 223150 477978
rect 223218 477922 223274 477978
rect 223342 477922 223398 477978
rect 222970 460294 223026 460350
rect 223094 460294 223150 460350
rect 223218 460294 223274 460350
rect 223342 460294 223398 460350
rect 222970 460170 223026 460226
rect 223094 460170 223150 460226
rect 223218 460170 223274 460226
rect 223342 460170 223398 460226
rect 222970 460046 223026 460102
rect 223094 460046 223150 460102
rect 223218 460046 223274 460102
rect 223342 460046 223398 460102
rect 222970 459922 223026 459978
rect 223094 459922 223150 459978
rect 223218 459922 223274 459978
rect 223342 459922 223398 459978
rect 222970 442294 223026 442350
rect 223094 442294 223150 442350
rect 223218 442294 223274 442350
rect 223342 442294 223398 442350
rect 222970 442170 223026 442226
rect 223094 442170 223150 442226
rect 223218 442170 223274 442226
rect 223342 442170 223398 442226
rect 222970 442046 223026 442102
rect 223094 442046 223150 442102
rect 223218 442046 223274 442102
rect 223342 442046 223398 442102
rect 222970 441922 223026 441978
rect 223094 441922 223150 441978
rect 223218 441922 223274 441978
rect 223342 441922 223398 441978
rect 222970 424294 223026 424350
rect 223094 424294 223150 424350
rect 223218 424294 223274 424350
rect 223342 424294 223398 424350
rect 222970 424170 223026 424226
rect 223094 424170 223150 424226
rect 223218 424170 223274 424226
rect 223342 424170 223398 424226
rect 222970 424046 223026 424102
rect 223094 424046 223150 424102
rect 223218 424046 223274 424102
rect 223342 424046 223398 424102
rect 222970 423922 223026 423978
rect 223094 423922 223150 423978
rect 223218 423922 223274 423978
rect 223342 423922 223398 423978
rect 222970 406294 223026 406350
rect 223094 406294 223150 406350
rect 223218 406294 223274 406350
rect 223342 406294 223398 406350
rect 222970 406170 223026 406226
rect 223094 406170 223150 406226
rect 223218 406170 223274 406226
rect 223342 406170 223398 406226
rect 222970 406046 223026 406102
rect 223094 406046 223150 406102
rect 223218 406046 223274 406102
rect 223342 406046 223398 406102
rect 222970 405922 223026 405978
rect 223094 405922 223150 405978
rect 223218 405922 223274 405978
rect 223342 405922 223398 405978
rect 222970 388294 223026 388350
rect 223094 388294 223150 388350
rect 223218 388294 223274 388350
rect 223342 388294 223398 388350
rect 222970 388170 223026 388226
rect 223094 388170 223150 388226
rect 223218 388170 223274 388226
rect 223342 388170 223398 388226
rect 222970 388046 223026 388102
rect 223094 388046 223150 388102
rect 223218 388046 223274 388102
rect 223342 388046 223398 388102
rect 222970 387922 223026 387978
rect 223094 387922 223150 387978
rect 223218 387922 223274 387978
rect 223342 387922 223398 387978
rect 222970 370294 223026 370350
rect 223094 370294 223150 370350
rect 223218 370294 223274 370350
rect 223342 370294 223398 370350
rect 222970 370170 223026 370226
rect 223094 370170 223150 370226
rect 223218 370170 223274 370226
rect 223342 370170 223398 370226
rect 222970 370046 223026 370102
rect 223094 370046 223150 370102
rect 223218 370046 223274 370102
rect 223342 370046 223398 370102
rect 222970 369922 223026 369978
rect 223094 369922 223150 369978
rect 223218 369922 223274 369978
rect 223342 369922 223398 369978
rect 222970 352294 223026 352350
rect 223094 352294 223150 352350
rect 223218 352294 223274 352350
rect 223342 352294 223398 352350
rect 222970 352170 223026 352226
rect 223094 352170 223150 352226
rect 223218 352170 223274 352226
rect 223342 352170 223398 352226
rect 222970 352046 223026 352102
rect 223094 352046 223150 352102
rect 223218 352046 223274 352102
rect 223342 352046 223398 352102
rect 222970 351922 223026 351978
rect 223094 351922 223150 351978
rect 223218 351922 223274 351978
rect 223342 351922 223398 351978
rect 222970 334294 223026 334350
rect 223094 334294 223150 334350
rect 223218 334294 223274 334350
rect 223342 334294 223398 334350
rect 222970 334170 223026 334226
rect 223094 334170 223150 334226
rect 223218 334170 223274 334226
rect 223342 334170 223398 334226
rect 222970 334046 223026 334102
rect 223094 334046 223150 334102
rect 223218 334046 223274 334102
rect 223342 334046 223398 334102
rect 222970 333922 223026 333978
rect 223094 333922 223150 333978
rect 223218 333922 223274 333978
rect 223342 333922 223398 333978
rect 222970 316294 223026 316350
rect 223094 316294 223150 316350
rect 223218 316294 223274 316350
rect 223342 316294 223398 316350
rect 222970 316170 223026 316226
rect 223094 316170 223150 316226
rect 223218 316170 223274 316226
rect 223342 316170 223398 316226
rect 222970 316046 223026 316102
rect 223094 316046 223150 316102
rect 223218 316046 223274 316102
rect 223342 316046 223398 316102
rect 222970 315922 223026 315978
rect 223094 315922 223150 315978
rect 223218 315922 223274 315978
rect 223342 315922 223398 315978
rect 222970 298294 223026 298350
rect 223094 298294 223150 298350
rect 223218 298294 223274 298350
rect 223342 298294 223398 298350
rect 222970 298170 223026 298226
rect 223094 298170 223150 298226
rect 223218 298170 223274 298226
rect 223342 298170 223398 298226
rect 222970 298046 223026 298102
rect 223094 298046 223150 298102
rect 223218 298046 223274 298102
rect 223342 298046 223398 298102
rect 222970 297922 223026 297978
rect 223094 297922 223150 297978
rect 223218 297922 223274 297978
rect 223342 297922 223398 297978
rect 222970 280294 223026 280350
rect 223094 280294 223150 280350
rect 223218 280294 223274 280350
rect 223342 280294 223398 280350
rect 222970 280170 223026 280226
rect 223094 280170 223150 280226
rect 223218 280170 223274 280226
rect 223342 280170 223398 280226
rect 222970 280046 223026 280102
rect 223094 280046 223150 280102
rect 223218 280046 223274 280102
rect 223342 280046 223398 280102
rect 222970 279922 223026 279978
rect 223094 279922 223150 279978
rect 223218 279922 223274 279978
rect 223342 279922 223398 279978
rect 222970 262294 223026 262350
rect 223094 262294 223150 262350
rect 223218 262294 223274 262350
rect 223342 262294 223398 262350
rect 222970 262170 223026 262226
rect 223094 262170 223150 262226
rect 223218 262170 223274 262226
rect 223342 262170 223398 262226
rect 222970 262046 223026 262102
rect 223094 262046 223150 262102
rect 223218 262046 223274 262102
rect 223342 262046 223398 262102
rect 222970 261922 223026 261978
rect 223094 261922 223150 261978
rect 223218 261922 223274 261978
rect 223342 261922 223398 261978
rect 222970 244294 223026 244350
rect 223094 244294 223150 244350
rect 223218 244294 223274 244350
rect 223342 244294 223398 244350
rect 222970 244170 223026 244226
rect 223094 244170 223150 244226
rect 223218 244170 223274 244226
rect 223342 244170 223398 244226
rect 222970 244046 223026 244102
rect 223094 244046 223150 244102
rect 223218 244046 223274 244102
rect 223342 244046 223398 244102
rect 222970 243922 223026 243978
rect 223094 243922 223150 243978
rect 223218 243922 223274 243978
rect 223342 243922 223398 243978
rect 237250 597156 237306 597212
rect 237374 597156 237430 597212
rect 237498 597156 237554 597212
rect 237622 597156 237678 597212
rect 237250 597032 237306 597088
rect 237374 597032 237430 597088
rect 237498 597032 237554 597088
rect 237622 597032 237678 597088
rect 237250 596908 237306 596964
rect 237374 596908 237430 596964
rect 237498 596908 237554 596964
rect 237622 596908 237678 596964
rect 237250 596784 237306 596840
rect 237374 596784 237430 596840
rect 237498 596784 237554 596840
rect 237622 596784 237678 596840
rect 237250 580294 237306 580350
rect 237374 580294 237430 580350
rect 237498 580294 237554 580350
rect 237622 580294 237678 580350
rect 237250 580170 237306 580226
rect 237374 580170 237430 580226
rect 237498 580170 237554 580226
rect 237622 580170 237678 580226
rect 237250 580046 237306 580102
rect 237374 580046 237430 580102
rect 237498 580046 237554 580102
rect 237622 580046 237678 580102
rect 237250 579922 237306 579978
rect 237374 579922 237430 579978
rect 237498 579922 237554 579978
rect 237622 579922 237678 579978
rect 237250 562294 237306 562350
rect 237374 562294 237430 562350
rect 237498 562294 237554 562350
rect 237622 562294 237678 562350
rect 237250 562170 237306 562226
rect 237374 562170 237430 562226
rect 237498 562170 237554 562226
rect 237622 562170 237678 562226
rect 237250 562046 237306 562102
rect 237374 562046 237430 562102
rect 237498 562046 237554 562102
rect 237622 562046 237678 562102
rect 237250 561922 237306 561978
rect 237374 561922 237430 561978
rect 237498 561922 237554 561978
rect 237622 561922 237678 561978
rect 237250 544294 237306 544350
rect 237374 544294 237430 544350
rect 237498 544294 237554 544350
rect 237622 544294 237678 544350
rect 237250 544170 237306 544226
rect 237374 544170 237430 544226
rect 237498 544170 237554 544226
rect 237622 544170 237678 544226
rect 237250 544046 237306 544102
rect 237374 544046 237430 544102
rect 237498 544046 237554 544102
rect 237622 544046 237678 544102
rect 237250 543922 237306 543978
rect 237374 543922 237430 543978
rect 237498 543922 237554 543978
rect 237622 543922 237678 543978
rect 237250 526294 237306 526350
rect 237374 526294 237430 526350
rect 237498 526294 237554 526350
rect 237622 526294 237678 526350
rect 237250 526170 237306 526226
rect 237374 526170 237430 526226
rect 237498 526170 237554 526226
rect 237622 526170 237678 526226
rect 237250 526046 237306 526102
rect 237374 526046 237430 526102
rect 237498 526046 237554 526102
rect 237622 526046 237678 526102
rect 237250 525922 237306 525978
rect 237374 525922 237430 525978
rect 237498 525922 237554 525978
rect 237622 525922 237678 525978
rect 237250 508294 237306 508350
rect 237374 508294 237430 508350
rect 237498 508294 237554 508350
rect 237622 508294 237678 508350
rect 237250 508170 237306 508226
rect 237374 508170 237430 508226
rect 237498 508170 237554 508226
rect 237622 508170 237678 508226
rect 237250 508046 237306 508102
rect 237374 508046 237430 508102
rect 237498 508046 237554 508102
rect 237622 508046 237678 508102
rect 237250 507922 237306 507978
rect 237374 507922 237430 507978
rect 237498 507922 237554 507978
rect 237622 507922 237678 507978
rect 237250 490294 237306 490350
rect 237374 490294 237430 490350
rect 237498 490294 237554 490350
rect 237622 490294 237678 490350
rect 237250 490170 237306 490226
rect 237374 490170 237430 490226
rect 237498 490170 237554 490226
rect 237622 490170 237678 490226
rect 237250 490046 237306 490102
rect 237374 490046 237430 490102
rect 237498 490046 237554 490102
rect 237622 490046 237678 490102
rect 237250 489922 237306 489978
rect 237374 489922 237430 489978
rect 237498 489922 237554 489978
rect 237622 489922 237678 489978
rect 237250 472294 237306 472350
rect 237374 472294 237430 472350
rect 237498 472294 237554 472350
rect 237622 472294 237678 472350
rect 237250 472170 237306 472226
rect 237374 472170 237430 472226
rect 237498 472170 237554 472226
rect 237622 472170 237678 472226
rect 237250 472046 237306 472102
rect 237374 472046 237430 472102
rect 237498 472046 237554 472102
rect 237622 472046 237678 472102
rect 237250 471922 237306 471978
rect 237374 471922 237430 471978
rect 237498 471922 237554 471978
rect 237622 471922 237678 471978
rect 237250 454294 237306 454350
rect 237374 454294 237430 454350
rect 237498 454294 237554 454350
rect 237622 454294 237678 454350
rect 237250 454170 237306 454226
rect 237374 454170 237430 454226
rect 237498 454170 237554 454226
rect 237622 454170 237678 454226
rect 237250 454046 237306 454102
rect 237374 454046 237430 454102
rect 237498 454046 237554 454102
rect 237622 454046 237678 454102
rect 237250 453922 237306 453978
rect 237374 453922 237430 453978
rect 237498 453922 237554 453978
rect 237622 453922 237678 453978
rect 237250 436294 237306 436350
rect 237374 436294 237430 436350
rect 237498 436294 237554 436350
rect 237622 436294 237678 436350
rect 237250 436170 237306 436226
rect 237374 436170 237430 436226
rect 237498 436170 237554 436226
rect 237622 436170 237678 436226
rect 237250 436046 237306 436102
rect 237374 436046 237430 436102
rect 237498 436046 237554 436102
rect 237622 436046 237678 436102
rect 237250 435922 237306 435978
rect 237374 435922 237430 435978
rect 237498 435922 237554 435978
rect 237622 435922 237678 435978
rect 237250 418294 237306 418350
rect 237374 418294 237430 418350
rect 237498 418294 237554 418350
rect 237622 418294 237678 418350
rect 237250 418170 237306 418226
rect 237374 418170 237430 418226
rect 237498 418170 237554 418226
rect 237622 418170 237678 418226
rect 237250 418046 237306 418102
rect 237374 418046 237430 418102
rect 237498 418046 237554 418102
rect 237622 418046 237678 418102
rect 237250 417922 237306 417978
rect 237374 417922 237430 417978
rect 237498 417922 237554 417978
rect 237622 417922 237678 417978
rect 237250 400294 237306 400350
rect 237374 400294 237430 400350
rect 237498 400294 237554 400350
rect 237622 400294 237678 400350
rect 237250 400170 237306 400226
rect 237374 400170 237430 400226
rect 237498 400170 237554 400226
rect 237622 400170 237678 400226
rect 237250 400046 237306 400102
rect 237374 400046 237430 400102
rect 237498 400046 237554 400102
rect 237622 400046 237678 400102
rect 237250 399922 237306 399978
rect 237374 399922 237430 399978
rect 237498 399922 237554 399978
rect 237622 399922 237678 399978
rect 237250 382294 237306 382350
rect 237374 382294 237430 382350
rect 237498 382294 237554 382350
rect 237622 382294 237678 382350
rect 237250 382170 237306 382226
rect 237374 382170 237430 382226
rect 237498 382170 237554 382226
rect 237622 382170 237678 382226
rect 237250 382046 237306 382102
rect 237374 382046 237430 382102
rect 237498 382046 237554 382102
rect 237622 382046 237678 382102
rect 237250 381922 237306 381978
rect 237374 381922 237430 381978
rect 237498 381922 237554 381978
rect 237622 381922 237678 381978
rect 237250 364294 237306 364350
rect 237374 364294 237430 364350
rect 237498 364294 237554 364350
rect 237622 364294 237678 364350
rect 237250 364170 237306 364226
rect 237374 364170 237430 364226
rect 237498 364170 237554 364226
rect 237622 364170 237678 364226
rect 237250 364046 237306 364102
rect 237374 364046 237430 364102
rect 237498 364046 237554 364102
rect 237622 364046 237678 364102
rect 237250 363922 237306 363978
rect 237374 363922 237430 363978
rect 237498 363922 237554 363978
rect 237622 363922 237678 363978
rect 237250 346294 237306 346350
rect 237374 346294 237430 346350
rect 237498 346294 237554 346350
rect 237622 346294 237678 346350
rect 237250 346170 237306 346226
rect 237374 346170 237430 346226
rect 237498 346170 237554 346226
rect 237622 346170 237678 346226
rect 237250 346046 237306 346102
rect 237374 346046 237430 346102
rect 237498 346046 237554 346102
rect 237622 346046 237678 346102
rect 237250 345922 237306 345978
rect 237374 345922 237430 345978
rect 237498 345922 237554 345978
rect 237622 345922 237678 345978
rect 237250 328294 237306 328350
rect 237374 328294 237430 328350
rect 237498 328294 237554 328350
rect 237622 328294 237678 328350
rect 237250 328170 237306 328226
rect 237374 328170 237430 328226
rect 237498 328170 237554 328226
rect 237622 328170 237678 328226
rect 237250 328046 237306 328102
rect 237374 328046 237430 328102
rect 237498 328046 237554 328102
rect 237622 328046 237678 328102
rect 237250 327922 237306 327978
rect 237374 327922 237430 327978
rect 237498 327922 237554 327978
rect 237622 327922 237678 327978
rect 237250 310294 237306 310350
rect 237374 310294 237430 310350
rect 237498 310294 237554 310350
rect 237622 310294 237678 310350
rect 237250 310170 237306 310226
rect 237374 310170 237430 310226
rect 237498 310170 237554 310226
rect 237622 310170 237678 310226
rect 237250 310046 237306 310102
rect 237374 310046 237430 310102
rect 237498 310046 237554 310102
rect 237622 310046 237678 310102
rect 237250 309922 237306 309978
rect 237374 309922 237430 309978
rect 237498 309922 237554 309978
rect 237622 309922 237678 309978
rect 237250 292294 237306 292350
rect 237374 292294 237430 292350
rect 237498 292294 237554 292350
rect 237622 292294 237678 292350
rect 237250 292170 237306 292226
rect 237374 292170 237430 292226
rect 237498 292170 237554 292226
rect 237622 292170 237678 292226
rect 237250 292046 237306 292102
rect 237374 292046 237430 292102
rect 237498 292046 237554 292102
rect 237622 292046 237678 292102
rect 237250 291922 237306 291978
rect 237374 291922 237430 291978
rect 237498 291922 237554 291978
rect 237622 291922 237678 291978
rect 237250 274294 237306 274350
rect 237374 274294 237430 274350
rect 237498 274294 237554 274350
rect 237622 274294 237678 274350
rect 237250 274170 237306 274226
rect 237374 274170 237430 274226
rect 237498 274170 237554 274226
rect 237622 274170 237678 274226
rect 237250 274046 237306 274102
rect 237374 274046 237430 274102
rect 237498 274046 237554 274102
rect 237622 274046 237678 274102
rect 237250 273922 237306 273978
rect 237374 273922 237430 273978
rect 237498 273922 237554 273978
rect 237622 273922 237678 273978
rect 237250 256294 237306 256350
rect 237374 256294 237430 256350
rect 237498 256294 237554 256350
rect 237622 256294 237678 256350
rect 237250 256170 237306 256226
rect 237374 256170 237430 256226
rect 237498 256170 237554 256226
rect 237622 256170 237678 256226
rect 237250 256046 237306 256102
rect 237374 256046 237430 256102
rect 237498 256046 237554 256102
rect 237622 256046 237678 256102
rect 237250 255922 237306 255978
rect 237374 255922 237430 255978
rect 237498 255922 237554 255978
rect 237622 255922 237678 255978
rect 237250 238294 237306 238350
rect 237374 238294 237430 238350
rect 237498 238294 237554 238350
rect 237622 238294 237678 238350
rect 237250 238170 237306 238226
rect 237374 238170 237430 238226
rect 237498 238170 237554 238226
rect 237622 238170 237678 238226
rect 237250 238046 237306 238102
rect 237374 238046 237430 238102
rect 237498 238046 237554 238102
rect 237622 238046 237678 238102
rect 237250 237922 237306 237978
rect 237374 237922 237430 237978
rect 237498 237922 237554 237978
rect 237622 237922 237678 237978
rect 222970 226294 223026 226350
rect 223094 226294 223150 226350
rect 223218 226294 223274 226350
rect 223342 226294 223398 226350
rect 222970 226170 223026 226226
rect 223094 226170 223150 226226
rect 223218 226170 223274 226226
rect 223342 226170 223398 226226
rect 222970 226046 223026 226102
rect 223094 226046 223150 226102
rect 223218 226046 223274 226102
rect 223342 226046 223398 226102
rect 222970 225922 223026 225978
rect 223094 225922 223150 225978
rect 223218 225922 223274 225978
rect 223342 225922 223398 225978
rect 233478 226294 233534 226350
rect 233602 226294 233658 226350
rect 233478 226170 233534 226226
rect 233602 226170 233658 226226
rect 233478 226046 233534 226102
rect 233602 226046 233658 226102
rect 233478 225922 233534 225978
rect 233602 225922 233658 225978
rect 237250 220294 237306 220350
rect 237374 220294 237430 220350
rect 237498 220294 237554 220350
rect 237622 220294 237678 220350
rect 237250 220170 237306 220226
rect 237374 220170 237430 220226
rect 237498 220170 237554 220226
rect 237622 220170 237678 220226
rect 237250 220046 237306 220102
rect 237374 220046 237430 220102
rect 237498 220046 237554 220102
rect 237622 220046 237678 220102
rect 237250 219922 237306 219978
rect 237374 219922 237430 219978
rect 237498 219922 237554 219978
rect 237622 219922 237678 219978
rect 240970 598116 241026 598172
rect 241094 598116 241150 598172
rect 241218 598116 241274 598172
rect 241342 598116 241398 598172
rect 240970 597992 241026 598048
rect 241094 597992 241150 598048
rect 241218 597992 241274 598048
rect 241342 597992 241398 598048
rect 240970 597868 241026 597924
rect 241094 597868 241150 597924
rect 241218 597868 241274 597924
rect 241342 597868 241398 597924
rect 240970 597744 241026 597800
rect 241094 597744 241150 597800
rect 241218 597744 241274 597800
rect 241342 597744 241398 597800
rect 240970 586294 241026 586350
rect 241094 586294 241150 586350
rect 241218 586294 241274 586350
rect 241342 586294 241398 586350
rect 240970 586170 241026 586226
rect 241094 586170 241150 586226
rect 241218 586170 241274 586226
rect 241342 586170 241398 586226
rect 240970 586046 241026 586102
rect 241094 586046 241150 586102
rect 241218 586046 241274 586102
rect 241342 586046 241398 586102
rect 240970 585922 241026 585978
rect 241094 585922 241150 585978
rect 241218 585922 241274 585978
rect 241342 585922 241398 585978
rect 240970 568294 241026 568350
rect 241094 568294 241150 568350
rect 241218 568294 241274 568350
rect 241342 568294 241398 568350
rect 240970 568170 241026 568226
rect 241094 568170 241150 568226
rect 241218 568170 241274 568226
rect 241342 568170 241398 568226
rect 240970 568046 241026 568102
rect 241094 568046 241150 568102
rect 241218 568046 241274 568102
rect 241342 568046 241398 568102
rect 240970 567922 241026 567978
rect 241094 567922 241150 567978
rect 241218 567922 241274 567978
rect 241342 567922 241398 567978
rect 240970 550294 241026 550350
rect 241094 550294 241150 550350
rect 241218 550294 241274 550350
rect 241342 550294 241398 550350
rect 240970 550170 241026 550226
rect 241094 550170 241150 550226
rect 241218 550170 241274 550226
rect 241342 550170 241398 550226
rect 240970 550046 241026 550102
rect 241094 550046 241150 550102
rect 241218 550046 241274 550102
rect 241342 550046 241398 550102
rect 240970 549922 241026 549978
rect 241094 549922 241150 549978
rect 241218 549922 241274 549978
rect 241342 549922 241398 549978
rect 240970 532294 241026 532350
rect 241094 532294 241150 532350
rect 241218 532294 241274 532350
rect 241342 532294 241398 532350
rect 240970 532170 241026 532226
rect 241094 532170 241150 532226
rect 241218 532170 241274 532226
rect 241342 532170 241398 532226
rect 240970 532046 241026 532102
rect 241094 532046 241150 532102
rect 241218 532046 241274 532102
rect 241342 532046 241398 532102
rect 240970 531922 241026 531978
rect 241094 531922 241150 531978
rect 241218 531922 241274 531978
rect 241342 531922 241398 531978
rect 240970 514294 241026 514350
rect 241094 514294 241150 514350
rect 241218 514294 241274 514350
rect 241342 514294 241398 514350
rect 240970 514170 241026 514226
rect 241094 514170 241150 514226
rect 241218 514170 241274 514226
rect 241342 514170 241398 514226
rect 240970 514046 241026 514102
rect 241094 514046 241150 514102
rect 241218 514046 241274 514102
rect 241342 514046 241398 514102
rect 240970 513922 241026 513978
rect 241094 513922 241150 513978
rect 241218 513922 241274 513978
rect 241342 513922 241398 513978
rect 240970 496294 241026 496350
rect 241094 496294 241150 496350
rect 241218 496294 241274 496350
rect 241342 496294 241398 496350
rect 240970 496170 241026 496226
rect 241094 496170 241150 496226
rect 241218 496170 241274 496226
rect 241342 496170 241398 496226
rect 240970 496046 241026 496102
rect 241094 496046 241150 496102
rect 241218 496046 241274 496102
rect 241342 496046 241398 496102
rect 240970 495922 241026 495978
rect 241094 495922 241150 495978
rect 241218 495922 241274 495978
rect 241342 495922 241398 495978
rect 240970 478294 241026 478350
rect 241094 478294 241150 478350
rect 241218 478294 241274 478350
rect 241342 478294 241398 478350
rect 240970 478170 241026 478226
rect 241094 478170 241150 478226
rect 241218 478170 241274 478226
rect 241342 478170 241398 478226
rect 240970 478046 241026 478102
rect 241094 478046 241150 478102
rect 241218 478046 241274 478102
rect 241342 478046 241398 478102
rect 240970 477922 241026 477978
rect 241094 477922 241150 477978
rect 241218 477922 241274 477978
rect 241342 477922 241398 477978
rect 240970 460294 241026 460350
rect 241094 460294 241150 460350
rect 241218 460294 241274 460350
rect 241342 460294 241398 460350
rect 240970 460170 241026 460226
rect 241094 460170 241150 460226
rect 241218 460170 241274 460226
rect 241342 460170 241398 460226
rect 240970 460046 241026 460102
rect 241094 460046 241150 460102
rect 241218 460046 241274 460102
rect 241342 460046 241398 460102
rect 240970 459922 241026 459978
rect 241094 459922 241150 459978
rect 241218 459922 241274 459978
rect 241342 459922 241398 459978
rect 240970 442294 241026 442350
rect 241094 442294 241150 442350
rect 241218 442294 241274 442350
rect 241342 442294 241398 442350
rect 240970 442170 241026 442226
rect 241094 442170 241150 442226
rect 241218 442170 241274 442226
rect 241342 442170 241398 442226
rect 240970 442046 241026 442102
rect 241094 442046 241150 442102
rect 241218 442046 241274 442102
rect 241342 442046 241398 442102
rect 240970 441922 241026 441978
rect 241094 441922 241150 441978
rect 241218 441922 241274 441978
rect 241342 441922 241398 441978
rect 240970 424294 241026 424350
rect 241094 424294 241150 424350
rect 241218 424294 241274 424350
rect 241342 424294 241398 424350
rect 240970 424170 241026 424226
rect 241094 424170 241150 424226
rect 241218 424170 241274 424226
rect 241342 424170 241398 424226
rect 240970 424046 241026 424102
rect 241094 424046 241150 424102
rect 241218 424046 241274 424102
rect 241342 424046 241398 424102
rect 240970 423922 241026 423978
rect 241094 423922 241150 423978
rect 241218 423922 241274 423978
rect 241342 423922 241398 423978
rect 240970 406294 241026 406350
rect 241094 406294 241150 406350
rect 241218 406294 241274 406350
rect 241342 406294 241398 406350
rect 240970 406170 241026 406226
rect 241094 406170 241150 406226
rect 241218 406170 241274 406226
rect 241342 406170 241398 406226
rect 240970 406046 241026 406102
rect 241094 406046 241150 406102
rect 241218 406046 241274 406102
rect 241342 406046 241398 406102
rect 240970 405922 241026 405978
rect 241094 405922 241150 405978
rect 241218 405922 241274 405978
rect 241342 405922 241398 405978
rect 240970 388294 241026 388350
rect 241094 388294 241150 388350
rect 241218 388294 241274 388350
rect 241342 388294 241398 388350
rect 240970 388170 241026 388226
rect 241094 388170 241150 388226
rect 241218 388170 241274 388226
rect 241342 388170 241398 388226
rect 240970 388046 241026 388102
rect 241094 388046 241150 388102
rect 241218 388046 241274 388102
rect 241342 388046 241398 388102
rect 240970 387922 241026 387978
rect 241094 387922 241150 387978
rect 241218 387922 241274 387978
rect 241342 387922 241398 387978
rect 240970 370294 241026 370350
rect 241094 370294 241150 370350
rect 241218 370294 241274 370350
rect 241342 370294 241398 370350
rect 240970 370170 241026 370226
rect 241094 370170 241150 370226
rect 241218 370170 241274 370226
rect 241342 370170 241398 370226
rect 240970 370046 241026 370102
rect 241094 370046 241150 370102
rect 241218 370046 241274 370102
rect 241342 370046 241398 370102
rect 240970 369922 241026 369978
rect 241094 369922 241150 369978
rect 241218 369922 241274 369978
rect 241342 369922 241398 369978
rect 240970 352294 241026 352350
rect 241094 352294 241150 352350
rect 241218 352294 241274 352350
rect 241342 352294 241398 352350
rect 240970 352170 241026 352226
rect 241094 352170 241150 352226
rect 241218 352170 241274 352226
rect 241342 352170 241398 352226
rect 240970 352046 241026 352102
rect 241094 352046 241150 352102
rect 241218 352046 241274 352102
rect 241342 352046 241398 352102
rect 240970 351922 241026 351978
rect 241094 351922 241150 351978
rect 241218 351922 241274 351978
rect 241342 351922 241398 351978
rect 240970 334294 241026 334350
rect 241094 334294 241150 334350
rect 241218 334294 241274 334350
rect 241342 334294 241398 334350
rect 240970 334170 241026 334226
rect 241094 334170 241150 334226
rect 241218 334170 241274 334226
rect 241342 334170 241398 334226
rect 240970 334046 241026 334102
rect 241094 334046 241150 334102
rect 241218 334046 241274 334102
rect 241342 334046 241398 334102
rect 240970 333922 241026 333978
rect 241094 333922 241150 333978
rect 241218 333922 241274 333978
rect 241342 333922 241398 333978
rect 240970 316294 241026 316350
rect 241094 316294 241150 316350
rect 241218 316294 241274 316350
rect 241342 316294 241398 316350
rect 240970 316170 241026 316226
rect 241094 316170 241150 316226
rect 241218 316170 241274 316226
rect 241342 316170 241398 316226
rect 240970 316046 241026 316102
rect 241094 316046 241150 316102
rect 241218 316046 241274 316102
rect 241342 316046 241398 316102
rect 240970 315922 241026 315978
rect 241094 315922 241150 315978
rect 241218 315922 241274 315978
rect 241342 315922 241398 315978
rect 240970 298294 241026 298350
rect 241094 298294 241150 298350
rect 241218 298294 241274 298350
rect 241342 298294 241398 298350
rect 240970 298170 241026 298226
rect 241094 298170 241150 298226
rect 241218 298170 241274 298226
rect 241342 298170 241398 298226
rect 240970 298046 241026 298102
rect 241094 298046 241150 298102
rect 241218 298046 241274 298102
rect 241342 298046 241398 298102
rect 240970 297922 241026 297978
rect 241094 297922 241150 297978
rect 241218 297922 241274 297978
rect 241342 297922 241398 297978
rect 240970 280294 241026 280350
rect 241094 280294 241150 280350
rect 241218 280294 241274 280350
rect 241342 280294 241398 280350
rect 240970 280170 241026 280226
rect 241094 280170 241150 280226
rect 241218 280170 241274 280226
rect 241342 280170 241398 280226
rect 240970 280046 241026 280102
rect 241094 280046 241150 280102
rect 241218 280046 241274 280102
rect 241342 280046 241398 280102
rect 240970 279922 241026 279978
rect 241094 279922 241150 279978
rect 241218 279922 241274 279978
rect 241342 279922 241398 279978
rect 240970 262294 241026 262350
rect 241094 262294 241150 262350
rect 241218 262294 241274 262350
rect 241342 262294 241398 262350
rect 240970 262170 241026 262226
rect 241094 262170 241150 262226
rect 241218 262170 241274 262226
rect 241342 262170 241398 262226
rect 240970 262046 241026 262102
rect 241094 262046 241150 262102
rect 241218 262046 241274 262102
rect 241342 262046 241398 262102
rect 240970 261922 241026 261978
rect 241094 261922 241150 261978
rect 241218 261922 241274 261978
rect 241342 261922 241398 261978
rect 240970 244294 241026 244350
rect 241094 244294 241150 244350
rect 241218 244294 241274 244350
rect 241342 244294 241398 244350
rect 240970 244170 241026 244226
rect 241094 244170 241150 244226
rect 241218 244170 241274 244226
rect 241342 244170 241398 244226
rect 240970 244046 241026 244102
rect 241094 244046 241150 244102
rect 241218 244046 241274 244102
rect 241342 244046 241398 244102
rect 240970 243922 241026 243978
rect 241094 243922 241150 243978
rect 241218 243922 241274 243978
rect 241342 243922 241398 243978
rect 258970 598116 259026 598172
rect 259094 598116 259150 598172
rect 259218 598116 259274 598172
rect 259342 598116 259398 598172
rect 258970 597992 259026 598048
rect 259094 597992 259150 598048
rect 259218 597992 259274 598048
rect 259342 597992 259398 598048
rect 258970 597868 259026 597924
rect 259094 597868 259150 597924
rect 259218 597868 259274 597924
rect 259342 597868 259398 597924
rect 258970 597744 259026 597800
rect 259094 597744 259150 597800
rect 259218 597744 259274 597800
rect 259342 597744 259398 597800
rect 258970 586294 259026 586350
rect 259094 586294 259150 586350
rect 259218 586294 259274 586350
rect 259342 586294 259398 586350
rect 258970 586170 259026 586226
rect 259094 586170 259150 586226
rect 259218 586170 259274 586226
rect 259342 586170 259398 586226
rect 258970 586046 259026 586102
rect 259094 586046 259150 586102
rect 259218 586046 259274 586102
rect 259342 586046 259398 586102
rect 258970 585922 259026 585978
rect 259094 585922 259150 585978
rect 259218 585922 259274 585978
rect 259342 585922 259398 585978
rect 258970 568294 259026 568350
rect 259094 568294 259150 568350
rect 259218 568294 259274 568350
rect 259342 568294 259398 568350
rect 258970 568170 259026 568226
rect 259094 568170 259150 568226
rect 259218 568170 259274 568226
rect 259342 568170 259398 568226
rect 258970 568046 259026 568102
rect 259094 568046 259150 568102
rect 259218 568046 259274 568102
rect 259342 568046 259398 568102
rect 258970 567922 259026 567978
rect 259094 567922 259150 567978
rect 259218 567922 259274 567978
rect 259342 567922 259398 567978
rect 258970 550294 259026 550350
rect 259094 550294 259150 550350
rect 259218 550294 259274 550350
rect 259342 550294 259398 550350
rect 258970 550170 259026 550226
rect 259094 550170 259150 550226
rect 259218 550170 259274 550226
rect 259342 550170 259398 550226
rect 258970 550046 259026 550102
rect 259094 550046 259150 550102
rect 259218 550046 259274 550102
rect 259342 550046 259398 550102
rect 258970 549922 259026 549978
rect 259094 549922 259150 549978
rect 259218 549922 259274 549978
rect 259342 549922 259398 549978
rect 258970 532294 259026 532350
rect 259094 532294 259150 532350
rect 259218 532294 259274 532350
rect 259342 532294 259398 532350
rect 258970 532170 259026 532226
rect 259094 532170 259150 532226
rect 259218 532170 259274 532226
rect 259342 532170 259398 532226
rect 258970 532046 259026 532102
rect 259094 532046 259150 532102
rect 259218 532046 259274 532102
rect 259342 532046 259398 532102
rect 258970 531922 259026 531978
rect 259094 531922 259150 531978
rect 259218 531922 259274 531978
rect 259342 531922 259398 531978
rect 258970 514294 259026 514350
rect 259094 514294 259150 514350
rect 259218 514294 259274 514350
rect 259342 514294 259398 514350
rect 258970 514170 259026 514226
rect 259094 514170 259150 514226
rect 259218 514170 259274 514226
rect 259342 514170 259398 514226
rect 258970 514046 259026 514102
rect 259094 514046 259150 514102
rect 259218 514046 259274 514102
rect 259342 514046 259398 514102
rect 258970 513922 259026 513978
rect 259094 513922 259150 513978
rect 259218 513922 259274 513978
rect 259342 513922 259398 513978
rect 258970 496294 259026 496350
rect 259094 496294 259150 496350
rect 259218 496294 259274 496350
rect 259342 496294 259398 496350
rect 258970 496170 259026 496226
rect 259094 496170 259150 496226
rect 259218 496170 259274 496226
rect 259342 496170 259398 496226
rect 258970 496046 259026 496102
rect 259094 496046 259150 496102
rect 259218 496046 259274 496102
rect 259342 496046 259398 496102
rect 258970 495922 259026 495978
rect 259094 495922 259150 495978
rect 259218 495922 259274 495978
rect 259342 495922 259398 495978
rect 258970 478294 259026 478350
rect 259094 478294 259150 478350
rect 259218 478294 259274 478350
rect 259342 478294 259398 478350
rect 258970 478170 259026 478226
rect 259094 478170 259150 478226
rect 259218 478170 259274 478226
rect 259342 478170 259398 478226
rect 258970 478046 259026 478102
rect 259094 478046 259150 478102
rect 259218 478046 259274 478102
rect 259342 478046 259398 478102
rect 258970 477922 259026 477978
rect 259094 477922 259150 477978
rect 259218 477922 259274 477978
rect 259342 477922 259398 477978
rect 258970 460294 259026 460350
rect 259094 460294 259150 460350
rect 259218 460294 259274 460350
rect 259342 460294 259398 460350
rect 258970 460170 259026 460226
rect 259094 460170 259150 460226
rect 259218 460170 259274 460226
rect 259342 460170 259398 460226
rect 258970 460046 259026 460102
rect 259094 460046 259150 460102
rect 259218 460046 259274 460102
rect 259342 460046 259398 460102
rect 258970 459922 259026 459978
rect 259094 459922 259150 459978
rect 259218 459922 259274 459978
rect 259342 459922 259398 459978
rect 258970 442294 259026 442350
rect 259094 442294 259150 442350
rect 259218 442294 259274 442350
rect 259342 442294 259398 442350
rect 258970 442170 259026 442226
rect 259094 442170 259150 442226
rect 259218 442170 259274 442226
rect 259342 442170 259398 442226
rect 258970 442046 259026 442102
rect 259094 442046 259150 442102
rect 259218 442046 259274 442102
rect 259342 442046 259398 442102
rect 258970 441922 259026 441978
rect 259094 441922 259150 441978
rect 259218 441922 259274 441978
rect 259342 441922 259398 441978
rect 258970 424294 259026 424350
rect 259094 424294 259150 424350
rect 259218 424294 259274 424350
rect 259342 424294 259398 424350
rect 258970 424170 259026 424226
rect 259094 424170 259150 424226
rect 259218 424170 259274 424226
rect 259342 424170 259398 424226
rect 258970 424046 259026 424102
rect 259094 424046 259150 424102
rect 259218 424046 259274 424102
rect 259342 424046 259398 424102
rect 258970 423922 259026 423978
rect 259094 423922 259150 423978
rect 259218 423922 259274 423978
rect 259342 423922 259398 423978
rect 258970 406294 259026 406350
rect 259094 406294 259150 406350
rect 259218 406294 259274 406350
rect 259342 406294 259398 406350
rect 258970 406170 259026 406226
rect 259094 406170 259150 406226
rect 259218 406170 259274 406226
rect 259342 406170 259398 406226
rect 258970 406046 259026 406102
rect 259094 406046 259150 406102
rect 259218 406046 259274 406102
rect 259342 406046 259398 406102
rect 258970 405922 259026 405978
rect 259094 405922 259150 405978
rect 259218 405922 259274 405978
rect 259342 405922 259398 405978
rect 258970 388294 259026 388350
rect 259094 388294 259150 388350
rect 259218 388294 259274 388350
rect 259342 388294 259398 388350
rect 258970 388170 259026 388226
rect 259094 388170 259150 388226
rect 259218 388170 259274 388226
rect 259342 388170 259398 388226
rect 258970 388046 259026 388102
rect 259094 388046 259150 388102
rect 259218 388046 259274 388102
rect 259342 388046 259398 388102
rect 258970 387922 259026 387978
rect 259094 387922 259150 387978
rect 259218 387922 259274 387978
rect 259342 387922 259398 387978
rect 258970 370294 259026 370350
rect 259094 370294 259150 370350
rect 259218 370294 259274 370350
rect 259342 370294 259398 370350
rect 258970 370170 259026 370226
rect 259094 370170 259150 370226
rect 259218 370170 259274 370226
rect 259342 370170 259398 370226
rect 258970 370046 259026 370102
rect 259094 370046 259150 370102
rect 259218 370046 259274 370102
rect 259342 370046 259398 370102
rect 258970 369922 259026 369978
rect 259094 369922 259150 369978
rect 259218 369922 259274 369978
rect 259342 369922 259398 369978
rect 258970 352294 259026 352350
rect 259094 352294 259150 352350
rect 259218 352294 259274 352350
rect 259342 352294 259398 352350
rect 258970 352170 259026 352226
rect 259094 352170 259150 352226
rect 259218 352170 259274 352226
rect 259342 352170 259398 352226
rect 258970 352046 259026 352102
rect 259094 352046 259150 352102
rect 259218 352046 259274 352102
rect 259342 352046 259398 352102
rect 258970 351922 259026 351978
rect 259094 351922 259150 351978
rect 259218 351922 259274 351978
rect 259342 351922 259398 351978
rect 258970 334294 259026 334350
rect 259094 334294 259150 334350
rect 259218 334294 259274 334350
rect 259342 334294 259398 334350
rect 258970 334170 259026 334226
rect 259094 334170 259150 334226
rect 259218 334170 259274 334226
rect 259342 334170 259398 334226
rect 258970 334046 259026 334102
rect 259094 334046 259150 334102
rect 259218 334046 259274 334102
rect 259342 334046 259398 334102
rect 258970 333922 259026 333978
rect 259094 333922 259150 333978
rect 259218 333922 259274 333978
rect 259342 333922 259398 333978
rect 258970 316294 259026 316350
rect 259094 316294 259150 316350
rect 259218 316294 259274 316350
rect 259342 316294 259398 316350
rect 258970 316170 259026 316226
rect 259094 316170 259150 316226
rect 259218 316170 259274 316226
rect 259342 316170 259398 316226
rect 258970 316046 259026 316102
rect 259094 316046 259150 316102
rect 259218 316046 259274 316102
rect 259342 316046 259398 316102
rect 258970 315922 259026 315978
rect 259094 315922 259150 315978
rect 259218 315922 259274 315978
rect 259342 315922 259398 315978
rect 258970 298294 259026 298350
rect 259094 298294 259150 298350
rect 259218 298294 259274 298350
rect 259342 298294 259398 298350
rect 258970 298170 259026 298226
rect 259094 298170 259150 298226
rect 259218 298170 259274 298226
rect 259342 298170 259398 298226
rect 258970 298046 259026 298102
rect 259094 298046 259150 298102
rect 259218 298046 259274 298102
rect 259342 298046 259398 298102
rect 258970 297922 259026 297978
rect 259094 297922 259150 297978
rect 259218 297922 259274 297978
rect 259342 297922 259398 297978
rect 258970 280294 259026 280350
rect 259094 280294 259150 280350
rect 259218 280294 259274 280350
rect 259342 280294 259398 280350
rect 258970 280170 259026 280226
rect 259094 280170 259150 280226
rect 259218 280170 259274 280226
rect 259342 280170 259398 280226
rect 258970 280046 259026 280102
rect 259094 280046 259150 280102
rect 259218 280046 259274 280102
rect 259342 280046 259398 280102
rect 258970 279922 259026 279978
rect 259094 279922 259150 279978
rect 259218 279922 259274 279978
rect 259342 279922 259398 279978
rect 258970 262294 259026 262350
rect 259094 262294 259150 262350
rect 259218 262294 259274 262350
rect 259342 262294 259398 262350
rect 258970 262170 259026 262226
rect 259094 262170 259150 262226
rect 259218 262170 259274 262226
rect 259342 262170 259398 262226
rect 258970 262046 259026 262102
rect 259094 262046 259150 262102
rect 259218 262046 259274 262102
rect 259342 262046 259398 262102
rect 258970 261922 259026 261978
rect 259094 261922 259150 261978
rect 259218 261922 259274 261978
rect 259342 261922 259398 261978
rect 258970 244294 259026 244350
rect 259094 244294 259150 244350
rect 259218 244294 259274 244350
rect 259342 244294 259398 244350
rect 258970 244170 259026 244226
rect 259094 244170 259150 244226
rect 259218 244170 259274 244226
rect 259342 244170 259398 244226
rect 258970 244046 259026 244102
rect 259094 244046 259150 244102
rect 259218 244046 259274 244102
rect 259342 244046 259398 244102
rect 258970 243922 259026 243978
rect 259094 243922 259150 243978
rect 259218 243922 259274 243978
rect 259342 243922 259398 243978
rect 240970 226294 241026 226350
rect 241094 226294 241150 226350
rect 241218 226294 241274 226350
rect 241342 226294 241398 226350
rect 240970 226170 241026 226226
rect 241094 226170 241150 226226
rect 241218 226170 241274 226226
rect 241342 226170 241398 226226
rect 240970 226046 241026 226102
rect 241094 226046 241150 226102
rect 241218 226046 241274 226102
rect 241342 226046 241398 226102
rect 240970 225922 241026 225978
rect 241094 225922 241150 225978
rect 241218 225922 241274 225978
rect 241342 225922 241398 225978
rect 79878 208294 79934 208350
rect 80002 208294 80058 208350
rect 79878 208170 79934 208226
rect 80002 208170 80058 208226
rect 79878 208046 79934 208102
rect 80002 208046 80058 208102
rect 79878 207922 79934 207978
rect 80002 207922 80058 207978
rect 110598 208294 110654 208350
rect 110722 208294 110778 208350
rect 110598 208170 110654 208226
rect 110722 208170 110778 208226
rect 110598 208046 110654 208102
rect 110722 208046 110778 208102
rect 110598 207922 110654 207978
rect 110722 207922 110778 207978
rect 141318 208294 141374 208350
rect 141442 208294 141498 208350
rect 141318 208170 141374 208226
rect 141442 208170 141498 208226
rect 141318 208046 141374 208102
rect 141442 208046 141498 208102
rect 141318 207922 141374 207978
rect 141442 207922 141498 207978
rect 172038 208294 172094 208350
rect 172162 208294 172218 208350
rect 172038 208170 172094 208226
rect 172162 208170 172218 208226
rect 172038 208046 172094 208102
rect 172162 208046 172218 208102
rect 172038 207922 172094 207978
rect 172162 207922 172218 207978
rect 202758 208294 202814 208350
rect 202882 208294 202938 208350
rect 202758 208170 202814 208226
rect 202882 208170 202938 208226
rect 202758 208046 202814 208102
rect 202882 208046 202938 208102
rect 202758 207922 202814 207978
rect 202882 207922 202938 207978
rect 233478 208294 233534 208350
rect 233602 208294 233658 208350
rect 233478 208170 233534 208226
rect 233602 208170 233658 208226
rect 233478 208046 233534 208102
rect 233602 208046 233658 208102
rect 233478 207922 233534 207978
rect 233602 207922 233658 207978
rect 255250 238294 255306 238350
rect 255374 238294 255430 238350
rect 255498 238294 255554 238350
rect 255622 238294 255678 238350
rect 255250 238170 255306 238226
rect 255374 238170 255430 238226
rect 255498 238170 255554 238226
rect 255622 238170 255678 238226
rect 255250 238046 255306 238102
rect 255374 238046 255430 238102
rect 255498 238046 255554 238102
rect 255622 238046 255678 238102
rect 255250 237922 255306 237978
rect 255374 237922 255430 237978
rect 255498 237922 255554 237978
rect 255622 237922 255678 237978
rect 255250 220294 255306 220350
rect 255374 220294 255430 220350
rect 255498 220294 255554 220350
rect 255622 220294 255678 220350
rect 255250 220170 255306 220226
rect 255374 220170 255430 220226
rect 255498 220170 255554 220226
rect 255622 220170 255678 220226
rect 255250 220046 255306 220102
rect 255374 220046 255430 220102
rect 255498 220046 255554 220102
rect 255622 220046 255678 220102
rect 255250 219922 255306 219978
rect 255374 219922 255430 219978
rect 255498 219922 255554 219978
rect 255622 219922 255678 219978
rect 240970 208294 241026 208350
rect 241094 208294 241150 208350
rect 241218 208294 241274 208350
rect 241342 208294 241398 208350
rect 240970 208170 241026 208226
rect 241094 208170 241150 208226
rect 241218 208170 241274 208226
rect 241342 208170 241398 208226
rect 240970 208046 241026 208102
rect 241094 208046 241150 208102
rect 241218 208046 241274 208102
rect 241342 208046 241398 208102
rect 240970 207922 241026 207978
rect 241094 207922 241150 207978
rect 241218 207922 241274 207978
rect 241342 207922 241398 207978
rect 57250 202294 57306 202350
rect 57374 202294 57430 202350
rect 57498 202294 57554 202350
rect 57622 202294 57678 202350
rect 57250 202170 57306 202226
rect 57374 202170 57430 202226
rect 57498 202170 57554 202226
rect 57622 202170 57678 202226
rect 57250 202046 57306 202102
rect 57374 202046 57430 202102
rect 57498 202046 57554 202102
rect 57622 202046 57678 202102
rect 57250 201922 57306 201978
rect 57374 201922 57430 201978
rect 57498 201922 57554 201978
rect 57622 201922 57678 201978
rect 64518 202294 64574 202350
rect 64642 202294 64698 202350
rect 64518 202170 64574 202226
rect 64642 202170 64698 202226
rect 64518 202046 64574 202102
rect 64642 202046 64698 202102
rect 64518 201922 64574 201978
rect 64642 201922 64698 201978
rect 95238 202294 95294 202350
rect 95362 202294 95418 202350
rect 95238 202170 95294 202226
rect 95362 202170 95418 202226
rect 95238 202046 95294 202102
rect 95362 202046 95418 202102
rect 95238 201922 95294 201978
rect 95362 201922 95418 201978
rect 125958 202294 126014 202350
rect 126082 202294 126138 202350
rect 125958 202170 126014 202226
rect 126082 202170 126138 202226
rect 125958 202046 126014 202102
rect 126082 202046 126138 202102
rect 125958 201922 126014 201978
rect 126082 201922 126138 201978
rect 156678 202294 156734 202350
rect 156802 202294 156858 202350
rect 156678 202170 156734 202226
rect 156802 202170 156858 202226
rect 156678 202046 156734 202102
rect 156802 202046 156858 202102
rect 156678 201922 156734 201978
rect 156802 201922 156858 201978
rect 187398 202294 187454 202350
rect 187522 202294 187578 202350
rect 187398 202170 187454 202226
rect 187522 202170 187578 202226
rect 187398 202046 187454 202102
rect 187522 202046 187578 202102
rect 187398 201922 187454 201978
rect 187522 201922 187578 201978
rect 218118 202294 218174 202350
rect 218242 202294 218298 202350
rect 218118 202170 218174 202226
rect 218242 202170 218298 202226
rect 218118 202046 218174 202102
rect 218242 202046 218298 202102
rect 218118 201922 218174 201978
rect 218242 201922 218298 201978
rect 240970 190294 241026 190350
rect 241094 190294 241150 190350
rect 241218 190294 241274 190350
rect 241342 190294 241398 190350
rect 240970 190170 241026 190226
rect 241094 190170 241150 190226
rect 241218 190170 241274 190226
rect 241342 190170 241398 190226
rect 240970 190046 241026 190102
rect 241094 190046 241150 190102
rect 241218 190046 241274 190102
rect 241342 190046 241398 190102
rect 240970 189922 241026 189978
rect 241094 189922 241150 189978
rect 241218 189922 241274 189978
rect 241342 189922 241398 189978
rect 57250 184294 57306 184350
rect 57374 184294 57430 184350
rect 57498 184294 57554 184350
rect 57622 184294 57678 184350
rect 57250 184170 57306 184226
rect 57374 184170 57430 184226
rect 57498 184170 57554 184226
rect 57622 184170 57678 184226
rect 57250 184046 57306 184102
rect 57374 184046 57430 184102
rect 57498 184046 57554 184102
rect 57622 184046 57678 184102
rect 57250 183922 57306 183978
rect 57374 183922 57430 183978
rect 57498 183922 57554 183978
rect 57622 183922 57678 183978
rect 64518 184294 64574 184350
rect 64642 184294 64698 184350
rect 64518 184170 64574 184226
rect 64642 184170 64698 184226
rect 64518 184046 64574 184102
rect 64642 184046 64698 184102
rect 64518 183922 64574 183978
rect 64642 183922 64698 183978
rect 240970 172294 241026 172350
rect 241094 172294 241150 172350
rect 241218 172294 241274 172350
rect 241342 172294 241398 172350
rect 240970 172170 241026 172226
rect 241094 172170 241150 172226
rect 241218 172170 241274 172226
rect 241342 172170 241398 172226
rect 240970 172046 241026 172102
rect 241094 172046 241150 172102
rect 241218 172046 241274 172102
rect 241342 172046 241398 172102
rect 240970 171922 241026 171978
rect 241094 171922 241150 171978
rect 241218 171922 241274 171978
rect 241342 171922 241398 171978
rect 57250 166294 57306 166350
rect 57374 166294 57430 166350
rect 57498 166294 57554 166350
rect 57622 166294 57678 166350
rect 57250 166170 57306 166226
rect 57374 166170 57430 166226
rect 57498 166170 57554 166226
rect 57622 166170 57678 166226
rect 57250 166046 57306 166102
rect 57374 166046 57430 166102
rect 57498 166046 57554 166102
rect 57622 166046 57678 166102
rect 57250 165922 57306 165978
rect 57374 165922 57430 165978
rect 57498 165922 57554 165978
rect 57622 165922 57678 165978
rect 64518 166294 64574 166350
rect 64642 166294 64698 166350
rect 64518 166170 64574 166226
rect 64642 166170 64698 166226
rect 64518 166046 64574 166102
rect 64642 166046 64698 166102
rect 64518 165922 64574 165978
rect 64642 165922 64698 165978
rect 240970 154294 241026 154350
rect 241094 154294 241150 154350
rect 241218 154294 241274 154350
rect 241342 154294 241398 154350
rect 240970 154170 241026 154226
rect 241094 154170 241150 154226
rect 241218 154170 241274 154226
rect 241342 154170 241398 154226
rect 240970 154046 241026 154102
rect 241094 154046 241150 154102
rect 241218 154046 241274 154102
rect 241342 154046 241398 154102
rect 240970 153922 241026 153978
rect 241094 153922 241150 153978
rect 241218 153922 241274 153978
rect 241342 153922 241398 153978
rect 57250 148294 57306 148350
rect 57374 148294 57430 148350
rect 57498 148294 57554 148350
rect 57622 148294 57678 148350
rect 57250 148170 57306 148226
rect 57374 148170 57430 148226
rect 57498 148170 57554 148226
rect 57622 148170 57678 148226
rect 57250 148046 57306 148102
rect 57374 148046 57430 148102
rect 57498 148046 57554 148102
rect 57622 148046 57678 148102
rect 57250 147922 57306 147978
rect 57374 147922 57430 147978
rect 57498 147922 57554 147978
rect 57622 147922 57678 147978
rect 64518 148294 64574 148350
rect 64642 148294 64698 148350
rect 64518 148170 64574 148226
rect 64642 148170 64698 148226
rect 64518 148046 64574 148102
rect 64642 148046 64698 148102
rect 64518 147922 64574 147978
rect 64642 147922 64698 147978
rect 240970 136294 241026 136350
rect 241094 136294 241150 136350
rect 241218 136294 241274 136350
rect 241342 136294 241398 136350
rect 240970 136170 241026 136226
rect 241094 136170 241150 136226
rect 241218 136170 241274 136226
rect 241342 136170 241398 136226
rect 240970 136046 241026 136102
rect 241094 136046 241150 136102
rect 241218 136046 241274 136102
rect 241342 136046 241398 136102
rect 240970 135922 241026 135978
rect 241094 135922 241150 135978
rect 241218 135922 241274 135978
rect 241342 135922 241398 135978
rect 57250 130294 57306 130350
rect 57374 130294 57430 130350
rect 57498 130294 57554 130350
rect 57622 130294 57678 130350
rect 57250 130170 57306 130226
rect 57374 130170 57430 130226
rect 57498 130170 57554 130226
rect 57622 130170 57678 130226
rect 57250 130046 57306 130102
rect 57374 130046 57430 130102
rect 57498 130046 57554 130102
rect 57622 130046 57678 130102
rect 57250 129922 57306 129978
rect 57374 129922 57430 129978
rect 57498 129922 57554 129978
rect 57622 129922 57678 129978
rect 64518 130294 64574 130350
rect 64642 130294 64698 130350
rect 64518 130170 64574 130226
rect 64642 130170 64698 130226
rect 64518 130046 64574 130102
rect 64642 130046 64698 130102
rect 64518 129922 64574 129978
rect 64642 129922 64698 129978
rect 240970 118294 241026 118350
rect 241094 118294 241150 118350
rect 241218 118294 241274 118350
rect 241342 118294 241398 118350
rect 240970 118170 241026 118226
rect 241094 118170 241150 118226
rect 241218 118170 241274 118226
rect 241342 118170 241398 118226
rect 240970 118046 241026 118102
rect 241094 118046 241150 118102
rect 241218 118046 241274 118102
rect 241342 118046 241398 118102
rect 240970 117922 241026 117978
rect 241094 117922 241150 117978
rect 241218 117922 241274 117978
rect 241342 117922 241398 117978
rect 57250 112294 57306 112350
rect 57374 112294 57430 112350
rect 57498 112294 57554 112350
rect 57622 112294 57678 112350
rect 57250 112170 57306 112226
rect 57374 112170 57430 112226
rect 57498 112170 57554 112226
rect 57622 112170 57678 112226
rect 57250 112046 57306 112102
rect 57374 112046 57430 112102
rect 57498 112046 57554 112102
rect 57622 112046 57678 112102
rect 57250 111922 57306 111978
rect 57374 111922 57430 111978
rect 57498 111922 57554 111978
rect 57622 111922 57678 111978
rect 64518 112294 64574 112350
rect 64642 112294 64698 112350
rect 64518 112170 64574 112226
rect 64642 112170 64698 112226
rect 64518 112046 64574 112102
rect 64642 112046 64698 112102
rect 64518 111922 64574 111978
rect 64642 111922 64698 111978
rect 240970 100294 241026 100350
rect 241094 100294 241150 100350
rect 241218 100294 241274 100350
rect 241342 100294 241398 100350
rect 240970 100170 241026 100226
rect 241094 100170 241150 100226
rect 241218 100170 241274 100226
rect 241342 100170 241398 100226
rect 240970 100046 241026 100102
rect 241094 100046 241150 100102
rect 241218 100046 241274 100102
rect 241342 100046 241398 100102
rect 240970 99922 241026 99978
rect 241094 99922 241150 99978
rect 241218 99922 241274 99978
rect 241342 99922 241398 99978
rect 57250 94294 57306 94350
rect 57374 94294 57430 94350
rect 57498 94294 57554 94350
rect 57622 94294 57678 94350
rect 57250 94170 57306 94226
rect 57374 94170 57430 94226
rect 57498 94170 57554 94226
rect 57622 94170 57678 94226
rect 57250 94046 57306 94102
rect 57374 94046 57430 94102
rect 57498 94046 57554 94102
rect 57622 94046 57678 94102
rect 57250 93922 57306 93978
rect 57374 93922 57430 93978
rect 57498 93922 57554 93978
rect 57622 93922 57678 93978
rect 42970 82294 43026 82350
rect 43094 82294 43150 82350
rect 43218 82294 43274 82350
rect 43342 82294 43398 82350
rect 42970 82170 43026 82226
rect 43094 82170 43150 82226
rect 43218 82170 43274 82226
rect 43342 82170 43398 82226
rect 42970 82046 43026 82102
rect 43094 82046 43150 82102
rect 43218 82046 43274 82102
rect 43342 82046 43398 82102
rect 42970 81922 43026 81978
rect 43094 81922 43150 81978
rect 43218 81922 43274 81978
rect 43342 81922 43398 81978
rect 64518 94294 64574 94350
rect 64642 94294 64698 94350
rect 64518 94170 64574 94226
rect 64642 94170 64698 94226
rect 64518 94046 64574 94102
rect 64642 94046 64698 94102
rect 64518 93922 64574 93978
rect 64642 93922 64698 93978
rect 240970 82294 241026 82350
rect 241094 82294 241150 82350
rect 241218 82294 241274 82350
rect 241342 82294 241398 82350
rect 240970 82170 241026 82226
rect 241094 82170 241150 82226
rect 241218 82170 241274 82226
rect 241342 82170 241398 82226
rect 240970 82046 241026 82102
rect 241094 82046 241150 82102
rect 241218 82046 241274 82102
rect 241342 82046 241398 82102
rect 240970 81922 241026 81978
rect 241094 81922 241150 81978
rect 241218 81922 241274 81978
rect 241342 81922 241398 81978
rect 57250 76294 57306 76350
rect 57374 76294 57430 76350
rect 57498 76294 57554 76350
rect 57622 76294 57678 76350
rect 57250 76170 57306 76226
rect 57374 76170 57430 76226
rect 57498 76170 57554 76226
rect 57622 76170 57678 76226
rect 57250 76046 57306 76102
rect 57374 76046 57430 76102
rect 57498 76046 57554 76102
rect 57622 76046 57678 76102
rect 57250 75922 57306 75978
rect 57374 75922 57430 75978
rect 57498 75922 57554 75978
rect 57622 75922 57678 75978
rect 42970 64294 43026 64350
rect 43094 64294 43150 64350
rect 43218 64294 43274 64350
rect 43342 64294 43398 64350
rect 42970 64170 43026 64226
rect 43094 64170 43150 64226
rect 43218 64170 43274 64226
rect 43342 64170 43398 64226
rect 42970 64046 43026 64102
rect 43094 64046 43150 64102
rect 43218 64046 43274 64102
rect 43342 64046 43398 64102
rect 42970 63922 43026 63978
rect 43094 63922 43150 63978
rect 43218 63922 43274 63978
rect 43342 63922 43398 63978
rect 64518 76294 64574 76350
rect 64642 76294 64698 76350
rect 64518 76170 64574 76226
rect 64642 76170 64698 76226
rect 64518 76046 64574 76102
rect 64642 76046 64698 76102
rect 64518 75922 64574 75978
rect 64642 75922 64698 75978
rect 240970 64294 241026 64350
rect 241094 64294 241150 64350
rect 241218 64294 241274 64350
rect 241342 64294 241398 64350
rect 240970 64170 241026 64226
rect 241094 64170 241150 64226
rect 241218 64170 241274 64226
rect 241342 64170 241398 64226
rect 240970 64046 241026 64102
rect 241094 64046 241150 64102
rect 241218 64046 241274 64102
rect 241342 64046 241398 64102
rect 240970 63922 241026 63978
rect 241094 63922 241150 63978
rect 241218 63922 241274 63978
rect 241342 63922 241398 63978
rect 57250 58294 57306 58350
rect 57374 58294 57430 58350
rect 57498 58294 57554 58350
rect 57622 58294 57678 58350
rect 57250 58170 57306 58226
rect 57374 58170 57430 58226
rect 57498 58170 57554 58226
rect 57622 58170 57678 58226
rect 57250 58046 57306 58102
rect 57374 58046 57430 58102
rect 57498 58046 57554 58102
rect 57622 58046 57678 58102
rect 57250 57922 57306 57978
rect 57374 57922 57430 57978
rect 57498 57922 57554 57978
rect 57622 57922 57678 57978
rect 42970 46294 43026 46350
rect 43094 46294 43150 46350
rect 43218 46294 43274 46350
rect 43342 46294 43398 46350
rect 42970 46170 43026 46226
rect 43094 46170 43150 46226
rect 43218 46170 43274 46226
rect 43342 46170 43398 46226
rect 42970 46046 43026 46102
rect 43094 46046 43150 46102
rect 43218 46046 43274 46102
rect 43342 46046 43398 46102
rect 42970 45922 43026 45978
rect 43094 45922 43150 45978
rect 43218 45922 43274 45978
rect 43342 45922 43398 45978
rect 42970 28294 43026 28350
rect 43094 28294 43150 28350
rect 43218 28294 43274 28350
rect 43342 28294 43398 28350
rect 42970 28170 43026 28226
rect 43094 28170 43150 28226
rect 43218 28170 43274 28226
rect 43342 28170 43398 28226
rect 42970 28046 43026 28102
rect 43094 28046 43150 28102
rect 43218 28046 43274 28102
rect 43342 28046 43398 28102
rect 42970 27922 43026 27978
rect 43094 27922 43150 27978
rect 43218 27922 43274 27978
rect 43342 27922 43398 27978
rect 42970 10294 43026 10350
rect 43094 10294 43150 10350
rect 43218 10294 43274 10350
rect 43342 10294 43398 10350
rect 42970 10170 43026 10226
rect 43094 10170 43150 10226
rect 43218 10170 43274 10226
rect 43342 10170 43398 10226
rect 42970 10046 43026 10102
rect 43094 10046 43150 10102
rect 43218 10046 43274 10102
rect 43342 10046 43398 10102
rect 42970 9922 43026 9978
rect 43094 9922 43150 9978
rect 43218 9922 43274 9978
rect 43342 9922 43398 9978
rect 42970 -1176 43026 -1120
rect 43094 -1176 43150 -1120
rect 43218 -1176 43274 -1120
rect 43342 -1176 43398 -1120
rect 42970 -1300 43026 -1244
rect 43094 -1300 43150 -1244
rect 43218 -1300 43274 -1244
rect 43342 -1300 43398 -1244
rect 42970 -1424 43026 -1368
rect 43094 -1424 43150 -1368
rect 43218 -1424 43274 -1368
rect 43342 -1424 43398 -1368
rect 42970 -1548 43026 -1492
rect 43094 -1548 43150 -1492
rect 43218 -1548 43274 -1492
rect 43342 -1548 43398 -1492
rect 64518 58294 64574 58350
rect 64642 58294 64698 58350
rect 64518 58170 64574 58226
rect 64642 58170 64698 58226
rect 64518 58046 64574 58102
rect 64642 58046 64698 58102
rect 64518 57922 64574 57978
rect 64642 57922 64698 57978
rect 240970 46294 241026 46350
rect 241094 46294 241150 46350
rect 241218 46294 241274 46350
rect 241342 46294 241398 46350
rect 240970 46170 241026 46226
rect 241094 46170 241150 46226
rect 241218 46170 241274 46226
rect 241342 46170 241398 46226
rect 240970 46046 241026 46102
rect 241094 46046 241150 46102
rect 241218 46046 241274 46102
rect 241342 46046 241398 46102
rect 240970 45922 241026 45978
rect 241094 45922 241150 45978
rect 241218 45922 241274 45978
rect 241342 45922 241398 45978
rect 57250 40294 57306 40350
rect 57374 40294 57430 40350
rect 57498 40294 57554 40350
rect 57622 40294 57678 40350
rect 57250 40170 57306 40226
rect 57374 40170 57430 40226
rect 57498 40170 57554 40226
rect 57622 40170 57678 40226
rect 57250 40046 57306 40102
rect 57374 40046 57430 40102
rect 57498 40046 57554 40102
rect 57622 40046 57678 40102
rect 57250 39922 57306 39978
rect 57374 39922 57430 39978
rect 57498 39922 57554 39978
rect 57622 39922 57678 39978
rect 64518 40294 64574 40350
rect 64642 40294 64698 40350
rect 64518 40170 64574 40226
rect 64642 40170 64698 40226
rect 64518 40046 64574 40102
rect 64642 40046 64698 40102
rect 64518 39922 64574 39978
rect 64642 39922 64698 39978
rect 238476 34442 238532 34498
rect 153468 33182 153524 33238
rect 57250 22294 57306 22350
rect 57374 22294 57430 22350
rect 57498 22294 57554 22350
rect 57622 22294 57678 22350
rect 57250 22170 57306 22226
rect 57374 22170 57430 22226
rect 57498 22170 57554 22226
rect 57622 22170 57678 22226
rect 57250 22046 57306 22102
rect 57374 22046 57430 22102
rect 57498 22046 57554 22102
rect 57622 22046 57678 22102
rect 57250 21922 57306 21978
rect 57374 21922 57430 21978
rect 57498 21922 57554 21978
rect 57622 21922 57678 21978
rect 57250 4294 57306 4350
rect 57374 4294 57430 4350
rect 57498 4294 57554 4350
rect 57622 4294 57678 4350
rect 57250 4170 57306 4226
rect 57374 4170 57430 4226
rect 57498 4170 57554 4226
rect 57622 4170 57678 4226
rect 57250 4046 57306 4102
rect 57374 4046 57430 4102
rect 57498 4046 57554 4102
rect 57622 4046 57678 4102
rect 57250 3922 57306 3978
rect 57374 3922 57430 3978
rect 57498 3922 57554 3978
rect 57622 3922 57678 3978
rect 57250 -216 57306 -160
rect 57374 -216 57430 -160
rect 57498 -216 57554 -160
rect 57622 -216 57678 -160
rect 57250 -340 57306 -284
rect 57374 -340 57430 -284
rect 57498 -340 57554 -284
rect 57622 -340 57678 -284
rect 57250 -464 57306 -408
rect 57374 -464 57430 -408
rect 57498 -464 57554 -408
rect 57622 -464 57678 -408
rect 57250 -588 57306 -532
rect 57374 -588 57430 -532
rect 57498 -588 57554 -532
rect 57622 -588 57678 -532
rect 60970 28294 61026 28350
rect 61094 28294 61150 28350
rect 61218 28294 61274 28350
rect 61342 28294 61398 28350
rect 60970 28170 61026 28226
rect 61094 28170 61150 28226
rect 61218 28170 61274 28226
rect 61342 28170 61398 28226
rect 60970 28046 61026 28102
rect 61094 28046 61150 28102
rect 61218 28046 61274 28102
rect 61342 28046 61398 28102
rect 60970 27922 61026 27978
rect 61094 27922 61150 27978
rect 61218 27922 61274 27978
rect 61342 27922 61398 27978
rect 73836 20042 73892 20098
rect 75250 22294 75306 22350
rect 75374 22294 75430 22350
rect 75498 22294 75554 22350
rect 75622 22294 75678 22350
rect 75250 22170 75306 22226
rect 75374 22170 75430 22226
rect 75498 22170 75554 22226
rect 75622 22170 75678 22226
rect 75250 22046 75306 22102
rect 75374 22046 75430 22102
rect 75498 22046 75554 22102
rect 75622 22046 75678 22102
rect 75250 21922 75306 21978
rect 75374 21922 75430 21978
rect 75498 21922 75554 21978
rect 75622 21922 75678 21978
rect 60970 10294 61026 10350
rect 61094 10294 61150 10350
rect 61218 10294 61274 10350
rect 61342 10294 61398 10350
rect 60970 10170 61026 10226
rect 61094 10170 61150 10226
rect 61218 10170 61274 10226
rect 61342 10170 61398 10226
rect 60970 10046 61026 10102
rect 61094 10046 61150 10102
rect 61218 10046 61274 10102
rect 61342 10046 61398 10102
rect 60970 9922 61026 9978
rect 61094 9922 61150 9978
rect 61218 9922 61274 9978
rect 61342 9922 61398 9978
rect 60970 -1176 61026 -1120
rect 61094 -1176 61150 -1120
rect 61218 -1176 61274 -1120
rect 61342 -1176 61398 -1120
rect 60970 -1300 61026 -1244
rect 61094 -1300 61150 -1244
rect 61218 -1300 61274 -1244
rect 61342 -1300 61398 -1244
rect 60970 -1424 61026 -1368
rect 61094 -1424 61150 -1368
rect 61218 -1424 61274 -1368
rect 61342 -1424 61398 -1368
rect 60970 -1548 61026 -1492
rect 61094 -1548 61150 -1492
rect 61218 -1548 61274 -1492
rect 61342 -1548 61398 -1492
rect 75250 4294 75306 4350
rect 75374 4294 75430 4350
rect 75498 4294 75554 4350
rect 75622 4294 75678 4350
rect 75250 4170 75306 4226
rect 75374 4170 75430 4226
rect 75498 4170 75554 4226
rect 75622 4170 75678 4226
rect 75250 4046 75306 4102
rect 75374 4046 75430 4102
rect 75498 4046 75554 4102
rect 75622 4046 75678 4102
rect 75250 3922 75306 3978
rect 75374 3922 75430 3978
rect 75498 3922 75554 3978
rect 75622 3922 75678 3978
rect 75250 -216 75306 -160
rect 75374 -216 75430 -160
rect 75498 -216 75554 -160
rect 75622 -216 75678 -160
rect 75250 -340 75306 -284
rect 75374 -340 75430 -284
rect 75498 -340 75554 -284
rect 75622 -340 75678 -284
rect 75250 -464 75306 -408
rect 75374 -464 75430 -408
rect 75498 -464 75554 -408
rect 75622 -464 75678 -408
rect 75250 -588 75306 -532
rect 75374 -588 75430 -532
rect 75498 -588 75554 -532
rect 75622 -588 75678 -532
rect 78970 28294 79026 28350
rect 79094 28294 79150 28350
rect 79218 28294 79274 28350
rect 79342 28294 79398 28350
rect 78970 28170 79026 28226
rect 79094 28170 79150 28226
rect 79218 28170 79274 28226
rect 79342 28170 79398 28226
rect 78970 28046 79026 28102
rect 79094 28046 79150 28102
rect 79218 28046 79274 28102
rect 79342 28046 79398 28102
rect 78970 27922 79026 27978
rect 79094 27922 79150 27978
rect 79218 27922 79274 27978
rect 79342 27922 79398 27978
rect 78970 10294 79026 10350
rect 79094 10294 79150 10350
rect 79218 10294 79274 10350
rect 79342 10294 79398 10350
rect 78970 10170 79026 10226
rect 79094 10170 79150 10226
rect 79218 10170 79274 10226
rect 79342 10170 79398 10226
rect 78970 10046 79026 10102
rect 79094 10046 79150 10102
rect 79218 10046 79274 10102
rect 79342 10046 79398 10102
rect 78970 9922 79026 9978
rect 79094 9922 79150 9978
rect 79218 9922 79274 9978
rect 79342 9922 79398 9978
rect 93250 22294 93306 22350
rect 93374 22294 93430 22350
rect 93498 22294 93554 22350
rect 93622 22294 93678 22350
rect 93250 22170 93306 22226
rect 93374 22170 93430 22226
rect 93498 22170 93554 22226
rect 93622 22170 93678 22226
rect 93250 22046 93306 22102
rect 93374 22046 93430 22102
rect 93498 22046 93554 22102
rect 93622 22046 93678 22102
rect 93250 21922 93306 21978
rect 93374 21922 93430 21978
rect 93498 21922 93554 21978
rect 93622 21922 93678 21978
rect 78970 -1176 79026 -1120
rect 79094 -1176 79150 -1120
rect 79218 -1176 79274 -1120
rect 79342 -1176 79398 -1120
rect 78970 -1300 79026 -1244
rect 79094 -1300 79150 -1244
rect 79218 -1300 79274 -1244
rect 79342 -1300 79398 -1244
rect 78970 -1424 79026 -1368
rect 79094 -1424 79150 -1368
rect 79218 -1424 79274 -1368
rect 79342 -1424 79398 -1368
rect 78970 -1548 79026 -1492
rect 79094 -1548 79150 -1492
rect 79218 -1548 79274 -1492
rect 79342 -1548 79398 -1492
rect 93250 4294 93306 4350
rect 93374 4294 93430 4350
rect 93498 4294 93554 4350
rect 93622 4294 93678 4350
rect 93250 4170 93306 4226
rect 93374 4170 93430 4226
rect 93498 4170 93554 4226
rect 93622 4170 93678 4226
rect 93250 4046 93306 4102
rect 93374 4046 93430 4102
rect 93498 4046 93554 4102
rect 93622 4046 93678 4102
rect 93250 3922 93306 3978
rect 93374 3922 93430 3978
rect 93498 3922 93554 3978
rect 93622 3922 93678 3978
rect 93250 -216 93306 -160
rect 93374 -216 93430 -160
rect 93498 -216 93554 -160
rect 93622 -216 93678 -160
rect 93250 -340 93306 -284
rect 93374 -340 93430 -284
rect 93498 -340 93554 -284
rect 93622 -340 93678 -284
rect 93250 -464 93306 -408
rect 93374 -464 93430 -408
rect 93498 -464 93554 -408
rect 93622 -464 93678 -408
rect 93250 -588 93306 -532
rect 93374 -588 93430 -532
rect 93498 -588 93554 -532
rect 93622 -588 93678 -532
rect 140812 31742 140868 31798
rect 139132 31562 139188 31618
rect 96970 28294 97026 28350
rect 97094 28294 97150 28350
rect 97218 28294 97274 28350
rect 97342 28294 97398 28350
rect 96970 28170 97026 28226
rect 97094 28170 97150 28226
rect 97218 28170 97274 28226
rect 97342 28170 97398 28226
rect 96970 28046 97026 28102
rect 97094 28046 97150 28102
rect 97218 28046 97274 28102
rect 97342 28046 97398 28102
rect 96970 27922 97026 27978
rect 97094 27922 97150 27978
rect 97218 27922 97274 27978
rect 97342 27922 97398 27978
rect 96970 10294 97026 10350
rect 97094 10294 97150 10350
rect 97218 10294 97274 10350
rect 97342 10294 97398 10350
rect 96970 10170 97026 10226
rect 97094 10170 97150 10226
rect 97218 10170 97274 10226
rect 97342 10170 97398 10226
rect 96970 10046 97026 10102
rect 97094 10046 97150 10102
rect 97218 10046 97274 10102
rect 97342 10046 97398 10102
rect 96970 9922 97026 9978
rect 97094 9922 97150 9978
rect 97218 9922 97274 9978
rect 97342 9922 97398 9978
rect 110460 26882 110516 26938
rect 112252 27602 112308 27658
rect 114970 28294 115026 28350
rect 115094 28294 115150 28350
rect 115218 28294 115274 28350
rect 115342 28294 115398 28350
rect 114970 28170 115026 28226
rect 115094 28170 115150 28226
rect 115218 28170 115274 28226
rect 115342 28170 115398 28226
rect 114970 28046 115026 28102
rect 115094 28046 115150 28102
rect 115218 28046 115274 28102
rect 115342 28046 115398 28102
rect 114970 27922 115026 27978
rect 115094 27922 115150 27978
rect 115218 27922 115274 27978
rect 115342 27922 115398 27978
rect 111250 22294 111306 22350
rect 111374 22294 111430 22350
rect 111498 22294 111554 22350
rect 111622 22294 111678 22350
rect 111250 22170 111306 22226
rect 111374 22170 111430 22226
rect 111498 22170 111554 22226
rect 111622 22170 111678 22226
rect 111250 22046 111306 22102
rect 111374 22046 111430 22102
rect 111498 22046 111554 22102
rect 111622 22046 111678 22102
rect 111250 21922 111306 21978
rect 111374 21922 111430 21978
rect 111498 21922 111554 21978
rect 111622 21922 111678 21978
rect 96970 -1176 97026 -1120
rect 97094 -1176 97150 -1120
rect 97218 -1176 97274 -1120
rect 97342 -1176 97398 -1120
rect 96970 -1300 97026 -1244
rect 97094 -1300 97150 -1244
rect 97218 -1300 97274 -1244
rect 97342 -1300 97398 -1244
rect 96970 -1424 97026 -1368
rect 97094 -1424 97150 -1368
rect 97218 -1424 97274 -1368
rect 97342 -1424 97398 -1368
rect 96970 -1548 97026 -1492
rect 97094 -1548 97150 -1492
rect 97218 -1548 97274 -1492
rect 97342 -1548 97398 -1492
rect 111250 4294 111306 4350
rect 111374 4294 111430 4350
rect 111498 4294 111554 4350
rect 111622 4294 111678 4350
rect 111250 4170 111306 4226
rect 111374 4170 111430 4226
rect 111498 4170 111554 4226
rect 111622 4170 111678 4226
rect 111250 4046 111306 4102
rect 111374 4046 111430 4102
rect 111498 4046 111554 4102
rect 111622 4046 111678 4102
rect 111250 3922 111306 3978
rect 111374 3922 111430 3978
rect 111498 3922 111554 3978
rect 111622 3922 111678 3978
rect 111250 -216 111306 -160
rect 111374 -216 111430 -160
rect 111498 -216 111554 -160
rect 111622 -216 111678 -160
rect 111250 -340 111306 -284
rect 111374 -340 111430 -284
rect 111498 -340 111554 -284
rect 111622 -340 111678 -284
rect 111250 -464 111306 -408
rect 111374 -464 111430 -408
rect 111498 -464 111554 -408
rect 111622 -464 111678 -408
rect 111250 -588 111306 -532
rect 111374 -588 111430 -532
rect 111498 -588 111554 -532
rect 111622 -588 111678 -532
rect 114970 10294 115026 10350
rect 115094 10294 115150 10350
rect 115218 10294 115274 10350
rect 115342 10294 115398 10350
rect 114970 10170 115026 10226
rect 115094 10170 115150 10226
rect 115218 10170 115274 10226
rect 115342 10170 115398 10226
rect 114970 10046 115026 10102
rect 115094 10046 115150 10102
rect 115218 10046 115274 10102
rect 115342 10046 115398 10102
rect 114970 9922 115026 9978
rect 115094 9922 115150 9978
rect 115218 9922 115274 9978
rect 115342 9922 115398 9978
rect 114970 -1176 115026 -1120
rect 115094 -1176 115150 -1120
rect 115218 -1176 115274 -1120
rect 115342 -1176 115398 -1120
rect 114970 -1300 115026 -1244
rect 115094 -1300 115150 -1244
rect 115218 -1300 115274 -1244
rect 115342 -1300 115398 -1244
rect 114970 -1424 115026 -1368
rect 115094 -1424 115150 -1368
rect 115218 -1424 115274 -1368
rect 115342 -1424 115398 -1368
rect 114970 -1548 115026 -1492
rect 115094 -1548 115150 -1492
rect 115218 -1548 115274 -1492
rect 115342 -1548 115398 -1492
rect 129250 22294 129306 22350
rect 129374 22294 129430 22350
rect 129498 22294 129554 22350
rect 129622 22294 129678 22350
rect 129250 22170 129306 22226
rect 129374 22170 129430 22226
rect 129498 22170 129554 22226
rect 129622 22170 129678 22226
rect 129250 22046 129306 22102
rect 129374 22046 129430 22102
rect 129498 22046 129554 22102
rect 129622 22046 129678 22102
rect 129250 21922 129306 21978
rect 129374 21922 129430 21978
rect 129498 21922 129554 21978
rect 129622 21922 129678 21978
rect 129250 4294 129306 4350
rect 129374 4294 129430 4350
rect 129498 4294 129554 4350
rect 129622 4294 129678 4350
rect 129250 4170 129306 4226
rect 129374 4170 129430 4226
rect 129498 4170 129554 4226
rect 129622 4170 129678 4226
rect 129250 4046 129306 4102
rect 129374 4046 129430 4102
rect 129498 4046 129554 4102
rect 129622 4046 129678 4102
rect 129250 3922 129306 3978
rect 129374 3922 129430 3978
rect 129498 3922 129554 3978
rect 129622 3922 129678 3978
rect 129250 -216 129306 -160
rect 129374 -216 129430 -160
rect 129498 -216 129554 -160
rect 129622 -216 129678 -160
rect 129250 -340 129306 -284
rect 129374 -340 129430 -284
rect 129498 -340 129554 -284
rect 129622 -340 129678 -284
rect 129250 -464 129306 -408
rect 129374 -464 129430 -408
rect 129498 -464 129554 -408
rect 129622 -464 129678 -408
rect 129250 -588 129306 -532
rect 129374 -588 129430 -532
rect 129498 -588 129554 -532
rect 129622 -588 129678 -532
rect 132970 28294 133026 28350
rect 133094 28294 133150 28350
rect 133218 28294 133274 28350
rect 133342 28294 133398 28350
rect 132970 28170 133026 28226
rect 133094 28170 133150 28226
rect 133218 28170 133274 28226
rect 133342 28170 133398 28226
rect 132970 28046 133026 28102
rect 133094 28046 133150 28102
rect 133218 28046 133274 28102
rect 133342 28046 133398 28102
rect 132970 27922 133026 27978
rect 133094 27922 133150 27978
rect 133218 27922 133274 27978
rect 133342 27922 133398 27978
rect 132970 10294 133026 10350
rect 133094 10294 133150 10350
rect 133218 10294 133274 10350
rect 133342 10294 133398 10350
rect 132970 10170 133026 10226
rect 133094 10170 133150 10226
rect 133218 10170 133274 10226
rect 133342 10170 133398 10226
rect 132970 10046 133026 10102
rect 133094 10046 133150 10102
rect 133218 10046 133274 10102
rect 133342 10046 133398 10102
rect 132970 9922 133026 9978
rect 133094 9922 133150 9978
rect 133218 9922 133274 9978
rect 133342 9922 133398 9978
rect 140924 31382 140980 31438
rect 142716 31202 142772 31258
rect 149884 31022 149940 31078
rect 147868 29764 147924 29818
rect 147868 29762 147924 29764
rect 147250 22294 147306 22350
rect 147374 22294 147430 22350
rect 147498 22294 147554 22350
rect 147622 22294 147678 22350
rect 147250 22170 147306 22226
rect 147374 22170 147430 22226
rect 147498 22170 147554 22226
rect 147622 22170 147678 22226
rect 147250 22046 147306 22102
rect 147374 22046 147430 22102
rect 147498 22046 147554 22102
rect 147622 22046 147678 22102
rect 147250 21922 147306 21978
rect 147374 21922 147430 21978
rect 147498 21922 147554 21978
rect 147622 21922 147678 21978
rect 132970 -1176 133026 -1120
rect 133094 -1176 133150 -1120
rect 133218 -1176 133274 -1120
rect 133342 -1176 133398 -1120
rect 132970 -1300 133026 -1244
rect 133094 -1300 133150 -1244
rect 133218 -1300 133274 -1244
rect 133342 -1300 133398 -1244
rect 132970 -1424 133026 -1368
rect 133094 -1424 133150 -1368
rect 133218 -1424 133274 -1368
rect 133342 -1424 133398 -1368
rect 132970 -1548 133026 -1492
rect 133094 -1548 133150 -1492
rect 133218 -1548 133274 -1492
rect 133342 -1548 133398 -1492
rect 158844 33002 158900 33058
rect 160636 32822 160692 32878
rect 162428 32642 162484 32698
rect 157052 30122 157108 30178
rect 150970 28294 151026 28350
rect 151094 28294 151150 28350
rect 151218 28294 151274 28350
rect 151342 28294 151398 28350
rect 150970 28170 151026 28226
rect 151094 28170 151150 28226
rect 151218 28170 151274 28226
rect 151342 28170 151398 28226
rect 150970 28046 151026 28102
rect 151094 28046 151150 28102
rect 151218 28046 151274 28102
rect 151342 28046 151398 28102
rect 150970 27922 151026 27978
rect 151094 27922 151150 27978
rect 151218 27922 151274 27978
rect 151342 27922 151398 27978
rect 147250 4294 147306 4350
rect 147374 4294 147430 4350
rect 147498 4294 147554 4350
rect 147622 4294 147678 4350
rect 147250 4170 147306 4226
rect 147374 4170 147430 4226
rect 147498 4170 147554 4226
rect 147622 4170 147678 4226
rect 147250 4046 147306 4102
rect 147374 4046 147430 4102
rect 147498 4046 147554 4102
rect 147622 4046 147678 4102
rect 147250 3922 147306 3978
rect 147374 3922 147430 3978
rect 147498 3922 147554 3978
rect 147622 3922 147678 3978
rect 147250 -216 147306 -160
rect 147374 -216 147430 -160
rect 147498 -216 147554 -160
rect 147622 -216 147678 -160
rect 147250 -340 147306 -284
rect 147374 -340 147430 -284
rect 147498 -340 147554 -284
rect 147622 -340 147678 -284
rect 147250 -464 147306 -408
rect 147374 -464 147430 -408
rect 147498 -464 147554 -408
rect 147622 -464 147678 -408
rect 147250 -588 147306 -532
rect 147374 -588 147430 -532
rect 147498 -588 147554 -532
rect 147622 -588 147678 -532
rect 155260 29942 155316 29998
rect 165250 22294 165306 22350
rect 165374 22294 165430 22350
rect 165498 22294 165554 22350
rect 165622 22294 165678 22350
rect 165250 22170 165306 22226
rect 165374 22170 165430 22226
rect 165498 22170 165554 22226
rect 165622 22170 165678 22226
rect 165250 22046 165306 22102
rect 165374 22046 165430 22102
rect 165498 22046 165554 22102
rect 165622 22046 165678 22102
rect 165250 21922 165306 21978
rect 165374 21922 165430 21978
rect 165498 21922 165554 21978
rect 165622 21922 165678 21978
rect 150970 10294 151026 10350
rect 151094 10294 151150 10350
rect 151218 10294 151274 10350
rect 151342 10294 151398 10350
rect 150970 10170 151026 10226
rect 151094 10170 151150 10226
rect 151218 10170 151274 10226
rect 151342 10170 151398 10226
rect 150970 10046 151026 10102
rect 151094 10046 151150 10102
rect 151218 10046 151274 10102
rect 151342 10046 151398 10102
rect 150970 9922 151026 9978
rect 151094 9922 151150 9978
rect 151218 9922 151274 9978
rect 151342 9922 151398 9978
rect 150970 -1176 151026 -1120
rect 151094 -1176 151150 -1120
rect 151218 -1176 151274 -1120
rect 151342 -1176 151398 -1120
rect 150970 -1300 151026 -1244
rect 151094 -1300 151150 -1244
rect 151218 -1300 151274 -1244
rect 151342 -1300 151398 -1244
rect 150970 -1424 151026 -1368
rect 151094 -1424 151150 -1368
rect 151218 -1424 151274 -1368
rect 151342 -1424 151398 -1368
rect 150970 -1548 151026 -1492
rect 151094 -1548 151150 -1492
rect 151218 -1548 151274 -1492
rect 151342 -1548 151398 -1492
rect 165250 4294 165306 4350
rect 165374 4294 165430 4350
rect 165498 4294 165554 4350
rect 165622 4294 165678 4350
rect 165250 4170 165306 4226
rect 165374 4170 165430 4226
rect 165498 4170 165554 4226
rect 165622 4170 165678 4226
rect 165250 4046 165306 4102
rect 165374 4046 165430 4102
rect 165498 4046 165554 4102
rect 165622 4046 165678 4102
rect 165250 3922 165306 3978
rect 165374 3922 165430 3978
rect 165498 3922 165554 3978
rect 165622 3922 165678 3978
rect 165250 -216 165306 -160
rect 165374 -216 165430 -160
rect 165498 -216 165554 -160
rect 165622 -216 165678 -160
rect 165250 -340 165306 -284
rect 165374 -340 165430 -284
rect 165498 -340 165554 -284
rect 165622 -340 165678 -284
rect 165250 -464 165306 -408
rect 165374 -464 165430 -408
rect 165498 -464 165554 -408
rect 165622 -464 165678 -408
rect 165250 -588 165306 -532
rect 165374 -588 165430 -532
rect 165498 -588 165554 -532
rect 165622 -588 165678 -532
rect 168970 28294 169026 28350
rect 169094 28294 169150 28350
rect 169218 28294 169274 28350
rect 169342 28294 169398 28350
rect 168970 28170 169026 28226
rect 169094 28170 169150 28226
rect 169218 28170 169274 28226
rect 169342 28170 169398 28226
rect 168970 28046 169026 28102
rect 169094 28046 169150 28102
rect 169218 28046 169274 28102
rect 169342 28046 169398 28102
rect 168970 27922 169026 27978
rect 169094 27922 169150 27978
rect 169218 27922 169274 27978
rect 169342 27922 169398 27978
rect 168970 10294 169026 10350
rect 169094 10294 169150 10350
rect 169218 10294 169274 10350
rect 169342 10294 169398 10350
rect 168970 10170 169026 10226
rect 169094 10170 169150 10226
rect 169218 10170 169274 10226
rect 169342 10170 169398 10226
rect 168970 10046 169026 10102
rect 169094 10046 169150 10102
rect 169218 10046 169274 10102
rect 169342 10046 169398 10102
rect 168970 9922 169026 9978
rect 169094 9922 169150 9978
rect 169218 9922 169274 9978
rect 169342 9922 169398 9978
rect 168970 -1176 169026 -1120
rect 169094 -1176 169150 -1120
rect 169218 -1176 169274 -1120
rect 169342 -1176 169398 -1120
rect 168970 -1300 169026 -1244
rect 169094 -1300 169150 -1244
rect 169218 -1300 169274 -1244
rect 169342 -1300 169398 -1244
rect 168970 -1424 169026 -1368
rect 169094 -1424 169150 -1368
rect 169218 -1424 169274 -1368
rect 169342 -1424 169398 -1368
rect 168970 -1548 169026 -1492
rect 169094 -1548 169150 -1492
rect 169218 -1548 169274 -1492
rect 169342 -1548 169398 -1492
rect 186508 29402 186564 29458
rect 186970 28294 187026 28350
rect 187094 28294 187150 28350
rect 187218 28294 187274 28350
rect 187342 28294 187398 28350
rect 186970 28170 187026 28226
rect 187094 28170 187150 28226
rect 187218 28170 187274 28226
rect 187342 28170 187398 28226
rect 186970 28046 187026 28102
rect 187094 28046 187150 28102
rect 187218 28046 187274 28102
rect 187342 28046 187398 28102
rect 186970 27922 187026 27978
rect 187094 27922 187150 27978
rect 187218 27922 187274 27978
rect 187342 27922 187398 27978
rect 183250 22294 183306 22350
rect 183374 22294 183430 22350
rect 183498 22294 183554 22350
rect 183622 22294 183678 22350
rect 183250 22170 183306 22226
rect 183374 22170 183430 22226
rect 183498 22170 183554 22226
rect 183622 22170 183678 22226
rect 183250 22046 183306 22102
rect 183374 22046 183430 22102
rect 183498 22046 183554 22102
rect 183622 22046 183678 22102
rect 183250 21922 183306 21978
rect 183374 21922 183430 21978
rect 183498 21922 183554 21978
rect 183622 21922 183678 21978
rect 183250 4294 183306 4350
rect 183374 4294 183430 4350
rect 183498 4294 183554 4350
rect 183622 4294 183678 4350
rect 183250 4170 183306 4226
rect 183374 4170 183430 4226
rect 183498 4170 183554 4226
rect 183622 4170 183678 4226
rect 183250 4046 183306 4102
rect 183374 4046 183430 4102
rect 183498 4046 183554 4102
rect 183622 4046 183678 4102
rect 183250 3922 183306 3978
rect 183374 3922 183430 3978
rect 183498 3922 183554 3978
rect 183622 3922 183678 3978
rect 183250 -216 183306 -160
rect 183374 -216 183430 -160
rect 183498 -216 183554 -160
rect 183622 -216 183678 -160
rect 183250 -340 183306 -284
rect 183374 -340 183430 -284
rect 183498 -340 183554 -284
rect 183622 -340 183678 -284
rect 183250 -464 183306 -408
rect 183374 -464 183430 -408
rect 183498 -464 183554 -408
rect 183622 -464 183678 -408
rect 183250 -588 183306 -532
rect 183374 -588 183430 -532
rect 183498 -588 183554 -532
rect 183622 -588 183678 -532
rect 186970 10294 187026 10350
rect 187094 10294 187150 10350
rect 187218 10294 187274 10350
rect 187342 10294 187398 10350
rect 186970 10170 187026 10226
rect 187094 10170 187150 10226
rect 187218 10170 187274 10226
rect 187342 10170 187398 10226
rect 186970 10046 187026 10102
rect 187094 10046 187150 10102
rect 187218 10046 187274 10102
rect 187342 10046 187398 10102
rect 186970 9922 187026 9978
rect 187094 9922 187150 9978
rect 187218 9922 187274 9978
rect 187342 9922 187398 9978
rect 186970 -1176 187026 -1120
rect 187094 -1176 187150 -1120
rect 187218 -1176 187274 -1120
rect 187342 -1176 187398 -1120
rect 186970 -1300 187026 -1244
rect 187094 -1300 187150 -1244
rect 187218 -1300 187274 -1244
rect 187342 -1300 187398 -1244
rect 186970 -1424 187026 -1368
rect 187094 -1424 187150 -1368
rect 187218 -1424 187274 -1368
rect 187342 -1424 187398 -1368
rect 186970 -1548 187026 -1492
rect 187094 -1548 187150 -1492
rect 187218 -1548 187274 -1492
rect 187342 -1548 187398 -1492
rect 204970 28294 205026 28350
rect 205094 28294 205150 28350
rect 205218 28294 205274 28350
rect 205342 28294 205398 28350
rect 204970 28170 205026 28226
rect 205094 28170 205150 28226
rect 205218 28170 205274 28226
rect 205342 28170 205398 28226
rect 204970 28046 205026 28102
rect 205094 28046 205150 28102
rect 205218 28046 205274 28102
rect 205342 28046 205398 28102
rect 204970 27922 205026 27978
rect 205094 27922 205150 27978
rect 205218 27922 205274 27978
rect 205342 27922 205398 27978
rect 203308 27636 203364 27658
rect 203308 27602 203364 27636
rect 201250 22294 201306 22350
rect 201374 22294 201430 22350
rect 201498 22294 201554 22350
rect 201622 22294 201678 22350
rect 201250 22170 201306 22226
rect 201374 22170 201430 22226
rect 201498 22170 201554 22226
rect 201622 22170 201678 22226
rect 201250 22046 201306 22102
rect 201374 22046 201430 22102
rect 201498 22046 201554 22102
rect 201622 22046 201678 22102
rect 201250 21922 201306 21978
rect 201374 21922 201430 21978
rect 201498 21922 201554 21978
rect 201622 21922 201678 21978
rect 201250 4294 201306 4350
rect 201374 4294 201430 4350
rect 201498 4294 201554 4350
rect 201622 4294 201678 4350
rect 201250 4170 201306 4226
rect 201374 4170 201430 4226
rect 201498 4170 201554 4226
rect 201622 4170 201678 4226
rect 201250 4046 201306 4102
rect 201374 4046 201430 4102
rect 201498 4046 201554 4102
rect 201622 4046 201678 4102
rect 201250 3922 201306 3978
rect 201374 3922 201430 3978
rect 201498 3922 201554 3978
rect 201622 3922 201678 3978
rect 201250 -216 201306 -160
rect 201374 -216 201430 -160
rect 201498 -216 201554 -160
rect 201622 -216 201678 -160
rect 201250 -340 201306 -284
rect 201374 -340 201430 -284
rect 201498 -340 201554 -284
rect 201622 -340 201678 -284
rect 201250 -464 201306 -408
rect 201374 -464 201430 -408
rect 201498 -464 201554 -408
rect 201622 -464 201678 -408
rect 201250 -588 201306 -532
rect 201374 -588 201430 -532
rect 201498 -588 201554 -532
rect 201622 -588 201678 -532
rect 215852 27602 215908 27658
rect 209356 26882 209412 26938
rect 218428 27422 218484 27478
rect 221564 29596 221620 29638
rect 221564 29582 221620 29596
rect 219884 27422 219940 27478
rect 219250 22294 219306 22350
rect 219374 22294 219430 22350
rect 219498 22294 219554 22350
rect 219622 22294 219678 22350
rect 219250 22170 219306 22226
rect 219374 22170 219430 22226
rect 219498 22170 219554 22226
rect 219622 22170 219678 22226
rect 219250 22046 219306 22102
rect 219374 22046 219430 22102
rect 219498 22046 219554 22102
rect 219622 22046 219678 22102
rect 219250 21922 219306 21978
rect 219374 21922 219430 21978
rect 219498 21922 219554 21978
rect 219622 21922 219678 21978
rect 204970 10294 205026 10350
rect 205094 10294 205150 10350
rect 205218 10294 205274 10350
rect 205342 10294 205398 10350
rect 204970 10170 205026 10226
rect 205094 10170 205150 10226
rect 205218 10170 205274 10226
rect 205342 10170 205398 10226
rect 204970 10046 205026 10102
rect 205094 10046 205150 10102
rect 205218 10046 205274 10102
rect 205342 10046 205398 10102
rect 204970 9922 205026 9978
rect 205094 9922 205150 9978
rect 205218 9922 205274 9978
rect 205342 9922 205398 9978
rect 204970 -1176 205026 -1120
rect 205094 -1176 205150 -1120
rect 205218 -1176 205274 -1120
rect 205342 -1176 205398 -1120
rect 204970 -1300 205026 -1244
rect 205094 -1300 205150 -1244
rect 205218 -1300 205274 -1244
rect 205342 -1300 205398 -1244
rect 204970 -1424 205026 -1368
rect 205094 -1424 205150 -1368
rect 205218 -1424 205274 -1368
rect 205342 -1424 205398 -1368
rect 204970 -1548 205026 -1492
rect 205094 -1548 205150 -1492
rect 205218 -1548 205274 -1492
rect 205342 -1548 205398 -1492
rect 222970 28294 223026 28350
rect 223094 28294 223150 28350
rect 223218 28294 223274 28350
rect 223342 28294 223398 28350
rect 222970 28170 223026 28226
rect 223094 28170 223150 28226
rect 223218 28170 223274 28226
rect 223342 28170 223398 28226
rect 222970 28046 223026 28102
rect 223094 28046 223150 28102
rect 223218 28046 223274 28102
rect 223342 28046 223398 28102
rect 222970 27922 223026 27978
rect 223094 27922 223150 27978
rect 223218 27922 223274 27978
rect 223342 27922 223398 27978
rect 219250 4294 219306 4350
rect 219374 4294 219430 4350
rect 219498 4294 219554 4350
rect 219622 4294 219678 4350
rect 219250 4170 219306 4226
rect 219374 4170 219430 4226
rect 219498 4170 219554 4226
rect 219622 4170 219678 4226
rect 219250 4046 219306 4102
rect 219374 4046 219430 4102
rect 219498 4046 219554 4102
rect 219622 4046 219678 4102
rect 219250 3922 219306 3978
rect 219374 3922 219430 3978
rect 219498 3922 219554 3978
rect 219622 3922 219678 3978
rect 219250 -216 219306 -160
rect 219374 -216 219430 -160
rect 219498 -216 219554 -160
rect 219622 -216 219678 -160
rect 219250 -340 219306 -284
rect 219374 -340 219430 -284
rect 219498 -340 219554 -284
rect 219622 -340 219678 -284
rect 219250 -464 219306 -408
rect 219374 -464 219430 -408
rect 219498 -464 219554 -408
rect 219622 -464 219678 -408
rect 219250 -588 219306 -532
rect 219374 -588 219430 -532
rect 219498 -588 219554 -532
rect 219622 -588 219678 -532
rect 222970 10294 223026 10350
rect 223094 10294 223150 10350
rect 223218 10294 223274 10350
rect 223342 10294 223398 10350
rect 222970 10170 223026 10226
rect 223094 10170 223150 10226
rect 223218 10170 223274 10226
rect 223342 10170 223398 10226
rect 222970 10046 223026 10102
rect 223094 10046 223150 10102
rect 223218 10046 223274 10102
rect 223342 10046 223398 10102
rect 222970 9922 223026 9978
rect 223094 9922 223150 9978
rect 223218 9922 223274 9978
rect 223342 9922 223398 9978
rect 222970 -1176 223026 -1120
rect 223094 -1176 223150 -1120
rect 223218 -1176 223274 -1120
rect 223342 -1176 223398 -1120
rect 222970 -1300 223026 -1244
rect 223094 -1300 223150 -1244
rect 223218 -1300 223274 -1244
rect 223342 -1300 223398 -1244
rect 222970 -1424 223026 -1368
rect 223094 -1424 223150 -1368
rect 223218 -1424 223274 -1368
rect 223342 -1424 223398 -1368
rect 222970 -1548 223026 -1492
rect 223094 -1548 223150 -1492
rect 223218 -1548 223274 -1492
rect 223342 -1548 223398 -1492
rect 255250 202294 255306 202350
rect 255374 202294 255430 202350
rect 255498 202294 255554 202350
rect 255622 202294 255678 202350
rect 255250 202170 255306 202226
rect 255374 202170 255430 202226
rect 255498 202170 255554 202226
rect 255622 202170 255678 202226
rect 255250 202046 255306 202102
rect 255374 202046 255430 202102
rect 255498 202046 255554 202102
rect 255622 202046 255678 202102
rect 255250 201922 255306 201978
rect 255374 201922 255430 201978
rect 255498 201922 255554 201978
rect 255622 201922 255678 201978
rect 258970 226294 259026 226350
rect 259094 226294 259150 226350
rect 259218 226294 259274 226350
rect 259342 226294 259398 226350
rect 258970 226170 259026 226226
rect 259094 226170 259150 226226
rect 259218 226170 259274 226226
rect 259342 226170 259398 226226
rect 258970 226046 259026 226102
rect 259094 226046 259150 226102
rect 259218 226046 259274 226102
rect 259342 226046 259398 226102
rect 258970 225922 259026 225978
rect 259094 225922 259150 225978
rect 259218 225922 259274 225978
rect 259342 225922 259398 225978
rect 273250 597156 273306 597212
rect 273374 597156 273430 597212
rect 273498 597156 273554 597212
rect 273622 597156 273678 597212
rect 273250 597032 273306 597088
rect 273374 597032 273430 597088
rect 273498 597032 273554 597088
rect 273622 597032 273678 597088
rect 273250 596908 273306 596964
rect 273374 596908 273430 596964
rect 273498 596908 273554 596964
rect 273622 596908 273678 596964
rect 273250 596784 273306 596840
rect 273374 596784 273430 596840
rect 273498 596784 273554 596840
rect 273622 596784 273678 596840
rect 273250 580294 273306 580350
rect 273374 580294 273430 580350
rect 273498 580294 273554 580350
rect 273622 580294 273678 580350
rect 273250 580170 273306 580226
rect 273374 580170 273430 580226
rect 273498 580170 273554 580226
rect 273622 580170 273678 580226
rect 273250 580046 273306 580102
rect 273374 580046 273430 580102
rect 273498 580046 273554 580102
rect 273622 580046 273678 580102
rect 273250 579922 273306 579978
rect 273374 579922 273430 579978
rect 273498 579922 273554 579978
rect 273622 579922 273678 579978
rect 273250 562294 273306 562350
rect 273374 562294 273430 562350
rect 273498 562294 273554 562350
rect 273622 562294 273678 562350
rect 273250 562170 273306 562226
rect 273374 562170 273430 562226
rect 273498 562170 273554 562226
rect 273622 562170 273678 562226
rect 273250 562046 273306 562102
rect 273374 562046 273430 562102
rect 273498 562046 273554 562102
rect 273622 562046 273678 562102
rect 273250 561922 273306 561978
rect 273374 561922 273430 561978
rect 273498 561922 273554 561978
rect 273622 561922 273678 561978
rect 273250 544294 273306 544350
rect 273374 544294 273430 544350
rect 273498 544294 273554 544350
rect 273622 544294 273678 544350
rect 273250 544170 273306 544226
rect 273374 544170 273430 544226
rect 273498 544170 273554 544226
rect 273622 544170 273678 544226
rect 273250 544046 273306 544102
rect 273374 544046 273430 544102
rect 273498 544046 273554 544102
rect 273622 544046 273678 544102
rect 273250 543922 273306 543978
rect 273374 543922 273430 543978
rect 273498 543922 273554 543978
rect 273622 543922 273678 543978
rect 273250 526294 273306 526350
rect 273374 526294 273430 526350
rect 273498 526294 273554 526350
rect 273622 526294 273678 526350
rect 273250 526170 273306 526226
rect 273374 526170 273430 526226
rect 273498 526170 273554 526226
rect 273622 526170 273678 526226
rect 273250 526046 273306 526102
rect 273374 526046 273430 526102
rect 273498 526046 273554 526102
rect 273622 526046 273678 526102
rect 273250 525922 273306 525978
rect 273374 525922 273430 525978
rect 273498 525922 273554 525978
rect 273622 525922 273678 525978
rect 273250 508294 273306 508350
rect 273374 508294 273430 508350
rect 273498 508294 273554 508350
rect 273622 508294 273678 508350
rect 273250 508170 273306 508226
rect 273374 508170 273430 508226
rect 273498 508170 273554 508226
rect 273622 508170 273678 508226
rect 273250 508046 273306 508102
rect 273374 508046 273430 508102
rect 273498 508046 273554 508102
rect 273622 508046 273678 508102
rect 273250 507922 273306 507978
rect 273374 507922 273430 507978
rect 273498 507922 273554 507978
rect 273622 507922 273678 507978
rect 273250 490294 273306 490350
rect 273374 490294 273430 490350
rect 273498 490294 273554 490350
rect 273622 490294 273678 490350
rect 273250 490170 273306 490226
rect 273374 490170 273430 490226
rect 273498 490170 273554 490226
rect 273622 490170 273678 490226
rect 273250 490046 273306 490102
rect 273374 490046 273430 490102
rect 273498 490046 273554 490102
rect 273622 490046 273678 490102
rect 273250 489922 273306 489978
rect 273374 489922 273430 489978
rect 273498 489922 273554 489978
rect 273622 489922 273678 489978
rect 273250 472294 273306 472350
rect 273374 472294 273430 472350
rect 273498 472294 273554 472350
rect 273622 472294 273678 472350
rect 273250 472170 273306 472226
rect 273374 472170 273430 472226
rect 273498 472170 273554 472226
rect 273622 472170 273678 472226
rect 273250 472046 273306 472102
rect 273374 472046 273430 472102
rect 273498 472046 273554 472102
rect 273622 472046 273678 472102
rect 273250 471922 273306 471978
rect 273374 471922 273430 471978
rect 273498 471922 273554 471978
rect 273622 471922 273678 471978
rect 273250 454294 273306 454350
rect 273374 454294 273430 454350
rect 273498 454294 273554 454350
rect 273622 454294 273678 454350
rect 273250 454170 273306 454226
rect 273374 454170 273430 454226
rect 273498 454170 273554 454226
rect 273622 454170 273678 454226
rect 273250 454046 273306 454102
rect 273374 454046 273430 454102
rect 273498 454046 273554 454102
rect 273622 454046 273678 454102
rect 273250 453922 273306 453978
rect 273374 453922 273430 453978
rect 273498 453922 273554 453978
rect 273622 453922 273678 453978
rect 273250 436294 273306 436350
rect 273374 436294 273430 436350
rect 273498 436294 273554 436350
rect 273622 436294 273678 436350
rect 273250 436170 273306 436226
rect 273374 436170 273430 436226
rect 273498 436170 273554 436226
rect 273622 436170 273678 436226
rect 273250 436046 273306 436102
rect 273374 436046 273430 436102
rect 273498 436046 273554 436102
rect 273622 436046 273678 436102
rect 273250 435922 273306 435978
rect 273374 435922 273430 435978
rect 273498 435922 273554 435978
rect 273622 435922 273678 435978
rect 273250 418294 273306 418350
rect 273374 418294 273430 418350
rect 273498 418294 273554 418350
rect 273622 418294 273678 418350
rect 273250 418170 273306 418226
rect 273374 418170 273430 418226
rect 273498 418170 273554 418226
rect 273622 418170 273678 418226
rect 273250 418046 273306 418102
rect 273374 418046 273430 418102
rect 273498 418046 273554 418102
rect 273622 418046 273678 418102
rect 273250 417922 273306 417978
rect 273374 417922 273430 417978
rect 273498 417922 273554 417978
rect 273622 417922 273678 417978
rect 273250 400294 273306 400350
rect 273374 400294 273430 400350
rect 273498 400294 273554 400350
rect 273622 400294 273678 400350
rect 273250 400170 273306 400226
rect 273374 400170 273430 400226
rect 273498 400170 273554 400226
rect 273622 400170 273678 400226
rect 273250 400046 273306 400102
rect 273374 400046 273430 400102
rect 273498 400046 273554 400102
rect 273622 400046 273678 400102
rect 273250 399922 273306 399978
rect 273374 399922 273430 399978
rect 273498 399922 273554 399978
rect 273622 399922 273678 399978
rect 273250 382294 273306 382350
rect 273374 382294 273430 382350
rect 273498 382294 273554 382350
rect 273622 382294 273678 382350
rect 273250 382170 273306 382226
rect 273374 382170 273430 382226
rect 273498 382170 273554 382226
rect 273622 382170 273678 382226
rect 273250 382046 273306 382102
rect 273374 382046 273430 382102
rect 273498 382046 273554 382102
rect 273622 382046 273678 382102
rect 273250 381922 273306 381978
rect 273374 381922 273430 381978
rect 273498 381922 273554 381978
rect 273622 381922 273678 381978
rect 273250 364294 273306 364350
rect 273374 364294 273430 364350
rect 273498 364294 273554 364350
rect 273622 364294 273678 364350
rect 273250 364170 273306 364226
rect 273374 364170 273430 364226
rect 273498 364170 273554 364226
rect 273622 364170 273678 364226
rect 273250 364046 273306 364102
rect 273374 364046 273430 364102
rect 273498 364046 273554 364102
rect 273622 364046 273678 364102
rect 273250 363922 273306 363978
rect 273374 363922 273430 363978
rect 273498 363922 273554 363978
rect 273622 363922 273678 363978
rect 273250 346294 273306 346350
rect 273374 346294 273430 346350
rect 273498 346294 273554 346350
rect 273622 346294 273678 346350
rect 273250 346170 273306 346226
rect 273374 346170 273430 346226
rect 273498 346170 273554 346226
rect 273622 346170 273678 346226
rect 273250 346046 273306 346102
rect 273374 346046 273430 346102
rect 273498 346046 273554 346102
rect 273622 346046 273678 346102
rect 273250 345922 273306 345978
rect 273374 345922 273430 345978
rect 273498 345922 273554 345978
rect 273622 345922 273678 345978
rect 273250 328294 273306 328350
rect 273374 328294 273430 328350
rect 273498 328294 273554 328350
rect 273622 328294 273678 328350
rect 273250 328170 273306 328226
rect 273374 328170 273430 328226
rect 273498 328170 273554 328226
rect 273622 328170 273678 328226
rect 273250 328046 273306 328102
rect 273374 328046 273430 328102
rect 273498 328046 273554 328102
rect 273622 328046 273678 328102
rect 273250 327922 273306 327978
rect 273374 327922 273430 327978
rect 273498 327922 273554 327978
rect 273622 327922 273678 327978
rect 273250 310294 273306 310350
rect 273374 310294 273430 310350
rect 273498 310294 273554 310350
rect 273622 310294 273678 310350
rect 273250 310170 273306 310226
rect 273374 310170 273430 310226
rect 273498 310170 273554 310226
rect 273622 310170 273678 310226
rect 273250 310046 273306 310102
rect 273374 310046 273430 310102
rect 273498 310046 273554 310102
rect 273622 310046 273678 310102
rect 273250 309922 273306 309978
rect 273374 309922 273430 309978
rect 273498 309922 273554 309978
rect 273622 309922 273678 309978
rect 273250 292294 273306 292350
rect 273374 292294 273430 292350
rect 273498 292294 273554 292350
rect 273622 292294 273678 292350
rect 273250 292170 273306 292226
rect 273374 292170 273430 292226
rect 273498 292170 273554 292226
rect 273622 292170 273678 292226
rect 273250 292046 273306 292102
rect 273374 292046 273430 292102
rect 273498 292046 273554 292102
rect 273622 292046 273678 292102
rect 273250 291922 273306 291978
rect 273374 291922 273430 291978
rect 273498 291922 273554 291978
rect 273622 291922 273678 291978
rect 273250 274294 273306 274350
rect 273374 274294 273430 274350
rect 273498 274294 273554 274350
rect 273622 274294 273678 274350
rect 273250 274170 273306 274226
rect 273374 274170 273430 274226
rect 273498 274170 273554 274226
rect 273622 274170 273678 274226
rect 273250 274046 273306 274102
rect 273374 274046 273430 274102
rect 273498 274046 273554 274102
rect 273622 274046 273678 274102
rect 273250 273922 273306 273978
rect 273374 273922 273430 273978
rect 273498 273922 273554 273978
rect 273622 273922 273678 273978
rect 273250 256294 273306 256350
rect 273374 256294 273430 256350
rect 273498 256294 273554 256350
rect 273622 256294 273678 256350
rect 273250 256170 273306 256226
rect 273374 256170 273430 256226
rect 273498 256170 273554 256226
rect 273622 256170 273678 256226
rect 273250 256046 273306 256102
rect 273374 256046 273430 256102
rect 273498 256046 273554 256102
rect 273622 256046 273678 256102
rect 273250 255922 273306 255978
rect 273374 255922 273430 255978
rect 273498 255922 273554 255978
rect 273622 255922 273678 255978
rect 273250 238294 273306 238350
rect 273374 238294 273430 238350
rect 273498 238294 273554 238350
rect 273622 238294 273678 238350
rect 273250 238170 273306 238226
rect 273374 238170 273430 238226
rect 273498 238170 273554 238226
rect 273622 238170 273678 238226
rect 273250 238046 273306 238102
rect 273374 238046 273430 238102
rect 273498 238046 273554 238102
rect 273622 238046 273678 238102
rect 273250 237922 273306 237978
rect 273374 237922 273430 237978
rect 273498 237922 273554 237978
rect 273622 237922 273678 237978
rect 273250 220294 273306 220350
rect 273374 220294 273430 220350
rect 273498 220294 273554 220350
rect 273622 220294 273678 220350
rect 273250 220170 273306 220226
rect 273374 220170 273430 220226
rect 273498 220170 273554 220226
rect 273622 220170 273678 220226
rect 273250 220046 273306 220102
rect 273374 220046 273430 220102
rect 273498 220046 273554 220102
rect 273622 220046 273678 220102
rect 273250 219922 273306 219978
rect 273374 219922 273430 219978
rect 273498 219922 273554 219978
rect 273622 219922 273678 219978
rect 258970 208294 259026 208350
rect 259094 208294 259150 208350
rect 259218 208294 259274 208350
rect 259342 208294 259398 208350
rect 258970 208170 259026 208226
rect 259094 208170 259150 208226
rect 259218 208170 259274 208226
rect 259342 208170 259398 208226
rect 258970 208046 259026 208102
rect 259094 208046 259150 208102
rect 259218 208046 259274 208102
rect 259342 208046 259398 208102
rect 258970 207922 259026 207978
rect 259094 207922 259150 207978
rect 259218 207922 259274 207978
rect 259342 207922 259398 207978
rect 255250 184294 255306 184350
rect 255374 184294 255430 184350
rect 255498 184294 255554 184350
rect 255622 184294 255678 184350
rect 255250 184170 255306 184226
rect 255374 184170 255430 184226
rect 255498 184170 255554 184226
rect 255622 184170 255678 184226
rect 255250 184046 255306 184102
rect 255374 184046 255430 184102
rect 255498 184046 255554 184102
rect 255622 184046 255678 184102
rect 255250 183922 255306 183978
rect 255374 183922 255430 183978
rect 255498 183922 255554 183978
rect 255622 183922 255678 183978
rect 255250 166294 255306 166350
rect 255374 166294 255430 166350
rect 255498 166294 255554 166350
rect 255622 166294 255678 166350
rect 255250 166170 255306 166226
rect 255374 166170 255430 166226
rect 255498 166170 255554 166226
rect 255622 166170 255678 166226
rect 255250 166046 255306 166102
rect 255374 166046 255430 166102
rect 255498 166046 255554 166102
rect 255622 166046 255678 166102
rect 255250 165922 255306 165978
rect 255374 165922 255430 165978
rect 255498 165922 255554 165978
rect 255622 165922 255678 165978
rect 258970 190294 259026 190350
rect 259094 190294 259150 190350
rect 259218 190294 259274 190350
rect 259342 190294 259398 190350
rect 258970 190170 259026 190226
rect 259094 190170 259150 190226
rect 259218 190170 259274 190226
rect 259342 190170 259398 190226
rect 258970 190046 259026 190102
rect 259094 190046 259150 190102
rect 259218 190046 259274 190102
rect 259342 190046 259398 190102
rect 258970 189922 259026 189978
rect 259094 189922 259150 189978
rect 259218 189922 259274 189978
rect 259342 189922 259398 189978
rect 258970 172294 259026 172350
rect 259094 172294 259150 172350
rect 259218 172294 259274 172350
rect 259342 172294 259398 172350
rect 258970 172170 259026 172226
rect 259094 172170 259150 172226
rect 259218 172170 259274 172226
rect 259342 172170 259398 172226
rect 258970 172046 259026 172102
rect 259094 172046 259150 172102
rect 259218 172046 259274 172102
rect 259342 172046 259398 172102
rect 258970 171922 259026 171978
rect 259094 171922 259150 171978
rect 259218 171922 259274 171978
rect 259342 171922 259398 171978
rect 255250 148294 255306 148350
rect 255374 148294 255430 148350
rect 255498 148294 255554 148350
rect 255622 148294 255678 148350
rect 255250 148170 255306 148226
rect 255374 148170 255430 148226
rect 255498 148170 255554 148226
rect 255622 148170 255678 148226
rect 255250 148046 255306 148102
rect 255374 148046 255430 148102
rect 255498 148046 255554 148102
rect 255622 148046 255678 148102
rect 255250 147922 255306 147978
rect 255374 147922 255430 147978
rect 255498 147922 255554 147978
rect 255622 147922 255678 147978
rect 258970 154294 259026 154350
rect 259094 154294 259150 154350
rect 259218 154294 259274 154350
rect 259342 154294 259398 154350
rect 258970 154170 259026 154226
rect 259094 154170 259150 154226
rect 259218 154170 259274 154226
rect 259342 154170 259398 154226
rect 258970 154046 259026 154102
rect 259094 154046 259150 154102
rect 259218 154046 259274 154102
rect 259342 154046 259398 154102
rect 258970 153922 259026 153978
rect 259094 153922 259150 153978
rect 259218 153922 259274 153978
rect 259342 153922 259398 153978
rect 258970 136294 259026 136350
rect 259094 136294 259150 136350
rect 259218 136294 259274 136350
rect 259342 136294 259398 136350
rect 258970 136170 259026 136226
rect 259094 136170 259150 136226
rect 259218 136170 259274 136226
rect 259342 136170 259398 136226
rect 258970 136046 259026 136102
rect 259094 136046 259150 136102
rect 259218 136046 259274 136102
rect 259342 136046 259398 136102
rect 258970 135922 259026 135978
rect 259094 135922 259150 135978
rect 259218 135922 259274 135978
rect 259342 135922 259398 135978
rect 255250 130294 255306 130350
rect 255374 130294 255430 130350
rect 255498 130294 255554 130350
rect 255622 130294 255678 130350
rect 255250 130170 255306 130226
rect 255374 130170 255430 130226
rect 255498 130170 255554 130226
rect 255622 130170 255678 130226
rect 255250 130046 255306 130102
rect 255374 130046 255430 130102
rect 255498 130046 255554 130102
rect 255622 130046 255678 130102
rect 255250 129922 255306 129978
rect 255374 129922 255430 129978
rect 255498 129922 255554 129978
rect 255622 129922 255678 129978
rect 276970 598116 277026 598172
rect 277094 598116 277150 598172
rect 277218 598116 277274 598172
rect 277342 598116 277398 598172
rect 276970 597992 277026 598048
rect 277094 597992 277150 598048
rect 277218 597992 277274 598048
rect 277342 597992 277398 598048
rect 276970 597868 277026 597924
rect 277094 597868 277150 597924
rect 277218 597868 277274 597924
rect 277342 597868 277398 597924
rect 276970 597744 277026 597800
rect 277094 597744 277150 597800
rect 277218 597744 277274 597800
rect 277342 597744 277398 597800
rect 276970 586294 277026 586350
rect 277094 586294 277150 586350
rect 277218 586294 277274 586350
rect 277342 586294 277398 586350
rect 276970 586170 277026 586226
rect 277094 586170 277150 586226
rect 277218 586170 277274 586226
rect 277342 586170 277398 586226
rect 276970 586046 277026 586102
rect 277094 586046 277150 586102
rect 277218 586046 277274 586102
rect 277342 586046 277398 586102
rect 276970 585922 277026 585978
rect 277094 585922 277150 585978
rect 277218 585922 277274 585978
rect 277342 585922 277398 585978
rect 276970 568294 277026 568350
rect 277094 568294 277150 568350
rect 277218 568294 277274 568350
rect 277342 568294 277398 568350
rect 276970 568170 277026 568226
rect 277094 568170 277150 568226
rect 277218 568170 277274 568226
rect 277342 568170 277398 568226
rect 276970 568046 277026 568102
rect 277094 568046 277150 568102
rect 277218 568046 277274 568102
rect 277342 568046 277398 568102
rect 276970 567922 277026 567978
rect 277094 567922 277150 567978
rect 277218 567922 277274 567978
rect 277342 567922 277398 567978
rect 276970 550294 277026 550350
rect 277094 550294 277150 550350
rect 277218 550294 277274 550350
rect 277342 550294 277398 550350
rect 276970 550170 277026 550226
rect 277094 550170 277150 550226
rect 277218 550170 277274 550226
rect 277342 550170 277398 550226
rect 276970 550046 277026 550102
rect 277094 550046 277150 550102
rect 277218 550046 277274 550102
rect 277342 550046 277398 550102
rect 276970 549922 277026 549978
rect 277094 549922 277150 549978
rect 277218 549922 277274 549978
rect 277342 549922 277398 549978
rect 276970 532294 277026 532350
rect 277094 532294 277150 532350
rect 277218 532294 277274 532350
rect 277342 532294 277398 532350
rect 276970 532170 277026 532226
rect 277094 532170 277150 532226
rect 277218 532170 277274 532226
rect 277342 532170 277398 532226
rect 276970 532046 277026 532102
rect 277094 532046 277150 532102
rect 277218 532046 277274 532102
rect 277342 532046 277398 532102
rect 276970 531922 277026 531978
rect 277094 531922 277150 531978
rect 277218 531922 277274 531978
rect 277342 531922 277398 531978
rect 276970 514294 277026 514350
rect 277094 514294 277150 514350
rect 277218 514294 277274 514350
rect 277342 514294 277398 514350
rect 276970 514170 277026 514226
rect 277094 514170 277150 514226
rect 277218 514170 277274 514226
rect 277342 514170 277398 514226
rect 276970 514046 277026 514102
rect 277094 514046 277150 514102
rect 277218 514046 277274 514102
rect 277342 514046 277398 514102
rect 276970 513922 277026 513978
rect 277094 513922 277150 513978
rect 277218 513922 277274 513978
rect 277342 513922 277398 513978
rect 276970 496294 277026 496350
rect 277094 496294 277150 496350
rect 277218 496294 277274 496350
rect 277342 496294 277398 496350
rect 276970 496170 277026 496226
rect 277094 496170 277150 496226
rect 277218 496170 277274 496226
rect 277342 496170 277398 496226
rect 276970 496046 277026 496102
rect 277094 496046 277150 496102
rect 277218 496046 277274 496102
rect 277342 496046 277398 496102
rect 276970 495922 277026 495978
rect 277094 495922 277150 495978
rect 277218 495922 277274 495978
rect 277342 495922 277398 495978
rect 276970 478294 277026 478350
rect 277094 478294 277150 478350
rect 277218 478294 277274 478350
rect 277342 478294 277398 478350
rect 276970 478170 277026 478226
rect 277094 478170 277150 478226
rect 277218 478170 277274 478226
rect 277342 478170 277398 478226
rect 276970 478046 277026 478102
rect 277094 478046 277150 478102
rect 277218 478046 277274 478102
rect 277342 478046 277398 478102
rect 276970 477922 277026 477978
rect 277094 477922 277150 477978
rect 277218 477922 277274 477978
rect 277342 477922 277398 477978
rect 276970 460294 277026 460350
rect 277094 460294 277150 460350
rect 277218 460294 277274 460350
rect 277342 460294 277398 460350
rect 276970 460170 277026 460226
rect 277094 460170 277150 460226
rect 277218 460170 277274 460226
rect 277342 460170 277398 460226
rect 276970 460046 277026 460102
rect 277094 460046 277150 460102
rect 277218 460046 277274 460102
rect 277342 460046 277398 460102
rect 276970 459922 277026 459978
rect 277094 459922 277150 459978
rect 277218 459922 277274 459978
rect 277342 459922 277398 459978
rect 276970 442294 277026 442350
rect 277094 442294 277150 442350
rect 277218 442294 277274 442350
rect 277342 442294 277398 442350
rect 276970 442170 277026 442226
rect 277094 442170 277150 442226
rect 277218 442170 277274 442226
rect 277342 442170 277398 442226
rect 276970 442046 277026 442102
rect 277094 442046 277150 442102
rect 277218 442046 277274 442102
rect 277342 442046 277398 442102
rect 276970 441922 277026 441978
rect 277094 441922 277150 441978
rect 277218 441922 277274 441978
rect 277342 441922 277398 441978
rect 276970 424294 277026 424350
rect 277094 424294 277150 424350
rect 277218 424294 277274 424350
rect 277342 424294 277398 424350
rect 276970 424170 277026 424226
rect 277094 424170 277150 424226
rect 277218 424170 277274 424226
rect 277342 424170 277398 424226
rect 276970 424046 277026 424102
rect 277094 424046 277150 424102
rect 277218 424046 277274 424102
rect 277342 424046 277398 424102
rect 276970 423922 277026 423978
rect 277094 423922 277150 423978
rect 277218 423922 277274 423978
rect 277342 423922 277398 423978
rect 276970 406294 277026 406350
rect 277094 406294 277150 406350
rect 277218 406294 277274 406350
rect 277342 406294 277398 406350
rect 276970 406170 277026 406226
rect 277094 406170 277150 406226
rect 277218 406170 277274 406226
rect 277342 406170 277398 406226
rect 276970 406046 277026 406102
rect 277094 406046 277150 406102
rect 277218 406046 277274 406102
rect 277342 406046 277398 406102
rect 276970 405922 277026 405978
rect 277094 405922 277150 405978
rect 277218 405922 277274 405978
rect 277342 405922 277398 405978
rect 276970 388294 277026 388350
rect 277094 388294 277150 388350
rect 277218 388294 277274 388350
rect 277342 388294 277398 388350
rect 276970 388170 277026 388226
rect 277094 388170 277150 388226
rect 277218 388170 277274 388226
rect 277342 388170 277398 388226
rect 276970 388046 277026 388102
rect 277094 388046 277150 388102
rect 277218 388046 277274 388102
rect 277342 388046 277398 388102
rect 276970 387922 277026 387978
rect 277094 387922 277150 387978
rect 277218 387922 277274 387978
rect 277342 387922 277398 387978
rect 276970 370294 277026 370350
rect 277094 370294 277150 370350
rect 277218 370294 277274 370350
rect 277342 370294 277398 370350
rect 276970 370170 277026 370226
rect 277094 370170 277150 370226
rect 277218 370170 277274 370226
rect 277342 370170 277398 370226
rect 276970 370046 277026 370102
rect 277094 370046 277150 370102
rect 277218 370046 277274 370102
rect 277342 370046 277398 370102
rect 276970 369922 277026 369978
rect 277094 369922 277150 369978
rect 277218 369922 277274 369978
rect 277342 369922 277398 369978
rect 276970 352294 277026 352350
rect 277094 352294 277150 352350
rect 277218 352294 277274 352350
rect 277342 352294 277398 352350
rect 276970 352170 277026 352226
rect 277094 352170 277150 352226
rect 277218 352170 277274 352226
rect 277342 352170 277398 352226
rect 276970 352046 277026 352102
rect 277094 352046 277150 352102
rect 277218 352046 277274 352102
rect 277342 352046 277398 352102
rect 276970 351922 277026 351978
rect 277094 351922 277150 351978
rect 277218 351922 277274 351978
rect 277342 351922 277398 351978
rect 276970 334294 277026 334350
rect 277094 334294 277150 334350
rect 277218 334294 277274 334350
rect 277342 334294 277398 334350
rect 276970 334170 277026 334226
rect 277094 334170 277150 334226
rect 277218 334170 277274 334226
rect 277342 334170 277398 334226
rect 276970 334046 277026 334102
rect 277094 334046 277150 334102
rect 277218 334046 277274 334102
rect 277342 334046 277398 334102
rect 276970 333922 277026 333978
rect 277094 333922 277150 333978
rect 277218 333922 277274 333978
rect 277342 333922 277398 333978
rect 276970 316294 277026 316350
rect 277094 316294 277150 316350
rect 277218 316294 277274 316350
rect 277342 316294 277398 316350
rect 276970 316170 277026 316226
rect 277094 316170 277150 316226
rect 277218 316170 277274 316226
rect 277342 316170 277398 316226
rect 276970 316046 277026 316102
rect 277094 316046 277150 316102
rect 277218 316046 277274 316102
rect 277342 316046 277398 316102
rect 276970 315922 277026 315978
rect 277094 315922 277150 315978
rect 277218 315922 277274 315978
rect 277342 315922 277398 315978
rect 276970 298294 277026 298350
rect 277094 298294 277150 298350
rect 277218 298294 277274 298350
rect 277342 298294 277398 298350
rect 276970 298170 277026 298226
rect 277094 298170 277150 298226
rect 277218 298170 277274 298226
rect 277342 298170 277398 298226
rect 276970 298046 277026 298102
rect 277094 298046 277150 298102
rect 277218 298046 277274 298102
rect 277342 298046 277398 298102
rect 276970 297922 277026 297978
rect 277094 297922 277150 297978
rect 277218 297922 277274 297978
rect 277342 297922 277398 297978
rect 276970 280294 277026 280350
rect 277094 280294 277150 280350
rect 277218 280294 277274 280350
rect 277342 280294 277398 280350
rect 276970 280170 277026 280226
rect 277094 280170 277150 280226
rect 277218 280170 277274 280226
rect 277342 280170 277398 280226
rect 276970 280046 277026 280102
rect 277094 280046 277150 280102
rect 277218 280046 277274 280102
rect 277342 280046 277398 280102
rect 276970 279922 277026 279978
rect 277094 279922 277150 279978
rect 277218 279922 277274 279978
rect 277342 279922 277398 279978
rect 276970 262294 277026 262350
rect 277094 262294 277150 262350
rect 277218 262294 277274 262350
rect 277342 262294 277398 262350
rect 276970 262170 277026 262226
rect 277094 262170 277150 262226
rect 277218 262170 277274 262226
rect 277342 262170 277398 262226
rect 276970 262046 277026 262102
rect 277094 262046 277150 262102
rect 277218 262046 277274 262102
rect 277342 262046 277398 262102
rect 276970 261922 277026 261978
rect 277094 261922 277150 261978
rect 277218 261922 277274 261978
rect 277342 261922 277398 261978
rect 276970 244294 277026 244350
rect 277094 244294 277150 244350
rect 277218 244294 277274 244350
rect 277342 244294 277398 244350
rect 276970 244170 277026 244226
rect 277094 244170 277150 244226
rect 277218 244170 277274 244226
rect 277342 244170 277398 244226
rect 276970 244046 277026 244102
rect 277094 244046 277150 244102
rect 277218 244046 277274 244102
rect 277342 244046 277398 244102
rect 276970 243922 277026 243978
rect 277094 243922 277150 243978
rect 277218 243922 277274 243978
rect 277342 243922 277398 243978
rect 276970 226294 277026 226350
rect 277094 226294 277150 226350
rect 277218 226294 277274 226350
rect 277342 226294 277398 226350
rect 276970 226170 277026 226226
rect 277094 226170 277150 226226
rect 277218 226170 277274 226226
rect 277342 226170 277398 226226
rect 276970 226046 277026 226102
rect 277094 226046 277150 226102
rect 277218 226046 277274 226102
rect 277342 226046 277398 226102
rect 276970 225922 277026 225978
rect 277094 225922 277150 225978
rect 277218 225922 277274 225978
rect 277342 225922 277398 225978
rect 273250 202294 273306 202350
rect 273374 202294 273430 202350
rect 273498 202294 273554 202350
rect 273622 202294 273678 202350
rect 273250 202170 273306 202226
rect 273374 202170 273430 202226
rect 273498 202170 273554 202226
rect 273622 202170 273678 202226
rect 273250 202046 273306 202102
rect 273374 202046 273430 202102
rect 273498 202046 273554 202102
rect 273622 202046 273678 202102
rect 273250 201922 273306 201978
rect 273374 201922 273430 201978
rect 273498 201922 273554 201978
rect 273622 201922 273678 201978
rect 273250 184294 273306 184350
rect 273374 184294 273430 184350
rect 273498 184294 273554 184350
rect 273622 184294 273678 184350
rect 273250 184170 273306 184226
rect 273374 184170 273430 184226
rect 273498 184170 273554 184226
rect 273622 184170 273678 184226
rect 273250 184046 273306 184102
rect 273374 184046 273430 184102
rect 273498 184046 273554 184102
rect 273622 184046 273678 184102
rect 273250 183922 273306 183978
rect 273374 183922 273430 183978
rect 273498 183922 273554 183978
rect 273622 183922 273678 183978
rect 273250 166294 273306 166350
rect 273374 166294 273430 166350
rect 273498 166294 273554 166350
rect 273622 166294 273678 166350
rect 273250 166170 273306 166226
rect 273374 166170 273430 166226
rect 273498 166170 273554 166226
rect 273622 166170 273678 166226
rect 273250 166046 273306 166102
rect 273374 166046 273430 166102
rect 273498 166046 273554 166102
rect 273622 166046 273678 166102
rect 273250 165922 273306 165978
rect 273374 165922 273430 165978
rect 273498 165922 273554 165978
rect 273622 165922 273678 165978
rect 276970 208294 277026 208350
rect 277094 208294 277150 208350
rect 277218 208294 277274 208350
rect 277342 208294 277398 208350
rect 276970 208170 277026 208226
rect 277094 208170 277150 208226
rect 277218 208170 277274 208226
rect 277342 208170 277398 208226
rect 276970 208046 277026 208102
rect 277094 208046 277150 208102
rect 277218 208046 277274 208102
rect 277342 208046 277398 208102
rect 276970 207922 277026 207978
rect 277094 207922 277150 207978
rect 277218 207922 277274 207978
rect 277342 207922 277398 207978
rect 276970 190294 277026 190350
rect 277094 190294 277150 190350
rect 277218 190294 277274 190350
rect 277342 190294 277398 190350
rect 276970 190170 277026 190226
rect 277094 190170 277150 190226
rect 277218 190170 277274 190226
rect 277342 190170 277398 190226
rect 276970 190046 277026 190102
rect 277094 190046 277150 190102
rect 277218 190046 277274 190102
rect 277342 190046 277398 190102
rect 276970 189922 277026 189978
rect 277094 189922 277150 189978
rect 277218 189922 277274 189978
rect 277342 189922 277398 189978
rect 273250 148294 273306 148350
rect 273374 148294 273430 148350
rect 273498 148294 273554 148350
rect 273622 148294 273678 148350
rect 273250 148170 273306 148226
rect 273374 148170 273430 148226
rect 273498 148170 273554 148226
rect 273622 148170 273678 148226
rect 273250 148046 273306 148102
rect 273374 148046 273430 148102
rect 273498 148046 273554 148102
rect 273622 148046 273678 148102
rect 273250 147922 273306 147978
rect 273374 147922 273430 147978
rect 273498 147922 273554 147978
rect 273622 147922 273678 147978
rect 273250 130294 273306 130350
rect 273374 130294 273430 130350
rect 273498 130294 273554 130350
rect 273622 130294 273678 130350
rect 273250 130170 273306 130226
rect 273374 130170 273430 130226
rect 273498 130170 273554 130226
rect 273622 130170 273678 130226
rect 273250 130046 273306 130102
rect 273374 130046 273430 130102
rect 273498 130046 273554 130102
rect 273622 130046 273678 130102
rect 273250 129922 273306 129978
rect 273374 129922 273430 129978
rect 273498 129922 273554 129978
rect 273622 129922 273678 129978
rect 258970 118294 259026 118350
rect 259094 118294 259150 118350
rect 259218 118294 259274 118350
rect 259342 118294 259398 118350
rect 258970 118170 259026 118226
rect 259094 118170 259150 118226
rect 259218 118170 259274 118226
rect 259342 118170 259398 118226
rect 258970 118046 259026 118102
rect 259094 118046 259150 118102
rect 259218 118046 259274 118102
rect 259342 118046 259398 118102
rect 258970 117922 259026 117978
rect 259094 117922 259150 117978
rect 259218 117922 259274 117978
rect 259342 117922 259398 117978
rect 255250 112294 255306 112350
rect 255374 112294 255430 112350
rect 255498 112294 255554 112350
rect 255622 112294 255678 112350
rect 255250 112170 255306 112226
rect 255374 112170 255430 112226
rect 255498 112170 255554 112226
rect 255622 112170 255678 112226
rect 255250 112046 255306 112102
rect 255374 112046 255430 112102
rect 255498 112046 255554 112102
rect 255622 112046 255678 112102
rect 255250 111922 255306 111978
rect 255374 111922 255430 111978
rect 255498 111922 255554 111978
rect 255622 111922 255678 111978
rect 255250 94294 255306 94350
rect 255374 94294 255430 94350
rect 255498 94294 255554 94350
rect 255622 94294 255678 94350
rect 255250 94170 255306 94226
rect 255374 94170 255430 94226
rect 255498 94170 255554 94226
rect 255622 94170 255678 94226
rect 255250 94046 255306 94102
rect 255374 94046 255430 94102
rect 255498 94046 255554 94102
rect 255622 94046 255678 94102
rect 255250 93922 255306 93978
rect 255374 93922 255430 93978
rect 255498 93922 255554 93978
rect 255622 93922 255678 93978
rect 255250 76294 255306 76350
rect 255374 76294 255430 76350
rect 255498 76294 255554 76350
rect 255622 76294 255678 76350
rect 255250 76170 255306 76226
rect 255374 76170 255430 76226
rect 255498 76170 255554 76226
rect 255622 76170 255678 76226
rect 255250 76046 255306 76102
rect 255374 76046 255430 76102
rect 255498 76046 255554 76102
rect 255622 76046 255678 76102
rect 255250 75922 255306 75978
rect 255374 75922 255430 75978
rect 255498 75922 255554 75978
rect 255622 75922 255678 75978
rect 244412 29582 244468 29638
rect 255250 58294 255306 58350
rect 255374 58294 255430 58350
rect 255498 58294 255554 58350
rect 255622 58294 255678 58350
rect 255250 58170 255306 58226
rect 255374 58170 255430 58226
rect 255498 58170 255554 58226
rect 255622 58170 255678 58226
rect 255250 58046 255306 58102
rect 255374 58046 255430 58102
rect 255498 58046 255554 58102
rect 255622 58046 255678 58102
rect 255250 57922 255306 57978
rect 255374 57922 255430 57978
rect 255498 57922 255554 57978
rect 255622 57922 255678 57978
rect 255250 40294 255306 40350
rect 255374 40294 255430 40350
rect 255498 40294 255554 40350
rect 255622 40294 255678 40350
rect 255250 40170 255306 40226
rect 255374 40170 255430 40226
rect 255498 40170 255554 40226
rect 255622 40170 255678 40226
rect 255250 40046 255306 40102
rect 255374 40046 255430 40102
rect 255498 40046 255554 40102
rect 255622 40046 255678 40102
rect 255250 39922 255306 39978
rect 255374 39922 255430 39978
rect 255498 39922 255554 39978
rect 255622 39922 255678 39978
rect 240970 28294 241026 28350
rect 241094 28294 241150 28350
rect 241218 28294 241274 28350
rect 241342 28294 241398 28350
rect 240970 28170 241026 28226
rect 241094 28170 241150 28226
rect 241218 28170 241274 28226
rect 241342 28170 241398 28226
rect 240970 28046 241026 28102
rect 241094 28046 241150 28102
rect 241218 28046 241274 28102
rect 241342 28046 241398 28102
rect 240970 27922 241026 27978
rect 241094 27922 241150 27978
rect 241218 27922 241274 27978
rect 241342 27922 241398 27978
rect 237250 22294 237306 22350
rect 237374 22294 237430 22350
rect 237498 22294 237554 22350
rect 237622 22294 237678 22350
rect 237250 22170 237306 22226
rect 237374 22170 237430 22226
rect 237498 22170 237554 22226
rect 237622 22170 237678 22226
rect 237250 22046 237306 22102
rect 237374 22046 237430 22102
rect 237498 22046 237554 22102
rect 237622 22046 237678 22102
rect 237250 21922 237306 21978
rect 237374 21922 237430 21978
rect 237498 21922 237554 21978
rect 237622 21922 237678 21978
rect 237250 4294 237306 4350
rect 237374 4294 237430 4350
rect 237498 4294 237554 4350
rect 237622 4294 237678 4350
rect 237250 4170 237306 4226
rect 237374 4170 237430 4226
rect 237498 4170 237554 4226
rect 237622 4170 237678 4226
rect 237250 4046 237306 4102
rect 237374 4046 237430 4102
rect 237498 4046 237554 4102
rect 237622 4046 237678 4102
rect 237250 3922 237306 3978
rect 237374 3922 237430 3978
rect 237498 3922 237554 3978
rect 237622 3922 237678 3978
rect 237250 -216 237306 -160
rect 237374 -216 237430 -160
rect 237498 -216 237554 -160
rect 237622 -216 237678 -160
rect 237250 -340 237306 -284
rect 237374 -340 237430 -284
rect 237498 -340 237554 -284
rect 237622 -340 237678 -284
rect 237250 -464 237306 -408
rect 237374 -464 237430 -408
rect 237498 -464 237554 -408
rect 237622 -464 237678 -408
rect 237250 -588 237306 -532
rect 237374 -588 237430 -532
rect 237498 -588 237554 -532
rect 237622 -588 237678 -532
rect 240970 10294 241026 10350
rect 241094 10294 241150 10350
rect 241218 10294 241274 10350
rect 241342 10294 241398 10350
rect 240970 10170 241026 10226
rect 241094 10170 241150 10226
rect 241218 10170 241274 10226
rect 241342 10170 241398 10226
rect 240970 10046 241026 10102
rect 241094 10046 241150 10102
rect 241218 10046 241274 10102
rect 241342 10046 241398 10102
rect 240970 9922 241026 9978
rect 241094 9922 241150 9978
rect 241218 9922 241274 9978
rect 241342 9922 241398 9978
rect 240970 -1176 241026 -1120
rect 241094 -1176 241150 -1120
rect 241218 -1176 241274 -1120
rect 241342 -1176 241398 -1120
rect 240970 -1300 241026 -1244
rect 241094 -1300 241150 -1244
rect 241218 -1300 241274 -1244
rect 241342 -1300 241398 -1244
rect 240970 -1424 241026 -1368
rect 241094 -1424 241150 -1368
rect 241218 -1424 241274 -1368
rect 241342 -1424 241398 -1368
rect 240970 -1548 241026 -1492
rect 241094 -1548 241150 -1492
rect 241218 -1548 241274 -1492
rect 241342 -1548 241398 -1492
rect 255250 22294 255306 22350
rect 255374 22294 255430 22350
rect 255498 22294 255554 22350
rect 255622 22294 255678 22350
rect 255250 22170 255306 22226
rect 255374 22170 255430 22226
rect 255498 22170 255554 22226
rect 255622 22170 255678 22226
rect 255250 22046 255306 22102
rect 255374 22046 255430 22102
rect 255498 22046 255554 22102
rect 255622 22046 255678 22102
rect 255250 21922 255306 21978
rect 255374 21922 255430 21978
rect 255498 21922 255554 21978
rect 255622 21922 255678 21978
rect 255250 4294 255306 4350
rect 255374 4294 255430 4350
rect 255498 4294 255554 4350
rect 255622 4294 255678 4350
rect 255250 4170 255306 4226
rect 255374 4170 255430 4226
rect 255498 4170 255554 4226
rect 255622 4170 255678 4226
rect 255250 4046 255306 4102
rect 255374 4046 255430 4102
rect 255498 4046 255554 4102
rect 255622 4046 255678 4102
rect 255250 3922 255306 3978
rect 255374 3922 255430 3978
rect 255498 3922 255554 3978
rect 255622 3922 255678 3978
rect 255250 -216 255306 -160
rect 255374 -216 255430 -160
rect 255498 -216 255554 -160
rect 255622 -216 255678 -160
rect 255250 -340 255306 -284
rect 255374 -340 255430 -284
rect 255498 -340 255554 -284
rect 255622 -340 255678 -284
rect 255250 -464 255306 -408
rect 255374 -464 255430 -408
rect 255498 -464 255554 -408
rect 255622 -464 255678 -408
rect 255250 -588 255306 -532
rect 255374 -588 255430 -532
rect 255498 -588 255554 -532
rect 255622 -588 255678 -532
rect 258970 100294 259026 100350
rect 259094 100294 259150 100350
rect 259218 100294 259274 100350
rect 259342 100294 259398 100350
rect 258970 100170 259026 100226
rect 259094 100170 259150 100226
rect 259218 100170 259274 100226
rect 259342 100170 259398 100226
rect 258970 100046 259026 100102
rect 259094 100046 259150 100102
rect 259218 100046 259274 100102
rect 259342 100046 259398 100102
rect 258970 99922 259026 99978
rect 259094 99922 259150 99978
rect 259218 99922 259274 99978
rect 259342 99922 259398 99978
rect 258970 82294 259026 82350
rect 259094 82294 259150 82350
rect 259218 82294 259274 82350
rect 259342 82294 259398 82350
rect 258970 82170 259026 82226
rect 259094 82170 259150 82226
rect 259218 82170 259274 82226
rect 259342 82170 259398 82226
rect 258970 82046 259026 82102
rect 259094 82046 259150 82102
rect 259218 82046 259274 82102
rect 259342 82046 259398 82102
rect 258970 81922 259026 81978
rect 259094 81922 259150 81978
rect 259218 81922 259274 81978
rect 259342 81922 259398 81978
rect 258970 64294 259026 64350
rect 259094 64294 259150 64350
rect 259218 64294 259274 64350
rect 259342 64294 259398 64350
rect 258970 64170 259026 64226
rect 259094 64170 259150 64226
rect 259218 64170 259274 64226
rect 259342 64170 259398 64226
rect 258970 64046 259026 64102
rect 259094 64046 259150 64102
rect 259218 64046 259274 64102
rect 259342 64046 259398 64102
rect 258970 63922 259026 63978
rect 259094 63922 259150 63978
rect 259218 63922 259274 63978
rect 259342 63922 259398 63978
rect 258970 46294 259026 46350
rect 259094 46294 259150 46350
rect 259218 46294 259274 46350
rect 259342 46294 259398 46350
rect 258970 46170 259026 46226
rect 259094 46170 259150 46226
rect 259218 46170 259274 46226
rect 259342 46170 259398 46226
rect 258970 46046 259026 46102
rect 259094 46046 259150 46102
rect 259218 46046 259274 46102
rect 259342 46046 259398 46102
rect 258970 45922 259026 45978
rect 259094 45922 259150 45978
rect 259218 45922 259274 45978
rect 259342 45922 259398 45978
rect 258970 28294 259026 28350
rect 259094 28294 259150 28350
rect 259218 28294 259274 28350
rect 259342 28294 259398 28350
rect 258970 28170 259026 28226
rect 259094 28170 259150 28226
rect 259218 28170 259274 28226
rect 259342 28170 259398 28226
rect 258970 28046 259026 28102
rect 259094 28046 259150 28102
rect 259218 28046 259274 28102
rect 259342 28046 259398 28102
rect 258970 27922 259026 27978
rect 259094 27922 259150 27978
rect 259218 27922 259274 27978
rect 259342 27922 259398 27978
rect 258970 10294 259026 10350
rect 259094 10294 259150 10350
rect 259218 10294 259274 10350
rect 259342 10294 259398 10350
rect 258970 10170 259026 10226
rect 259094 10170 259150 10226
rect 259218 10170 259274 10226
rect 259342 10170 259398 10226
rect 258970 10046 259026 10102
rect 259094 10046 259150 10102
rect 259218 10046 259274 10102
rect 259342 10046 259398 10102
rect 258970 9922 259026 9978
rect 259094 9922 259150 9978
rect 259218 9922 259274 9978
rect 259342 9922 259398 9978
rect 258970 -1176 259026 -1120
rect 259094 -1176 259150 -1120
rect 259218 -1176 259274 -1120
rect 259342 -1176 259398 -1120
rect 258970 -1300 259026 -1244
rect 259094 -1300 259150 -1244
rect 259218 -1300 259274 -1244
rect 259342 -1300 259398 -1244
rect 258970 -1424 259026 -1368
rect 259094 -1424 259150 -1368
rect 259218 -1424 259274 -1368
rect 259342 -1424 259398 -1368
rect 258970 -1548 259026 -1492
rect 259094 -1548 259150 -1492
rect 259218 -1548 259274 -1492
rect 259342 -1548 259398 -1492
rect 276970 172294 277026 172350
rect 277094 172294 277150 172350
rect 277218 172294 277274 172350
rect 277342 172294 277398 172350
rect 276970 172170 277026 172226
rect 277094 172170 277150 172226
rect 277218 172170 277274 172226
rect 277342 172170 277398 172226
rect 276970 172046 277026 172102
rect 277094 172046 277150 172102
rect 277218 172046 277274 172102
rect 277342 172046 277398 172102
rect 276970 171922 277026 171978
rect 277094 171922 277150 171978
rect 277218 171922 277274 171978
rect 277342 171922 277398 171978
rect 291250 597156 291306 597212
rect 291374 597156 291430 597212
rect 291498 597156 291554 597212
rect 291622 597156 291678 597212
rect 291250 597032 291306 597088
rect 291374 597032 291430 597088
rect 291498 597032 291554 597088
rect 291622 597032 291678 597088
rect 291250 596908 291306 596964
rect 291374 596908 291430 596964
rect 291498 596908 291554 596964
rect 291622 596908 291678 596964
rect 291250 596784 291306 596840
rect 291374 596784 291430 596840
rect 291498 596784 291554 596840
rect 291622 596784 291678 596840
rect 291250 580294 291306 580350
rect 291374 580294 291430 580350
rect 291498 580294 291554 580350
rect 291622 580294 291678 580350
rect 291250 580170 291306 580226
rect 291374 580170 291430 580226
rect 291498 580170 291554 580226
rect 291622 580170 291678 580226
rect 291250 580046 291306 580102
rect 291374 580046 291430 580102
rect 291498 580046 291554 580102
rect 291622 580046 291678 580102
rect 291250 579922 291306 579978
rect 291374 579922 291430 579978
rect 291498 579922 291554 579978
rect 291622 579922 291678 579978
rect 291250 562294 291306 562350
rect 291374 562294 291430 562350
rect 291498 562294 291554 562350
rect 291622 562294 291678 562350
rect 291250 562170 291306 562226
rect 291374 562170 291430 562226
rect 291498 562170 291554 562226
rect 291622 562170 291678 562226
rect 291250 562046 291306 562102
rect 291374 562046 291430 562102
rect 291498 562046 291554 562102
rect 291622 562046 291678 562102
rect 291250 561922 291306 561978
rect 291374 561922 291430 561978
rect 291498 561922 291554 561978
rect 291622 561922 291678 561978
rect 291250 544294 291306 544350
rect 291374 544294 291430 544350
rect 291498 544294 291554 544350
rect 291622 544294 291678 544350
rect 291250 544170 291306 544226
rect 291374 544170 291430 544226
rect 291498 544170 291554 544226
rect 291622 544170 291678 544226
rect 291250 544046 291306 544102
rect 291374 544046 291430 544102
rect 291498 544046 291554 544102
rect 291622 544046 291678 544102
rect 291250 543922 291306 543978
rect 291374 543922 291430 543978
rect 291498 543922 291554 543978
rect 291622 543922 291678 543978
rect 291250 526294 291306 526350
rect 291374 526294 291430 526350
rect 291498 526294 291554 526350
rect 291622 526294 291678 526350
rect 291250 526170 291306 526226
rect 291374 526170 291430 526226
rect 291498 526170 291554 526226
rect 291622 526170 291678 526226
rect 291250 526046 291306 526102
rect 291374 526046 291430 526102
rect 291498 526046 291554 526102
rect 291622 526046 291678 526102
rect 291250 525922 291306 525978
rect 291374 525922 291430 525978
rect 291498 525922 291554 525978
rect 291622 525922 291678 525978
rect 291250 508294 291306 508350
rect 291374 508294 291430 508350
rect 291498 508294 291554 508350
rect 291622 508294 291678 508350
rect 291250 508170 291306 508226
rect 291374 508170 291430 508226
rect 291498 508170 291554 508226
rect 291622 508170 291678 508226
rect 291250 508046 291306 508102
rect 291374 508046 291430 508102
rect 291498 508046 291554 508102
rect 291622 508046 291678 508102
rect 291250 507922 291306 507978
rect 291374 507922 291430 507978
rect 291498 507922 291554 507978
rect 291622 507922 291678 507978
rect 291250 490294 291306 490350
rect 291374 490294 291430 490350
rect 291498 490294 291554 490350
rect 291622 490294 291678 490350
rect 291250 490170 291306 490226
rect 291374 490170 291430 490226
rect 291498 490170 291554 490226
rect 291622 490170 291678 490226
rect 291250 490046 291306 490102
rect 291374 490046 291430 490102
rect 291498 490046 291554 490102
rect 291622 490046 291678 490102
rect 291250 489922 291306 489978
rect 291374 489922 291430 489978
rect 291498 489922 291554 489978
rect 291622 489922 291678 489978
rect 291250 472294 291306 472350
rect 291374 472294 291430 472350
rect 291498 472294 291554 472350
rect 291622 472294 291678 472350
rect 291250 472170 291306 472226
rect 291374 472170 291430 472226
rect 291498 472170 291554 472226
rect 291622 472170 291678 472226
rect 291250 472046 291306 472102
rect 291374 472046 291430 472102
rect 291498 472046 291554 472102
rect 291622 472046 291678 472102
rect 291250 471922 291306 471978
rect 291374 471922 291430 471978
rect 291498 471922 291554 471978
rect 291622 471922 291678 471978
rect 291250 454294 291306 454350
rect 291374 454294 291430 454350
rect 291498 454294 291554 454350
rect 291622 454294 291678 454350
rect 291250 454170 291306 454226
rect 291374 454170 291430 454226
rect 291498 454170 291554 454226
rect 291622 454170 291678 454226
rect 291250 454046 291306 454102
rect 291374 454046 291430 454102
rect 291498 454046 291554 454102
rect 291622 454046 291678 454102
rect 291250 453922 291306 453978
rect 291374 453922 291430 453978
rect 291498 453922 291554 453978
rect 291622 453922 291678 453978
rect 291250 436294 291306 436350
rect 291374 436294 291430 436350
rect 291498 436294 291554 436350
rect 291622 436294 291678 436350
rect 291250 436170 291306 436226
rect 291374 436170 291430 436226
rect 291498 436170 291554 436226
rect 291622 436170 291678 436226
rect 291250 436046 291306 436102
rect 291374 436046 291430 436102
rect 291498 436046 291554 436102
rect 291622 436046 291678 436102
rect 291250 435922 291306 435978
rect 291374 435922 291430 435978
rect 291498 435922 291554 435978
rect 291622 435922 291678 435978
rect 291250 418294 291306 418350
rect 291374 418294 291430 418350
rect 291498 418294 291554 418350
rect 291622 418294 291678 418350
rect 291250 418170 291306 418226
rect 291374 418170 291430 418226
rect 291498 418170 291554 418226
rect 291622 418170 291678 418226
rect 291250 418046 291306 418102
rect 291374 418046 291430 418102
rect 291498 418046 291554 418102
rect 291622 418046 291678 418102
rect 291250 417922 291306 417978
rect 291374 417922 291430 417978
rect 291498 417922 291554 417978
rect 291622 417922 291678 417978
rect 291250 400294 291306 400350
rect 291374 400294 291430 400350
rect 291498 400294 291554 400350
rect 291622 400294 291678 400350
rect 291250 400170 291306 400226
rect 291374 400170 291430 400226
rect 291498 400170 291554 400226
rect 291622 400170 291678 400226
rect 291250 400046 291306 400102
rect 291374 400046 291430 400102
rect 291498 400046 291554 400102
rect 291622 400046 291678 400102
rect 291250 399922 291306 399978
rect 291374 399922 291430 399978
rect 291498 399922 291554 399978
rect 291622 399922 291678 399978
rect 291250 382294 291306 382350
rect 291374 382294 291430 382350
rect 291498 382294 291554 382350
rect 291622 382294 291678 382350
rect 291250 382170 291306 382226
rect 291374 382170 291430 382226
rect 291498 382170 291554 382226
rect 291622 382170 291678 382226
rect 291250 382046 291306 382102
rect 291374 382046 291430 382102
rect 291498 382046 291554 382102
rect 291622 382046 291678 382102
rect 291250 381922 291306 381978
rect 291374 381922 291430 381978
rect 291498 381922 291554 381978
rect 291622 381922 291678 381978
rect 291250 364294 291306 364350
rect 291374 364294 291430 364350
rect 291498 364294 291554 364350
rect 291622 364294 291678 364350
rect 291250 364170 291306 364226
rect 291374 364170 291430 364226
rect 291498 364170 291554 364226
rect 291622 364170 291678 364226
rect 291250 364046 291306 364102
rect 291374 364046 291430 364102
rect 291498 364046 291554 364102
rect 291622 364046 291678 364102
rect 291250 363922 291306 363978
rect 291374 363922 291430 363978
rect 291498 363922 291554 363978
rect 291622 363922 291678 363978
rect 291250 346294 291306 346350
rect 291374 346294 291430 346350
rect 291498 346294 291554 346350
rect 291622 346294 291678 346350
rect 291250 346170 291306 346226
rect 291374 346170 291430 346226
rect 291498 346170 291554 346226
rect 291622 346170 291678 346226
rect 291250 346046 291306 346102
rect 291374 346046 291430 346102
rect 291498 346046 291554 346102
rect 291622 346046 291678 346102
rect 291250 345922 291306 345978
rect 291374 345922 291430 345978
rect 291498 345922 291554 345978
rect 291622 345922 291678 345978
rect 291250 328294 291306 328350
rect 291374 328294 291430 328350
rect 291498 328294 291554 328350
rect 291622 328294 291678 328350
rect 291250 328170 291306 328226
rect 291374 328170 291430 328226
rect 291498 328170 291554 328226
rect 291622 328170 291678 328226
rect 291250 328046 291306 328102
rect 291374 328046 291430 328102
rect 291498 328046 291554 328102
rect 291622 328046 291678 328102
rect 291250 327922 291306 327978
rect 291374 327922 291430 327978
rect 291498 327922 291554 327978
rect 291622 327922 291678 327978
rect 291250 310294 291306 310350
rect 291374 310294 291430 310350
rect 291498 310294 291554 310350
rect 291622 310294 291678 310350
rect 291250 310170 291306 310226
rect 291374 310170 291430 310226
rect 291498 310170 291554 310226
rect 291622 310170 291678 310226
rect 291250 310046 291306 310102
rect 291374 310046 291430 310102
rect 291498 310046 291554 310102
rect 291622 310046 291678 310102
rect 291250 309922 291306 309978
rect 291374 309922 291430 309978
rect 291498 309922 291554 309978
rect 291622 309922 291678 309978
rect 291250 292294 291306 292350
rect 291374 292294 291430 292350
rect 291498 292294 291554 292350
rect 291622 292294 291678 292350
rect 291250 292170 291306 292226
rect 291374 292170 291430 292226
rect 291498 292170 291554 292226
rect 291622 292170 291678 292226
rect 291250 292046 291306 292102
rect 291374 292046 291430 292102
rect 291498 292046 291554 292102
rect 291622 292046 291678 292102
rect 291250 291922 291306 291978
rect 291374 291922 291430 291978
rect 291498 291922 291554 291978
rect 291622 291922 291678 291978
rect 291250 274294 291306 274350
rect 291374 274294 291430 274350
rect 291498 274294 291554 274350
rect 291622 274294 291678 274350
rect 291250 274170 291306 274226
rect 291374 274170 291430 274226
rect 291498 274170 291554 274226
rect 291622 274170 291678 274226
rect 291250 274046 291306 274102
rect 291374 274046 291430 274102
rect 291498 274046 291554 274102
rect 291622 274046 291678 274102
rect 291250 273922 291306 273978
rect 291374 273922 291430 273978
rect 291498 273922 291554 273978
rect 291622 273922 291678 273978
rect 291250 256294 291306 256350
rect 291374 256294 291430 256350
rect 291498 256294 291554 256350
rect 291622 256294 291678 256350
rect 291250 256170 291306 256226
rect 291374 256170 291430 256226
rect 291498 256170 291554 256226
rect 291622 256170 291678 256226
rect 291250 256046 291306 256102
rect 291374 256046 291430 256102
rect 291498 256046 291554 256102
rect 291622 256046 291678 256102
rect 291250 255922 291306 255978
rect 291374 255922 291430 255978
rect 291498 255922 291554 255978
rect 291622 255922 291678 255978
rect 309250 597156 309306 597212
rect 309374 597156 309430 597212
rect 309498 597156 309554 597212
rect 309622 597156 309678 597212
rect 309250 597032 309306 597088
rect 309374 597032 309430 597088
rect 309498 597032 309554 597088
rect 309622 597032 309678 597088
rect 309250 596908 309306 596964
rect 309374 596908 309430 596964
rect 309498 596908 309554 596964
rect 309622 596908 309678 596964
rect 309250 596784 309306 596840
rect 309374 596784 309430 596840
rect 309498 596784 309554 596840
rect 309622 596784 309678 596840
rect 309250 580294 309306 580350
rect 309374 580294 309430 580350
rect 309498 580294 309554 580350
rect 309622 580294 309678 580350
rect 309250 580170 309306 580226
rect 309374 580170 309430 580226
rect 309498 580170 309554 580226
rect 309622 580170 309678 580226
rect 309250 580046 309306 580102
rect 309374 580046 309430 580102
rect 309498 580046 309554 580102
rect 309622 580046 309678 580102
rect 309250 579922 309306 579978
rect 309374 579922 309430 579978
rect 309498 579922 309554 579978
rect 309622 579922 309678 579978
rect 309250 562294 309306 562350
rect 309374 562294 309430 562350
rect 309498 562294 309554 562350
rect 309622 562294 309678 562350
rect 309250 562170 309306 562226
rect 309374 562170 309430 562226
rect 309498 562170 309554 562226
rect 309622 562170 309678 562226
rect 309250 562046 309306 562102
rect 309374 562046 309430 562102
rect 309498 562046 309554 562102
rect 309622 562046 309678 562102
rect 309250 561922 309306 561978
rect 309374 561922 309430 561978
rect 309498 561922 309554 561978
rect 309622 561922 309678 561978
rect 309250 544294 309306 544350
rect 309374 544294 309430 544350
rect 309498 544294 309554 544350
rect 309622 544294 309678 544350
rect 309250 544170 309306 544226
rect 309374 544170 309430 544226
rect 309498 544170 309554 544226
rect 309622 544170 309678 544226
rect 309250 544046 309306 544102
rect 309374 544046 309430 544102
rect 309498 544046 309554 544102
rect 309622 544046 309678 544102
rect 309250 543922 309306 543978
rect 309374 543922 309430 543978
rect 309498 543922 309554 543978
rect 309622 543922 309678 543978
rect 309250 526294 309306 526350
rect 309374 526294 309430 526350
rect 309498 526294 309554 526350
rect 309622 526294 309678 526350
rect 309250 526170 309306 526226
rect 309374 526170 309430 526226
rect 309498 526170 309554 526226
rect 309622 526170 309678 526226
rect 309250 526046 309306 526102
rect 309374 526046 309430 526102
rect 309498 526046 309554 526102
rect 309622 526046 309678 526102
rect 309250 525922 309306 525978
rect 309374 525922 309430 525978
rect 309498 525922 309554 525978
rect 309622 525922 309678 525978
rect 309250 508294 309306 508350
rect 309374 508294 309430 508350
rect 309498 508294 309554 508350
rect 309622 508294 309678 508350
rect 309250 508170 309306 508226
rect 309374 508170 309430 508226
rect 309498 508170 309554 508226
rect 309622 508170 309678 508226
rect 309250 508046 309306 508102
rect 309374 508046 309430 508102
rect 309498 508046 309554 508102
rect 309622 508046 309678 508102
rect 309250 507922 309306 507978
rect 309374 507922 309430 507978
rect 309498 507922 309554 507978
rect 309622 507922 309678 507978
rect 309250 490294 309306 490350
rect 309374 490294 309430 490350
rect 309498 490294 309554 490350
rect 309622 490294 309678 490350
rect 309250 490170 309306 490226
rect 309374 490170 309430 490226
rect 309498 490170 309554 490226
rect 309622 490170 309678 490226
rect 309250 490046 309306 490102
rect 309374 490046 309430 490102
rect 309498 490046 309554 490102
rect 309622 490046 309678 490102
rect 309250 489922 309306 489978
rect 309374 489922 309430 489978
rect 309498 489922 309554 489978
rect 309622 489922 309678 489978
rect 309250 472294 309306 472350
rect 309374 472294 309430 472350
rect 309498 472294 309554 472350
rect 309622 472294 309678 472350
rect 309250 472170 309306 472226
rect 309374 472170 309430 472226
rect 309498 472170 309554 472226
rect 309622 472170 309678 472226
rect 309250 472046 309306 472102
rect 309374 472046 309430 472102
rect 309498 472046 309554 472102
rect 309622 472046 309678 472102
rect 309250 471922 309306 471978
rect 309374 471922 309430 471978
rect 309498 471922 309554 471978
rect 309622 471922 309678 471978
rect 309250 454294 309306 454350
rect 309374 454294 309430 454350
rect 309498 454294 309554 454350
rect 309622 454294 309678 454350
rect 309250 454170 309306 454226
rect 309374 454170 309430 454226
rect 309498 454170 309554 454226
rect 309622 454170 309678 454226
rect 309250 454046 309306 454102
rect 309374 454046 309430 454102
rect 309498 454046 309554 454102
rect 309622 454046 309678 454102
rect 309250 453922 309306 453978
rect 309374 453922 309430 453978
rect 309498 453922 309554 453978
rect 309622 453922 309678 453978
rect 309250 436294 309306 436350
rect 309374 436294 309430 436350
rect 309498 436294 309554 436350
rect 309622 436294 309678 436350
rect 309250 436170 309306 436226
rect 309374 436170 309430 436226
rect 309498 436170 309554 436226
rect 309622 436170 309678 436226
rect 309250 436046 309306 436102
rect 309374 436046 309430 436102
rect 309498 436046 309554 436102
rect 309622 436046 309678 436102
rect 309250 435922 309306 435978
rect 309374 435922 309430 435978
rect 309498 435922 309554 435978
rect 309622 435922 309678 435978
rect 309250 418294 309306 418350
rect 309374 418294 309430 418350
rect 309498 418294 309554 418350
rect 309622 418294 309678 418350
rect 309250 418170 309306 418226
rect 309374 418170 309430 418226
rect 309498 418170 309554 418226
rect 309622 418170 309678 418226
rect 309250 418046 309306 418102
rect 309374 418046 309430 418102
rect 309498 418046 309554 418102
rect 309622 418046 309678 418102
rect 309250 417922 309306 417978
rect 309374 417922 309430 417978
rect 309498 417922 309554 417978
rect 309622 417922 309678 417978
rect 309250 400294 309306 400350
rect 309374 400294 309430 400350
rect 309498 400294 309554 400350
rect 309622 400294 309678 400350
rect 309250 400170 309306 400226
rect 309374 400170 309430 400226
rect 309498 400170 309554 400226
rect 309622 400170 309678 400226
rect 309250 400046 309306 400102
rect 309374 400046 309430 400102
rect 309498 400046 309554 400102
rect 309622 400046 309678 400102
rect 309250 399922 309306 399978
rect 309374 399922 309430 399978
rect 309498 399922 309554 399978
rect 309622 399922 309678 399978
rect 309250 382294 309306 382350
rect 309374 382294 309430 382350
rect 309498 382294 309554 382350
rect 309622 382294 309678 382350
rect 309250 382170 309306 382226
rect 309374 382170 309430 382226
rect 309498 382170 309554 382226
rect 309622 382170 309678 382226
rect 309250 382046 309306 382102
rect 309374 382046 309430 382102
rect 309498 382046 309554 382102
rect 309622 382046 309678 382102
rect 309250 381922 309306 381978
rect 309374 381922 309430 381978
rect 309498 381922 309554 381978
rect 309622 381922 309678 381978
rect 309250 364294 309306 364350
rect 309374 364294 309430 364350
rect 309498 364294 309554 364350
rect 309622 364294 309678 364350
rect 309250 364170 309306 364226
rect 309374 364170 309430 364226
rect 309498 364170 309554 364226
rect 309622 364170 309678 364226
rect 309250 364046 309306 364102
rect 309374 364046 309430 364102
rect 309498 364046 309554 364102
rect 309622 364046 309678 364102
rect 309250 363922 309306 363978
rect 309374 363922 309430 363978
rect 309498 363922 309554 363978
rect 309622 363922 309678 363978
rect 309250 346294 309306 346350
rect 309374 346294 309430 346350
rect 309498 346294 309554 346350
rect 309622 346294 309678 346350
rect 309250 346170 309306 346226
rect 309374 346170 309430 346226
rect 309498 346170 309554 346226
rect 309622 346170 309678 346226
rect 309250 346046 309306 346102
rect 309374 346046 309430 346102
rect 309498 346046 309554 346102
rect 309622 346046 309678 346102
rect 309250 345922 309306 345978
rect 309374 345922 309430 345978
rect 309498 345922 309554 345978
rect 309622 345922 309678 345978
rect 309250 328294 309306 328350
rect 309374 328294 309430 328350
rect 309498 328294 309554 328350
rect 309622 328294 309678 328350
rect 309250 328170 309306 328226
rect 309374 328170 309430 328226
rect 309498 328170 309554 328226
rect 309622 328170 309678 328226
rect 309250 328046 309306 328102
rect 309374 328046 309430 328102
rect 309498 328046 309554 328102
rect 309622 328046 309678 328102
rect 309250 327922 309306 327978
rect 309374 327922 309430 327978
rect 309498 327922 309554 327978
rect 309622 327922 309678 327978
rect 309250 310294 309306 310350
rect 309374 310294 309430 310350
rect 309498 310294 309554 310350
rect 309622 310294 309678 310350
rect 309250 310170 309306 310226
rect 309374 310170 309430 310226
rect 309498 310170 309554 310226
rect 309622 310170 309678 310226
rect 309250 310046 309306 310102
rect 309374 310046 309430 310102
rect 309498 310046 309554 310102
rect 309622 310046 309678 310102
rect 309250 309922 309306 309978
rect 309374 309922 309430 309978
rect 309498 309922 309554 309978
rect 309622 309922 309678 309978
rect 309250 292294 309306 292350
rect 309374 292294 309430 292350
rect 309498 292294 309554 292350
rect 309622 292294 309678 292350
rect 309250 292170 309306 292226
rect 309374 292170 309430 292226
rect 309498 292170 309554 292226
rect 309622 292170 309678 292226
rect 309250 292046 309306 292102
rect 309374 292046 309430 292102
rect 309498 292046 309554 292102
rect 309622 292046 309678 292102
rect 309250 291922 309306 291978
rect 309374 291922 309430 291978
rect 309498 291922 309554 291978
rect 309622 291922 309678 291978
rect 309250 274294 309306 274350
rect 309374 274294 309430 274350
rect 309498 274294 309554 274350
rect 309622 274294 309678 274350
rect 309250 274170 309306 274226
rect 309374 274170 309430 274226
rect 309498 274170 309554 274226
rect 309622 274170 309678 274226
rect 309250 274046 309306 274102
rect 309374 274046 309430 274102
rect 309498 274046 309554 274102
rect 309622 274046 309678 274102
rect 309250 273922 309306 273978
rect 309374 273922 309430 273978
rect 309498 273922 309554 273978
rect 309622 273922 309678 273978
rect 309250 256294 309306 256350
rect 309374 256294 309430 256350
rect 309498 256294 309554 256350
rect 309622 256294 309678 256350
rect 309250 256170 309306 256226
rect 309374 256170 309430 256226
rect 309498 256170 309554 256226
rect 309622 256170 309678 256226
rect 309250 256046 309306 256102
rect 309374 256046 309430 256102
rect 309498 256046 309554 256102
rect 309622 256046 309678 256102
rect 309250 255922 309306 255978
rect 309374 255922 309430 255978
rect 309498 255922 309554 255978
rect 309622 255922 309678 255978
rect 291250 238294 291306 238350
rect 291374 238294 291430 238350
rect 291498 238294 291554 238350
rect 291622 238294 291678 238350
rect 291250 238170 291306 238226
rect 291374 238170 291430 238226
rect 291498 238170 291554 238226
rect 291622 238170 291678 238226
rect 291250 238046 291306 238102
rect 291374 238046 291430 238102
rect 291498 238046 291554 238102
rect 291622 238046 291678 238102
rect 291250 237922 291306 237978
rect 291374 237922 291430 237978
rect 291498 237922 291554 237978
rect 291622 237922 291678 237978
rect 291250 220294 291306 220350
rect 291374 220294 291430 220350
rect 291498 220294 291554 220350
rect 291622 220294 291678 220350
rect 291250 220170 291306 220226
rect 291374 220170 291430 220226
rect 291498 220170 291554 220226
rect 291622 220170 291678 220226
rect 291250 220046 291306 220102
rect 291374 220046 291430 220102
rect 291498 220046 291554 220102
rect 291622 220046 291678 220102
rect 291250 219922 291306 219978
rect 291374 219922 291430 219978
rect 291498 219922 291554 219978
rect 291622 219922 291678 219978
rect 291250 202294 291306 202350
rect 291374 202294 291430 202350
rect 291498 202294 291554 202350
rect 291622 202294 291678 202350
rect 291250 202170 291306 202226
rect 291374 202170 291430 202226
rect 291498 202170 291554 202226
rect 291622 202170 291678 202226
rect 291250 202046 291306 202102
rect 291374 202046 291430 202102
rect 291498 202046 291554 202102
rect 291622 202046 291678 202102
rect 291250 201922 291306 201978
rect 291374 201922 291430 201978
rect 291498 201922 291554 201978
rect 291622 201922 291678 201978
rect 291250 184294 291306 184350
rect 291374 184294 291430 184350
rect 291498 184294 291554 184350
rect 291622 184294 291678 184350
rect 291250 184170 291306 184226
rect 291374 184170 291430 184226
rect 291498 184170 291554 184226
rect 291622 184170 291678 184226
rect 291250 184046 291306 184102
rect 291374 184046 291430 184102
rect 291498 184046 291554 184102
rect 291622 184046 291678 184102
rect 291250 183922 291306 183978
rect 291374 183922 291430 183978
rect 291498 183922 291554 183978
rect 291622 183922 291678 183978
rect 284022 166356 284078 166412
rect 284146 166356 284202 166412
rect 284270 166356 284326 166412
rect 284394 166356 284450 166412
rect 284518 166356 284574 166412
rect 284642 166356 284698 166412
rect 284766 166356 284822 166412
rect 284890 166356 284946 166412
rect 285014 166356 285070 166412
rect 285138 166356 285194 166412
rect 284022 166232 284078 166288
rect 284146 166232 284202 166288
rect 284270 166232 284326 166288
rect 284394 166232 284450 166288
rect 284518 166232 284574 166288
rect 284642 166232 284698 166288
rect 284766 166232 284822 166288
rect 284890 166232 284946 166288
rect 285014 166232 285070 166288
rect 285138 166232 285194 166288
rect 284022 166108 284078 166164
rect 284146 166108 284202 166164
rect 284270 166108 284326 166164
rect 284394 166108 284450 166164
rect 284518 166108 284574 166164
rect 284642 166108 284698 166164
rect 284766 166108 284822 166164
rect 284890 166108 284946 166164
rect 285014 166108 285070 166164
rect 285138 166108 285194 166164
rect 284022 165984 284078 166040
rect 284146 165984 284202 166040
rect 284270 165984 284326 166040
rect 284394 165984 284450 166040
rect 284518 165984 284574 166040
rect 284642 165984 284698 166040
rect 284766 165984 284822 166040
rect 284890 165984 284946 166040
rect 285014 165984 285070 166040
rect 285138 165984 285194 166040
rect 284022 165860 284078 165916
rect 284146 165860 284202 165916
rect 284270 165860 284326 165916
rect 284394 165860 284450 165916
rect 284518 165860 284574 165916
rect 284642 165860 284698 165916
rect 284766 165860 284822 165916
rect 284890 165860 284946 165916
rect 285014 165860 285070 165916
rect 285138 165860 285194 165916
rect 294970 226294 295026 226350
rect 295094 226294 295150 226350
rect 295218 226294 295274 226350
rect 295342 226294 295398 226350
rect 294970 226170 295026 226226
rect 295094 226170 295150 226226
rect 295218 226170 295274 226226
rect 295342 226170 295398 226226
rect 294970 226046 295026 226102
rect 295094 226046 295150 226102
rect 295218 226046 295274 226102
rect 295342 226046 295398 226102
rect 294970 225922 295026 225978
rect 295094 225922 295150 225978
rect 295218 225922 295274 225978
rect 295342 225922 295398 225978
rect 294970 208294 295026 208350
rect 295094 208294 295150 208350
rect 295218 208294 295274 208350
rect 295342 208294 295398 208350
rect 294970 208170 295026 208226
rect 295094 208170 295150 208226
rect 295218 208170 295274 208226
rect 295342 208170 295398 208226
rect 294970 208046 295026 208102
rect 295094 208046 295150 208102
rect 295218 208046 295274 208102
rect 295342 208046 295398 208102
rect 294970 207922 295026 207978
rect 295094 207922 295150 207978
rect 295218 207922 295274 207978
rect 295342 207922 295398 207978
rect 294970 190294 295026 190350
rect 295094 190294 295150 190350
rect 295218 190294 295274 190350
rect 295342 190294 295398 190350
rect 294970 190170 295026 190226
rect 295094 190170 295150 190226
rect 295218 190170 295274 190226
rect 295342 190170 295398 190226
rect 294970 190046 295026 190102
rect 295094 190046 295150 190102
rect 295218 190046 295274 190102
rect 295342 190046 295398 190102
rect 294970 189922 295026 189978
rect 295094 189922 295150 189978
rect 295218 189922 295274 189978
rect 295342 189922 295398 189978
rect 294970 172294 295026 172350
rect 295094 172294 295150 172350
rect 295218 172294 295274 172350
rect 295342 172294 295398 172350
rect 294970 172170 295026 172226
rect 295094 172170 295150 172226
rect 295218 172170 295274 172226
rect 295342 172170 295398 172226
rect 294970 172046 295026 172102
rect 295094 172046 295150 172102
rect 295218 172046 295274 172102
rect 295342 172046 295398 172102
rect 294970 171922 295026 171978
rect 295094 171922 295150 171978
rect 295218 171922 295274 171978
rect 295342 171922 295398 171978
rect 309250 238294 309306 238350
rect 309374 238294 309430 238350
rect 309498 238294 309554 238350
rect 309622 238294 309678 238350
rect 309250 238170 309306 238226
rect 309374 238170 309430 238226
rect 309498 238170 309554 238226
rect 309622 238170 309678 238226
rect 309250 238046 309306 238102
rect 309374 238046 309430 238102
rect 309498 238046 309554 238102
rect 309622 238046 309678 238102
rect 309250 237922 309306 237978
rect 309374 237922 309430 237978
rect 309498 237922 309554 237978
rect 309622 237922 309678 237978
rect 309250 220294 309306 220350
rect 309374 220294 309430 220350
rect 309498 220294 309554 220350
rect 309622 220294 309678 220350
rect 309250 220170 309306 220226
rect 309374 220170 309430 220226
rect 309498 220170 309554 220226
rect 309622 220170 309678 220226
rect 309250 220046 309306 220102
rect 309374 220046 309430 220102
rect 309498 220046 309554 220102
rect 309622 220046 309678 220102
rect 309250 219922 309306 219978
rect 309374 219922 309430 219978
rect 309498 219922 309554 219978
rect 309622 219922 309678 219978
rect 309250 202294 309306 202350
rect 309374 202294 309430 202350
rect 309498 202294 309554 202350
rect 309622 202294 309678 202350
rect 309250 202170 309306 202226
rect 309374 202170 309430 202226
rect 309498 202170 309554 202226
rect 309622 202170 309678 202226
rect 309250 202046 309306 202102
rect 309374 202046 309430 202102
rect 309498 202046 309554 202102
rect 309622 202046 309678 202102
rect 309250 201922 309306 201978
rect 309374 201922 309430 201978
rect 309498 201922 309554 201978
rect 309622 201922 309678 201978
rect 309250 184294 309306 184350
rect 309374 184294 309430 184350
rect 309498 184294 309554 184350
rect 309622 184294 309678 184350
rect 309250 184170 309306 184226
rect 309374 184170 309430 184226
rect 309498 184170 309554 184226
rect 309622 184170 309678 184226
rect 309250 184046 309306 184102
rect 309374 184046 309430 184102
rect 309498 184046 309554 184102
rect 309622 184046 309678 184102
rect 309250 183922 309306 183978
rect 309374 183922 309430 183978
rect 309498 183922 309554 183978
rect 309622 183922 309678 183978
rect 291250 166294 291306 166350
rect 291374 166294 291430 166350
rect 291498 166294 291554 166350
rect 291622 166294 291678 166350
rect 291250 166170 291306 166226
rect 291374 166170 291430 166226
rect 291498 166170 291554 166226
rect 291622 166170 291678 166226
rect 291250 166046 291306 166102
rect 291374 166046 291430 166102
rect 291498 166046 291554 166102
rect 291622 166046 291678 166102
rect 291250 165922 291306 165978
rect 291374 165922 291430 165978
rect 291498 165922 291554 165978
rect 291622 165922 291678 165978
rect 304022 166356 304078 166412
rect 304146 166356 304202 166412
rect 304270 166356 304326 166412
rect 304394 166356 304450 166412
rect 304518 166356 304574 166412
rect 304642 166356 304698 166412
rect 304766 166356 304822 166412
rect 304890 166356 304946 166412
rect 305014 166356 305070 166412
rect 305138 166356 305194 166412
rect 304022 166232 304078 166288
rect 304146 166232 304202 166288
rect 304270 166232 304326 166288
rect 304394 166232 304450 166288
rect 304518 166232 304574 166288
rect 304642 166232 304698 166288
rect 304766 166232 304822 166288
rect 304890 166232 304946 166288
rect 305014 166232 305070 166288
rect 305138 166232 305194 166288
rect 304022 166108 304078 166164
rect 304146 166108 304202 166164
rect 304270 166108 304326 166164
rect 304394 166108 304450 166164
rect 304518 166108 304574 166164
rect 304642 166108 304698 166164
rect 304766 166108 304822 166164
rect 304890 166108 304946 166164
rect 305014 166108 305070 166164
rect 305138 166108 305194 166164
rect 304022 165984 304078 166040
rect 304146 165984 304202 166040
rect 304270 165984 304326 166040
rect 304394 165984 304450 166040
rect 304518 165984 304574 166040
rect 304642 165984 304698 166040
rect 304766 165984 304822 166040
rect 304890 165984 304946 166040
rect 305014 165984 305070 166040
rect 305138 165984 305194 166040
rect 304022 165860 304078 165916
rect 304146 165860 304202 165916
rect 304270 165860 304326 165916
rect 304394 165860 304450 165916
rect 304518 165860 304574 165916
rect 304642 165860 304698 165916
rect 304766 165860 304822 165916
rect 304890 165860 304946 165916
rect 305014 165860 305070 165916
rect 305138 165860 305194 165916
rect 309250 166294 309306 166350
rect 309374 166294 309430 166350
rect 309498 166294 309554 166350
rect 309622 166294 309678 166350
rect 309250 166170 309306 166226
rect 309374 166170 309430 166226
rect 309498 166170 309554 166226
rect 309622 166170 309678 166226
rect 309250 166046 309306 166102
rect 309374 166046 309430 166102
rect 309498 166046 309554 166102
rect 309622 166046 309678 166102
rect 309250 165922 309306 165978
rect 309374 165922 309430 165978
rect 309498 165922 309554 165978
rect 309622 165922 309678 165978
rect 312970 598116 313026 598172
rect 313094 598116 313150 598172
rect 313218 598116 313274 598172
rect 313342 598116 313398 598172
rect 312970 597992 313026 598048
rect 313094 597992 313150 598048
rect 313218 597992 313274 598048
rect 313342 597992 313398 598048
rect 312970 597868 313026 597924
rect 313094 597868 313150 597924
rect 313218 597868 313274 597924
rect 313342 597868 313398 597924
rect 312970 597744 313026 597800
rect 313094 597744 313150 597800
rect 313218 597744 313274 597800
rect 313342 597744 313398 597800
rect 312970 586294 313026 586350
rect 313094 586294 313150 586350
rect 313218 586294 313274 586350
rect 313342 586294 313398 586350
rect 312970 586170 313026 586226
rect 313094 586170 313150 586226
rect 313218 586170 313274 586226
rect 313342 586170 313398 586226
rect 312970 586046 313026 586102
rect 313094 586046 313150 586102
rect 313218 586046 313274 586102
rect 313342 586046 313398 586102
rect 312970 585922 313026 585978
rect 313094 585922 313150 585978
rect 313218 585922 313274 585978
rect 313342 585922 313398 585978
rect 312970 568294 313026 568350
rect 313094 568294 313150 568350
rect 313218 568294 313274 568350
rect 313342 568294 313398 568350
rect 312970 568170 313026 568226
rect 313094 568170 313150 568226
rect 313218 568170 313274 568226
rect 313342 568170 313398 568226
rect 312970 568046 313026 568102
rect 313094 568046 313150 568102
rect 313218 568046 313274 568102
rect 313342 568046 313398 568102
rect 312970 567922 313026 567978
rect 313094 567922 313150 567978
rect 313218 567922 313274 567978
rect 313342 567922 313398 567978
rect 312970 550294 313026 550350
rect 313094 550294 313150 550350
rect 313218 550294 313274 550350
rect 313342 550294 313398 550350
rect 312970 550170 313026 550226
rect 313094 550170 313150 550226
rect 313218 550170 313274 550226
rect 313342 550170 313398 550226
rect 312970 550046 313026 550102
rect 313094 550046 313150 550102
rect 313218 550046 313274 550102
rect 313342 550046 313398 550102
rect 312970 549922 313026 549978
rect 313094 549922 313150 549978
rect 313218 549922 313274 549978
rect 313342 549922 313398 549978
rect 312970 532294 313026 532350
rect 313094 532294 313150 532350
rect 313218 532294 313274 532350
rect 313342 532294 313398 532350
rect 312970 532170 313026 532226
rect 313094 532170 313150 532226
rect 313218 532170 313274 532226
rect 313342 532170 313398 532226
rect 312970 532046 313026 532102
rect 313094 532046 313150 532102
rect 313218 532046 313274 532102
rect 313342 532046 313398 532102
rect 312970 531922 313026 531978
rect 313094 531922 313150 531978
rect 313218 531922 313274 531978
rect 313342 531922 313398 531978
rect 312970 514294 313026 514350
rect 313094 514294 313150 514350
rect 313218 514294 313274 514350
rect 313342 514294 313398 514350
rect 312970 514170 313026 514226
rect 313094 514170 313150 514226
rect 313218 514170 313274 514226
rect 313342 514170 313398 514226
rect 312970 514046 313026 514102
rect 313094 514046 313150 514102
rect 313218 514046 313274 514102
rect 313342 514046 313398 514102
rect 312970 513922 313026 513978
rect 313094 513922 313150 513978
rect 313218 513922 313274 513978
rect 313342 513922 313398 513978
rect 312970 496294 313026 496350
rect 313094 496294 313150 496350
rect 313218 496294 313274 496350
rect 313342 496294 313398 496350
rect 312970 496170 313026 496226
rect 313094 496170 313150 496226
rect 313218 496170 313274 496226
rect 313342 496170 313398 496226
rect 312970 496046 313026 496102
rect 313094 496046 313150 496102
rect 313218 496046 313274 496102
rect 313342 496046 313398 496102
rect 312970 495922 313026 495978
rect 313094 495922 313150 495978
rect 313218 495922 313274 495978
rect 313342 495922 313398 495978
rect 312970 478294 313026 478350
rect 313094 478294 313150 478350
rect 313218 478294 313274 478350
rect 313342 478294 313398 478350
rect 312970 478170 313026 478226
rect 313094 478170 313150 478226
rect 313218 478170 313274 478226
rect 313342 478170 313398 478226
rect 312970 478046 313026 478102
rect 313094 478046 313150 478102
rect 313218 478046 313274 478102
rect 313342 478046 313398 478102
rect 312970 477922 313026 477978
rect 313094 477922 313150 477978
rect 313218 477922 313274 477978
rect 313342 477922 313398 477978
rect 312970 460294 313026 460350
rect 313094 460294 313150 460350
rect 313218 460294 313274 460350
rect 313342 460294 313398 460350
rect 312970 460170 313026 460226
rect 313094 460170 313150 460226
rect 313218 460170 313274 460226
rect 313342 460170 313398 460226
rect 312970 460046 313026 460102
rect 313094 460046 313150 460102
rect 313218 460046 313274 460102
rect 313342 460046 313398 460102
rect 312970 459922 313026 459978
rect 313094 459922 313150 459978
rect 313218 459922 313274 459978
rect 313342 459922 313398 459978
rect 312970 442294 313026 442350
rect 313094 442294 313150 442350
rect 313218 442294 313274 442350
rect 313342 442294 313398 442350
rect 312970 442170 313026 442226
rect 313094 442170 313150 442226
rect 313218 442170 313274 442226
rect 313342 442170 313398 442226
rect 312970 442046 313026 442102
rect 313094 442046 313150 442102
rect 313218 442046 313274 442102
rect 313342 442046 313398 442102
rect 312970 441922 313026 441978
rect 313094 441922 313150 441978
rect 313218 441922 313274 441978
rect 313342 441922 313398 441978
rect 312970 424294 313026 424350
rect 313094 424294 313150 424350
rect 313218 424294 313274 424350
rect 313342 424294 313398 424350
rect 312970 424170 313026 424226
rect 313094 424170 313150 424226
rect 313218 424170 313274 424226
rect 313342 424170 313398 424226
rect 312970 424046 313026 424102
rect 313094 424046 313150 424102
rect 313218 424046 313274 424102
rect 313342 424046 313398 424102
rect 312970 423922 313026 423978
rect 313094 423922 313150 423978
rect 313218 423922 313274 423978
rect 313342 423922 313398 423978
rect 312970 406294 313026 406350
rect 313094 406294 313150 406350
rect 313218 406294 313274 406350
rect 313342 406294 313398 406350
rect 312970 406170 313026 406226
rect 313094 406170 313150 406226
rect 313218 406170 313274 406226
rect 313342 406170 313398 406226
rect 312970 406046 313026 406102
rect 313094 406046 313150 406102
rect 313218 406046 313274 406102
rect 313342 406046 313398 406102
rect 312970 405922 313026 405978
rect 313094 405922 313150 405978
rect 313218 405922 313274 405978
rect 313342 405922 313398 405978
rect 312970 388294 313026 388350
rect 313094 388294 313150 388350
rect 313218 388294 313274 388350
rect 313342 388294 313398 388350
rect 312970 388170 313026 388226
rect 313094 388170 313150 388226
rect 313218 388170 313274 388226
rect 313342 388170 313398 388226
rect 312970 388046 313026 388102
rect 313094 388046 313150 388102
rect 313218 388046 313274 388102
rect 313342 388046 313398 388102
rect 312970 387922 313026 387978
rect 313094 387922 313150 387978
rect 313218 387922 313274 387978
rect 313342 387922 313398 387978
rect 312970 370294 313026 370350
rect 313094 370294 313150 370350
rect 313218 370294 313274 370350
rect 313342 370294 313398 370350
rect 312970 370170 313026 370226
rect 313094 370170 313150 370226
rect 313218 370170 313274 370226
rect 313342 370170 313398 370226
rect 312970 370046 313026 370102
rect 313094 370046 313150 370102
rect 313218 370046 313274 370102
rect 313342 370046 313398 370102
rect 312970 369922 313026 369978
rect 313094 369922 313150 369978
rect 313218 369922 313274 369978
rect 313342 369922 313398 369978
rect 312970 352294 313026 352350
rect 313094 352294 313150 352350
rect 313218 352294 313274 352350
rect 313342 352294 313398 352350
rect 312970 352170 313026 352226
rect 313094 352170 313150 352226
rect 313218 352170 313274 352226
rect 313342 352170 313398 352226
rect 312970 352046 313026 352102
rect 313094 352046 313150 352102
rect 313218 352046 313274 352102
rect 313342 352046 313398 352102
rect 312970 351922 313026 351978
rect 313094 351922 313150 351978
rect 313218 351922 313274 351978
rect 313342 351922 313398 351978
rect 312970 334294 313026 334350
rect 313094 334294 313150 334350
rect 313218 334294 313274 334350
rect 313342 334294 313398 334350
rect 312970 334170 313026 334226
rect 313094 334170 313150 334226
rect 313218 334170 313274 334226
rect 313342 334170 313398 334226
rect 312970 334046 313026 334102
rect 313094 334046 313150 334102
rect 313218 334046 313274 334102
rect 313342 334046 313398 334102
rect 312970 333922 313026 333978
rect 313094 333922 313150 333978
rect 313218 333922 313274 333978
rect 313342 333922 313398 333978
rect 312970 316294 313026 316350
rect 313094 316294 313150 316350
rect 313218 316294 313274 316350
rect 313342 316294 313398 316350
rect 312970 316170 313026 316226
rect 313094 316170 313150 316226
rect 313218 316170 313274 316226
rect 313342 316170 313398 316226
rect 312970 316046 313026 316102
rect 313094 316046 313150 316102
rect 313218 316046 313274 316102
rect 313342 316046 313398 316102
rect 312970 315922 313026 315978
rect 313094 315922 313150 315978
rect 313218 315922 313274 315978
rect 313342 315922 313398 315978
rect 312970 298294 313026 298350
rect 313094 298294 313150 298350
rect 313218 298294 313274 298350
rect 313342 298294 313398 298350
rect 312970 298170 313026 298226
rect 313094 298170 313150 298226
rect 313218 298170 313274 298226
rect 313342 298170 313398 298226
rect 312970 298046 313026 298102
rect 313094 298046 313150 298102
rect 313218 298046 313274 298102
rect 313342 298046 313398 298102
rect 312970 297922 313026 297978
rect 313094 297922 313150 297978
rect 313218 297922 313274 297978
rect 313342 297922 313398 297978
rect 312970 280294 313026 280350
rect 313094 280294 313150 280350
rect 313218 280294 313274 280350
rect 313342 280294 313398 280350
rect 312970 280170 313026 280226
rect 313094 280170 313150 280226
rect 313218 280170 313274 280226
rect 313342 280170 313398 280226
rect 312970 280046 313026 280102
rect 313094 280046 313150 280102
rect 313218 280046 313274 280102
rect 313342 280046 313398 280102
rect 312970 279922 313026 279978
rect 313094 279922 313150 279978
rect 313218 279922 313274 279978
rect 313342 279922 313398 279978
rect 312970 262294 313026 262350
rect 313094 262294 313150 262350
rect 313218 262294 313274 262350
rect 313342 262294 313398 262350
rect 312970 262170 313026 262226
rect 313094 262170 313150 262226
rect 313218 262170 313274 262226
rect 313342 262170 313398 262226
rect 312970 262046 313026 262102
rect 313094 262046 313150 262102
rect 313218 262046 313274 262102
rect 313342 262046 313398 262102
rect 312970 261922 313026 261978
rect 313094 261922 313150 261978
rect 313218 261922 313274 261978
rect 313342 261922 313398 261978
rect 312970 244294 313026 244350
rect 313094 244294 313150 244350
rect 313218 244294 313274 244350
rect 313342 244294 313398 244350
rect 312970 244170 313026 244226
rect 313094 244170 313150 244226
rect 313218 244170 313274 244226
rect 313342 244170 313398 244226
rect 312970 244046 313026 244102
rect 313094 244046 313150 244102
rect 313218 244046 313274 244102
rect 313342 244046 313398 244102
rect 312970 243922 313026 243978
rect 313094 243922 313150 243978
rect 313218 243922 313274 243978
rect 313342 243922 313398 243978
rect 312970 226294 313026 226350
rect 313094 226294 313150 226350
rect 313218 226294 313274 226350
rect 313342 226294 313398 226350
rect 312970 226170 313026 226226
rect 313094 226170 313150 226226
rect 313218 226170 313274 226226
rect 313342 226170 313398 226226
rect 312970 226046 313026 226102
rect 313094 226046 313150 226102
rect 313218 226046 313274 226102
rect 313342 226046 313398 226102
rect 312970 225922 313026 225978
rect 313094 225922 313150 225978
rect 313218 225922 313274 225978
rect 313342 225922 313398 225978
rect 312970 208294 313026 208350
rect 313094 208294 313150 208350
rect 313218 208294 313274 208350
rect 313342 208294 313398 208350
rect 312970 208170 313026 208226
rect 313094 208170 313150 208226
rect 313218 208170 313274 208226
rect 313342 208170 313398 208226
rect 312970 208046 313026 208102
rect 313094 208046 313150 208102
rect 313218 208046 313274 208102
rect 313342 208046 313398 208102
rect 312970 207922 313026 207978
rect 313094 207922 313150 207978
rect 313218 207922 313274 207978
rect 313342 207922 313398 207978
rect 312970 190294 313026 190350
rect 313094 190294 313150 190350
rect 313218 190294 313274 190350
rect 313342 190294 313398 190350
rect 312970 190170 313026 190226
rect 313094 190170 313150 190226
rect 313218 190170 313274 190226
rect 313342 190170 313398 190226
rect 312970 190046 313026 190102
rect 313094 190046 313150 190102
rect 313218 190046 313274 190102
rect 313342 190046 313398 190102
rect 312970 189922 313026 189978
rect 313094 189922 313150 189978
rect 313218 189922 313274 189978
rect 313342 189922 313398 189978
rect 312970 172294 313026 172350
rect 313094 172294 313150 172350
rect 313218 172294 313274 172350
rect 313342 172294 313398 172350
rect 312970 172170 313026 172226
rect 313094 172170 313150 172226
rect 313218 172170 313274 172226
rect 313342 172170 313398 172226
rect 312970 172046 313026 172102
rect 313094 172046 313150 172102
rect 313218 172046 313274 172102
rect 313342 172046 313398 172102
rect 312970 171922 313026 171978
rect 313094 171922 313150 171978
rect 313218 171922 313274 171978
rect 313342 171922 313398 171978
rect 327250 597156 327306 597212
rect 327374 597156 327430 597212
rect 327498 597156 327554 597212
rect 327622 597156 327678 597212
rect 327250 597032 327306 597088
rect 327374 597032 327430 597088
rect 327498 597032 327554 597088
rect 327622 597032 327678 597088
rect 327250 596908 327306 596964
rect 327374 596908 327430 596964
rect 327498 596908 327554 596964
rect 327622 596908 327678 596964
rect 327250 596784 327306 596840
rect 327374 596784 327430 596840
rect 327498 596784 327554 596840
rect 327622 596784 327678 596840
rect 327250 580294 327306 580350
rect 327374 580294 327430 580350
rect 327498 580294 327554 580350
rect 327622 580294 327678 580350
rect 327250 580170 327306 580226
rect 327374 580170 327430 580226
rect 327498 580170 327554 580226
rect 327622 580170 327678 580226
rect 327250 580046 327306 580102
rect 327374 580046 327430 580102
rect 327498 580046 327554 580102
rect 327622 580046 327678 580102
rect 327250 579922 327306 579978
rect 327374 579922 327430 579978
rect 327498 579922 327554 579978
rect 327622 579922 327678 579978
rect 327250 562294 327306 562350
rect 327374 562294 327430 562350
rect 327498 562294 327554 562350
rect 327622 562294 327678 562350
rect 327250 562170 327306 562226
rect 327374 562170 327430 562226
rect 327498 562170 327554 562226
rect 327622 562170 327678 562226
rect 327250 562046 327306 562102
rect 327374 562046 327430 562102
rect 327498 562046 327554 562102
rect 327622 562046 327678 562102
rect 327250 561922 327306 561978
rect 327374 561922 327430 561978
rect 327498 561922 327554 561978
rect 327622 561922 327678 561978
rect 327250 544294 327306 544350
rect 327374 544294 327430 544350
rect 327498 544294 327554 544350
rect 327622 544294 327678 544350
rect 327250 544170 327306 544226
rect 327374 544170 327430 544226
rect 327498 544170 327554 544226
rect 327622 544170 327678 544226
rect 327250 544046 327306 544102
rect 327374 544046 327430 544102
rect 327498 544046 327554 544102
rect 327622 544046 327678 544102
rect 327250 543922 327306 543978
rect 327374 543922 327430 543978
rect 327498 543922 327554 543978
rect 327622 543922 327678 543978
rect 327250 526294 327306 526350
rect 327374 526294 327430 526350
rect 327498 526294 327554 526350
rect 327622 526294 327678 526350
rect 327250 526170 327306 526226
rect 327374 526170 327430 526226
rect 327498 526170 327554 526226
rect 327622 526170 327678 526226
rect 327250 526046 327306 526102
rect 327374 526046 327430 526102
rect 327498 526046 327554 526102
rect 327622 526046 327678 526102
rect 327250 525922 327306 525978
rect 327374 525922 327430 525978
rect 327498 525922 327554 525978
rect 327622 525922 327678 525978
rect 327250 508294 327306 508350
rect 327374 508294 327430 508350
rect 327498 508294 327554 508350
rect 327622 508294 327678 508350
rect 327250 508170 327306 508226
rect 327374 508170 327430 508226
rect 327498 508170 327554 508226
rect 327622 508170 327678 508226
rect 327250 508046 327306 508102
rect 327374 508046 327430 508102
rect 327498 508046 327554 508102
rect 327622 508046 327678 508102
rect 327250 507922 327306 507978
rect 327374 507922 327430 507978
rect 327498 507922 327554 507978
rect 327622 507922 327678 507978
rect 327250 490294 327306 490350
rect 327374 490294 327430 490350
rect 327498 490294 327554 490350
rect 327622 490294 327678 490350
rect 327250 490170 327306 490226
rect 327374 490170 327430 490226
rect 327498 490170 327554 490226
rect 327622 490170 327678 490226
rect 327250 490046 327306 490102
rect 327374 490046 327430 490102
rect 327498 490046 327554 490102
rect 327622 490046 327678 490102
rect 327250 489922 327306 489978
rect 327374 489922 327430 489978
rect 327498 489922 327554 489978
rect 327622 489922 327678 489978
rect 327250 472294 327306 472350
rect 327374 472294 327430 472350
rect 327498 472294 327554 472350
rect 327622 472294 327678 472350
rect 327250 472170 327306 472226
rect 327374 472170 327430 472226
rect 327498 472170 327554 472226
rect 327622 472170 327678 472226
rect 327250 472046 327306 472102
rect 327374 472046 327430 472102
rect 327498 472046 327554 472102
rect 327622 472046 327678 472102
rect 327250 471922 327306 471978
rect 327374 471922 327430 471978
rect 327498 471922 327554 471978
rect 327622 471922 327678 471978
rect 327250 454294 327306 454350
rect 327374 454294 327430 454350
rect 327498 454294 327554 454350
rect 327622 454294 327678 454350
rect 327250 454170 327306 454226
rect 327374 454170 327430 454226
rect 327498 454170 327554 454226
rect 327622 454170 327678 454226
rect 327250 454046 327306 454102
rect 327374 454046 327430 454102
rect 327498 454046 327554 454102
rect 327622 454046 327678 454102
rect 327250 453922 327306 453978
rect 327374 453922 327430 453978
rect 327498 453922 327554 453978
rect 327622 453922 327678 453978
rect 327250 436294 327306 436350
rect 327374 436294 327430 436350
rect 327498 436294 327554 436350
rect 327622 436294 327678 436350
rect 327250 436170 327306 436226
rect 327374 436170 327430 436226
rect 327498 436170 327554 436226
rect 327622 436170 327678 436226
rect 327250 436046 327306 436102
rect 327374 436046 327430 436102
rect 327498 436046 327554 436102
rect 327622 436046 327678 436102
rect 327250 435922 327306 435978
rect 327374 435922 327430 435978
rect 327498 435922 327554 435978
rect 327622 435922 327678 435978
rect 327250 418294 327306 418350
rect 327374 418294 327430 418350
rect 327498 418294 327554 418350
rect 327622 418294 327678 418350
rect 327250 418170 327306 418226
rect 327374 418170 327430 418226
rect 327498 418170 327554 418226
rect 327622 418170 327678 418226
rect 327250 418046 327306 418102
rect 327374 418046 327430 418102
rect 327498 418046 327554 418102
rect 327622 418046 327678 418102
rect 327250 417922 327306 417978
rect 327374 417922 327430 417978
rect 327498 417922 327554 417978
rect 327622 417922 327678 417978
rect 327250 400294 327306 400350
rect 327374 400294 327430 400350
rect 327498 400294 327554 400350
rect 327622 400294 327678 400350
rect 327250 400170 327306 400226
rect 327374 400170 327430 400226
rect 327498 400170 327554 400226
rect 327622 400170 327678 400226
rect 327250 400046 327306 400102
rect 327374 400046 327430 400102
rect 327498 400046 327554 400102
rect 327622 400046 327678 400102
rect 327250 399922 327306 399978
rect 327374 399922 327430 399978
rect 327498 399922 327554 399978
rect 327622 399922 327678 399978
rect 327250 382294 327306 382350
rect 327374 382294 327430 382350
rect 327498 382294 327554 382350
rect 327622 382294 327678 382350
rect 327250 382170 327306 382226
rect 327374 382170 327430 382226
rect 327498 382170 327554 382226
rect 327622 382170 327678 382226
rect 327250 382046 327306 382102
rect 327374 382046 327430 382102
rect 327498 382046 327554 382102
rect 327622 382046 327678 382102
rect 327250 381922 327306 381978
rect 327374 381922 327430 381978
rect 327498 381922 327554 381978
rect 327622 381922 327678 381978
rect 327250 364294 327306 364350
rect 327374 364294 327430 364350
rect 327498 364294 327554 364350
rect 327622 364294 327678 364350
rect 327250 364170 327306 364226
rect 327374 364170 327430 364226
rect 327498 364170 327554 364226
rect 327622 364170 327678 364226
rect 327250 364046 327306 364102
rect 327374 364046 327430 364102
rect 327498 364046 327554 364102
rect 327622 364046 327678 364102
rect 327250 363922 327306 363978
rect 327374 363922 327430 363978
rect 327498 363922 327554 363978
rect 327622 363922 327678 363978
rect 327250 346294 327306 346350
rect 327374 346294 327430 346350
rect 327498 346294 327554 346350
rect 327622 346294 327678 346350
rect 327250 346170 327306 346226
rect 327374 346170 327430 346226
rect 327498 346170 327554 346226
rect 327622 346170 327678 346226
rect 327250 346046 327306 346102
rect 327374 346046 327430 346102
rect 327498 346046 327554 346102
rect 327622 346046 327678 346102
rect 327250 345922 327306 345978
rect 327374 345922 327430 345978
rect 327498 345922 327554 345978
rect 327622 345922 327678 345978
rect 327250 328294 327306 328350
rect 327374 328294 327430 328350
rect 327498 328294 327554 328350
rect 327622 328294 327678 328350
rect 327250 328170 327306 328226
rect 327374 328170 327430 328226
rect 327498 328170 327554 328226
rect 327622 328170 327678 328226
rect 327250 328046 327306 328102
rect 327374 328046 327430 328102
rect 327498 328046 327554 328102
rect 327622 328046 327678 328102
rect 327250 327922 327306 327978
rect 327374 327922 327430 327978
rect 327498 327922 327554 327978
rect 327622 327922 327678 327978
rect 327250 310294 327306 310350
rect 327374 310294 327430 310350
rect 327498 310294 327554 310350
rect 327622 310294 327678 310350
rect 327250 310170 327306 310226
rect 327374 310170 327430 310226
rect 327498 310170 327554 310226
rect 327622 310170 327678 310226
rect 327250 310046 327306 310102
rect 327374 310046 327430 310102
rect 327498 310046 327554 310102
rect 327622 310046 327678 310102
rect 327250 309922 327306 309978
rect 327374 309922 327430 309978
rect 327498 309922 327554 309978
rect 327622 309922 327678 309978
rect 327250 292294 327306 292350
rect 327374 292294 327430 292350
rect 327498 292294 327554 292350
rect 327622 292294 327678 292350
rect 327250 292170 327306 292226
rect 327374 292170 327430 292226
rect 327498 292170 327554 292226
rect 327622 292170 327678 292226
rect 327250 292046 327306 292102
rect 327374 292046 327430 292102
rect 327498 292046 327554 292102
rect 327622 292046 327678 292102
rect 327250 291922 327306 291978
rect 327374 291922 327430 291978
rect 327498 291922 327554 291978
rect 327622 291922 327678 291978
rect 327250 274294 327306 274350
rect 327374 274294 327430 274350
rect 327498 274294 327554 274350
rect 327622 274294 327678 274350
rect 327250 274170 327306 274226
rect 327374 274170 327430 274226
rect 327498 274170 327554 274226
rect 327622 274170 327678 274226
rect 327250 274046 327306 274102
rect 327374 274046 327430 274102
rect 327498 274046 327554 274102
rect 327622 274046 327678 274102
rect 327250 273922 327306 273978
rect 327374 273922 327430 273978
rect 327498 273922 327554 273978
rect 327622 273922 327678 273978
rect 327250 256294 327306 256350
rect 327374 256294 327430 256350
rect 327498 256294 327554 256350
rect 327622 256294 327678 256350
rect 327250 256170 327306 256226
rect 327374 256170 327430 256226
rect 327498 256170 327554 256226
rect 327622 256170 327678 256226
rect 327250 256046 327306 256102
rect 327374 256046 327430 256102
rect 327498 256046 327554 256102
rect 327622 256046 327678 256102
rect 327250 255922 327306 255978
rect 327374 255922 327430 255978
rect 327498 255922 327554 255978
rect 327622 255922 327678 255978
rect 327250 238294 327306 238350
rect 327374 238294 327430 238350
rect 327498 238294 327554 238350
rect 327622 238294 327678 238350
rect 327250 238170 327306 238226
rect 327374 238170 327430 238226
rect 327498 238170 327554 238226
rect 327622 238170 327678 238226
rect 327250 238046 327306 238102
rect 327374 238046 327430 238102
rect 327498 238046 327554 238102
rect 327622 238046 327678 238102
rect 327250 237922 327306 237978
rect 327374 237922 327430 237978
rect 327498 237922 327554 237978
rect 327622 237922 327678 237978
rect 327250 220294 327306 220350
rect 327374 220294 327430 220350
rect 327498 220294 327554 220350
rect 327622 220294 327678 220350
rect 327250 220170 327306 220226
rect 327374 220170 327430 220226
rect 327498 220170 327554 220226
rect 327622 220170 327678 220226
rect 327250 220046 327306 220102
rect 327374 220046 327430 220102
rect 327498 220046 327554 220102
rect 327622 220046 327678 220102
rect 327250 219922 327306 219978
rect 327374 219922 327430 219978
rect 327498 219922 327554 219978
rect 327622 219922 327678 219978
rect 327250 202294 327306 202350
rect 327374 202294 327430 202350
rect 327498 202294 327554 202350
rect 327622 202294 327678 202350
rect 327250 202170 327306 202226
rect 327374 202170 327430 202226
rect 327498 202170 327554 202226
rect 327622 202170 327678 202226
rect 327250 202046 327306 202102
rect 327374 202046 327430 202102
rect 327498 202046 327554 202102
rect 327622 202046 327678 202102
rect 327250 201922 327306 201978
rect 327374 201922 327430 201978
rect 327498 201922 327554 201978
rect 327622 201922 327678 201978
rect 327250 184294 327306 184350
rect 327374 184294 327430 184350
rect 327498 184294 327554 184350
rect 327622 184294 327678 184350
rect 327250 184170 327306 184226
rect 327374 184170 327430 184226
rect 327498 184170 327554 184226
rect 327622 184170 327678 184226
rect 327250 184046 327306 184102
rect 327374 184046 327430 184102
rect 327498 184046 327554 184102
rect 327622 184046 327678 184102
rect 327250 183922 327306 183978
rect 327374 183922 327430 183978
rect 327498 183922 327554 183978
rect 327622 183922 327678 183978
rect 327250 166294 327306 166350
rect 327374 166294 327430 166350
rect 327498 166294 327554 166350
rect 327622 166294 327678 166350
rect 327250 166170 327306 166226
rect 327374 166170 327430 166226
rect 327498 166170 327554 166226
rect 327622 166170 327678 166226
rect 327250 166046 327306 166102
rect 327374 166046 327430 166102
rect 327498 166046 327554 166102
rect 327622 166046 327678 166102
rect 327250 165922 327306 165978
rect 327374 165922 327430 165978
rect 327498 165922 327554 165978
rect 327622 165922 327678 165978
rect 276970 154294 277026 154350
rect 277094 154294 277150 154350
rect 277218 154294 277274 154350
rect 277342 154294 277398 154350
rect 276970 154170 277026 154226
rect 277094 154170 277150 154226
rect 277218 154170 277274 154226
rect 277342 154170 277398 154226
rect 276970 154046 277026 154102
rect 277094 154046 277150 154102
rect 277218 154046 277274 154102
rect 277342 154046 277398 154102
rect 276970 153922 277026 153978
rect 277094 153922 277150 153978
rect 277218 153922 277274 153978
rect 277342 153922 277398 153978
rect 294022 154356 294078 154412
rect 294146 154356 294202 154412
rect 294270 154356 294326 154412
rect 294394 154356 294450 154412
rect 294518 154356 294574 154412
rect 294642 154356 294698 154412
rect 294766 154356 294822 154412
rect 294890 154356 294946 154412
rect 295014 154356 295070 154412
rect 295138 154356 295194 154412
rect 294022 154232 294078 154288
rect 294146 154232 294202 154288
rect 294270 154232 294326 154288
rect 294394 154232 294450 154288
rect 294518 154232 294574 154288
rect 294642 154232 294698 154288
rect 294766 154232 294822 154288
rect 294890 154232 294946 154288
rect 295014 154232 295070 154288
rect 295138 154232 295194 154288
rect 294022 154108 294078 154164
rect 294146 154108 294202 154164
rect 294270 154108 294326 154164
rect 294394 154108 294450 154164
rect 294518 154108 294574 154164
rect 294642 154108 294698 154164
rect 294766 154108 294822 154164
rect 294890 154108 294946 154164
rect 295014 154108 295070 154164
rect 295138 154108 295194 154164
rect 294022 153984 294078 154040
rect 294146 153984 294202 154040
rect 294270 153984 294326 154040
rect 294394 153984 294450 154040
rect 294518 153984 294574 154040
rect 294642 153984 294698 154040
rect 294766 153984 294822 154040
rect 294890 153984 294946 154040
rect 295014 153984 295070 154040
rect 295138 153984 295194 154040
rect 294022 153860 294078 153916
rect 294146 153860 294202 153916
rect 294270 153860 294326 153916
rect 294394 153860 294450 153916
rect 294518 153860 294574 153916
rect 294642 153860 294698 153916
rect 294766 153860 294822 153916
rect 294890 153860 294946 153916
rect 295014 153860 295070 153916
rect 295138 153860 295194 153916
rect 314022 154356 314078 154412
rect 314146 154356 314202 154412
rect 314270 154356 314326 154412
rect 314394 154356 314450 154412
rect 314518 154356 314574 154412
rect 314642 154356 314698 154412
rect 314766 154356 314822 154412
rect 314890 154356 314946 154412
rect 315014 154356 315070 154412
rect 315138 154356 315194 154412
rect 314022 154232 314078 154288
rect 314146 154232 314202 154288
rect 314270 154232 314326 154288
rect 314394 154232 314450 154288
rect 314518 154232 314574 154288
rect 314642 154232 314698 154288
rect 314766 154232 314822 154288
rect 314890 154232 314946 154288
rect 315014 154232 315070 154288
rect 315138 154232 315194 154288
rect 314022 154108 314078 154164
rect 314146 154108 314202 154164
rect 314270 154108 314326 154164
rect 314394 154108 314450 154164
rect 314518 154108 314574 154164
rect 314642 154108 314698 154164
rect 314766 154108 314822 154164
rect 314890 154108 314946 154164
rect 315014 154108 315070 154164
rect 315138 154108 315194 154164
rect 314022 153984 314078 154040
rect 314146 153984 314202 154040
rect 314270 153984 314326 154040
rect 314394 153984 314450 154040
rect 314518 153984 314574 154040
rect 314642 153984 314698 154040
rect 314766 153984 314822 154040
rect 314890 153984 314946 154040
rect 315014 153984 315070 154040
rect 315138 153984 315194 154040
rect 314022 153860 314078 153916
rect 314146 153860 314202 153916
rect 314270 153860 314326 153916
rect 314394 153860 314450 153916
rect 314518 153860 314574 153916
rect 314642 153860 314698 153916
rect 314766 153860 314822 153916
rect 314890 153860 314946 153916
rect 315014 153860 315070 153916
rect 315138 153860 315194 153916
rect 284022 148356 284078 148412
rect 284146 148356 284202 148412
rect 284270 148356 284326 148412
rect 284394 148356 284450 148412
rect 284518 148356 284574 148412
rect 284642 148356 284698 148412
rect 284766 148356 284822 148412
rect 284890 148356 284946 148412
rect 285014 148356 285070 148412
rect 285138 148356 285194 148412
rect 284022 148232 284078 148288
rect 284146 148232 284202 148288
rect 284270 148232 284326 148288
rect 284394 148232 284450 148288
rect 284518 148232 284574 148288
rect 284642 148232 284698 148288
rect 284766 148232 284822 148288
rect 284890 148232 284946 148288
rect 285014 148232 285070 148288
rect 285138 148232 285194 148288
rect 284022 148108 284078 148164
rect 284146 148108 284202 148164
rect 284270 148108 284326 148164
rect 284394 148108 284450 148164
rect 284518 148108 284574 148164
rect 284642 148108 284698 148164
rect 284766 148108 284822 148164
rect 284890 148108 284946 148164
rect 285014 148108 285070 148164
rect 285138 148108 285194 148164
rect 284022 147984 284078 148040
rect 284146 147984 284202 148040
rect 284270 147984 284326 148040
rect 284394 147984 284450 148040
rect 284518 147984 284574 148040
rect 284642 147984 284698 148040
rect 284766 147984 284822 148040
rect 284890 147984 284946 148040
rect 285014 147984 285070 148040
rect 285138 147984 285194 148040
rect 284022 147860 284078 147916
rect 284146 147860 284202 147916
rect 284270 147860 284326 147916
rect 284394 147860 284450 147916
rect 284518 147860 284574 147916
rect 284642 147860 284698 147916
rect 284766 147860 284822 147916
rect 284890 147860 284946 147916
rect 285014 147860 285070 147916
rect 285138 147860 285194 147916
rect 304022 148356 304078 148412
rect 304146 148356 304202 148412
rect 304270 148356 304326 148412
rect 304394 148356 304450 148412
rect 304518 148356 304574 148412
rect 304642 148356 304698 148412
rect 304766 148356 304822 148412
rect 304890 148356 304946 148412
rect 305014 148356 305070 148412
rect 305138 148356 305194 148412
rect 304022 148232 304078 148288
rect 304146 148232 304202 148288
rect 304270 148232 304326 148288
rect 304394 148232 304450 148288
rect 304518 148232 304574 148288
rect 304642 148232 304698 148288
rect 304766 148232 304822 148288
rect 304890 148232 304946 148288
rect 305014 148232 305070 148288
rect 305138 148232 305194 148288
rect 304022 148108 304078 148164
rect 304146 148108 304202 148164
rect 304270 148108 304326 148164
rect 304394 148108 304450 148164
rect 304518 148108 304574 148164
rect 304642 148108 304698 148164
rect 304766 148108 304822 148164
rect 304890 148108 304946 148164
rect 305014 148108 305070 148164
rect 305138 148108 305194 148164
rect 304022 147984 304078 148040
rect 304146 147984 304202 148040
rect 304270 147984 304326 148040
rect 304394 147984 304450 148040
rect 304518 147984 304574 148040
rect 304642 147984 304698 148040
rect 304766 147984 304822 148040
rect 304890 147984 304946 148040
rect 305014 147984 305070 148040
rect 305138 147984 305194 148040
rect 304022 147860 304078 147916
rect 304146 147860 304202 147916
rect 304270 147860 304326 147916
rect 304394 147860 304450 147916
rect 304518 147860 304574 147916
rect 304642 147860 304698 147916
rect 304766 147860 304822 147916
rect 304890 147860 304946 147916
rect 305014 147860 305070 147916
rect 305138 147860 305194 147916
rect 327250 148294 327306 148350
rect 327374 148294 327430 148350
rect 327498 148294 327554 148350
rect 327622 148294 327678 148350
rect 327250 148170 327306 148226
rect 327374 148170 327430 148226
rect 327498 148170 327554 148226
rect 327622 148170 327678 148226
rect 327250 148046 327306 148102
rect 327374 148046 327430 148102
rect 327498 148046 327554 148102
rect 327622 148046 327678 148102
rect 327250 147922 327306 147978
rect 327374 147922 327430 147978
rect 327498 147922 327554 147978
rect 327622 147922 327678 147978
rect 276970 136294 277026 136350
rect 277094 136294 277150 136350
rect 277218 136294 277274 136350
rect 277342 136294 277398 136350
rect 276970 136170 277026 136226
rect 277094 136170 277150 136226
rect 277218 136170 277274 136226
rect 277342 136170 277398 136226
rect 276970 136046 277026 136102
rect 277094 136046 277150 136102
rect 277218 136046 277274 136102
rect 277342 136046 277398 136102
rect 276970 135922 277026 135978
rect 277094 135922 277150 135978
rect 277218 135922 277274 135978
rect 277342 135922 277398 135978
rect 294022 136356 294078 136412
rect 294146 136356 294202 136412
rect 294270 136356 294326 136412
rect 294394 136356 294450 136412
rect 294518 136356 294574 136412
rect 294642 136356 294698 136412
rect 294766 136356 294822 136412
rect 294890 136356 294946 136412
rect 295014 136356 295070 136412
rect 295138 136356 295194 136412
rect 294022 136232 294078 136288
rect 294146 136232 294202 136288
rect 294270 136232 294326 136288
rect 294394 136232 294450 136288
rect 294518 136232 294574 136288
rect 294642 136232 294698 136288
rect 294766 136232 294822 136288
rect 294890 136232 294946 136288
rect 295014 136232 295070 136288
rect 295138 136232 295194 136288
rect 294022 136108 294078 136164
rect 294146 136108 294202 136164
rect 294270 136108 294326 136164
rect 294394 136108 294450 136164
rect 294518 136108 294574 136164
rect 294642 136108 294698 136164
rect 294766 136108 294822 136164
rect 294890 136108 294946 136164
rect 295014 136108 295070 136164
rect 295138 136108 295194 136164
rect 294022 135984 294078 136040
rect 294146 135984 294202 136040
rect 294270 135984 294326 136040
rect 294394 135984 294450 136040
rect 294518 135984 294574 136040
rect 294642 135984 294698 136040
rect 294766 135984 294822 136040
rect 294890 135984 294946 136040
rect 295014 135984 295070 136040
rect 295138 135984 295194 136040
rect 294022 135860 294078 135916
rect 294146 135860 294202 135916
rect 294270 135860 294326 135916
rect 294394 135860 294450 135916
rect 294518 135860 294574 135916
rect 294642 135860 294698 135916
rect 294766 135860 294822 135916
rect 294890 135860 294946 135916
rect 295014 135860 295070 135916
rect 295138 135860 295194 135916
rect 314022 136356 314078 136412
rect 314146 136356 314202 136412
rect 314270 136356 314326 136412
rect 314394 136356 314450 136412
rect 314518 136356 314574 136412
rect 314642 136356 314698 136412
rect 314766 136356 314822 136412
rect 314890 136356 314946 136412
rect 315014 136356 315070 136412
rect 315138 136356 315194 136412
rect 314022 136232 314078 136288
rect 314146 136232 314202 136288
rect 314270 136232 314326 136288
rect 314394 136232 314450 136288
rect 314518 136232 314574 136288
rect 314642 136232 314698 136288
rect 314766 136232 314822 136288
rect 314890 136232 314946 136288
rect 315014 136232 315070 136288
rect 315138 136232 315194 136288
rect 314022 136108 314078 136164
rect 314146 136108 314202 136164
rect 314270 136108 314326 136164
rect 314394 136108 314450 136164
rect 314518 136108 314574 136164
rect 314642 136108 314698 136164
rect 314766 136108 314822 136164
rect 314890 136108 314946 136164
rect 315014 136108 315070 136164
rect 315138 136108 315194 136164
rect 314022 135984 314078 136040
rect 314146 135984 314202 136040
rect 314270 135984 314326 136040
rect 314394 135984 314450 136040
rect 314518 135984 314574 136040
rect 314642 135984 314698 136040
rect 314766 135984 314822 136040
rect 314890 135984 314946 136040
rect 315014 135984 315070 136040
rect 315138 135984 315194 136040
rect 314022 135860 314078 135916
rect 314146 135860 314202 135916
rect 314270 135860 314326 135916
rect 314394 135860 314450 135916
rect 314518 135860 314574 135916
rect 314642 135860 314698 135916
rect 314766 135860 314822 135916
rect 314890 135860 314946 135916
rect 315014 135860 315070 135916
rect 315138 135860 315194 135916
rect 284022 130356 284078 130412
rect 284146 130356 284202 130412
rect 284270 130356 284326 130412
rect 284394 130356 284450 130412
rect 284518 130356 284574 130412
rect 284642 130356 284698 130412
rect 284766 130356 284822 130412
rect 284890 130356 284946 130412
rect 285014 130356 285070 130412
rect 285138 130356 285194 130412
rect 284022 130232 284078 130288
rect 284146 130232 284202 130288
rect 284270 130232 284326 130288
rect 284394 130232 284450 130288
rect 284518 130232 284574 130288
rect 284642 130232 284698 130288
rect 284766 130232 284822 130288
rect 284890 130232 284946 130288
rect 285014 130232 285070 130288
rect 285138 130232 285194 130288
rect 284022 130108 284078 130164
rect 284146 130108 284202 130164
rect 284270 130108 284326 130164
rect 284394 130108 284450 130164
rect 284518 130108 284574 130164
rect 284642 130108 284698 130164
rect 284766 130108 284822 130164
rect 284890 130108 284946 130164
rect 285014 130108 285070 130164
rect 285138 130108 285194 130164
rect 284022 129984 284078 130040
rect 284146 129984 284202 130040
rect 284270 129984 284326 130040
rect 284394 129984 284450 130040
rect 284518 129984 284574 130040
rect 284642 129984 284698 130040
rect 284766 129984 284822 130040
rect 284890 129984 284946 130040
rect 285014 129984 285070 130040
rect 285138 129984 285194 130040
rect 284022 129860 284078 129916
rect 284146 129860 284202 129916
rect 284270 129860 284326 129916
rect 284394 129860 284450 129916
rect 284518 129860 284574 129916
rect 284642 129860 284698 129916
rect 284766 129860 284822 129916
rect 284890 129860 284946 129916
rect 285014 129860 285070 129916
rect 285138 129860 285194 129916
rect 304022 130356 304078 130412
rect 304146 130356 304202 130412
rect 304270 130356 304326 130412
rect 304394 130356 304450 130412
rect 304518 130356 304574 130412
rect 304642 130356 304698 130412
rect 304766 130356 304822 130412
rect 304890 130356 304946 130412
rect 305014 130356 305070 130412
rect 305138 130356 305194 130412
rect 304022 130232 304078 130288
rect 304146 130232 304202 130288
rect 304270 130232 304326 130288
rect 304394 130232 304450 130288
rect 304518 130232 304574 130288
rect 304642 130232 304698 130288
rect 304766 130232 304822 130288
rect 304890 130232 304946 130288
rect 305014 130232 305070 130288
rect 305138 130232 305194 130288
rect 304022 130108 304078 130164
rect 304146 130108 304202 130164
rect 304270 130108 304326 130164
rect 304394 130108 304450 130164
rect 304518 130108 304574 130164
rect 304642 130108 304698 130164
rect 304766 130108 304822 130164
rect 304890 130108 304946 130164
rect 305014 130108 305070 130164
rect 305138 130108 305194 130164
rect 304022 129984 304078 130040
rect 304146 129984 304202 130040
rect 304270 129984 304326 130040
rect 304394 129984 304450 130040
rect 304518 129984 304574 130040
rect 304642 129984 304698 130040
rect 304766 129984 304822 130040
rect 304890 129984 304946 130040
rect 305014 129984 305070 130040
rect 305138 129984 305194 130040
rect 304022 129860 304078 129916
rect 304146 129860 304202 129916
rect 304270 129860 304326 129916
rect 304394 129860 304450 129916
rect 304518 129860 304574 129916
rect 304642 129860 304698 129916
rect 304766 129860 304822 129916
rect 304890 129860 304946 129916
rect 305014 129860 305070 129916
rect 305138 129860 305194 129916
rect 327250 130294 327306 130350
rect 327374 130294 327430 130350
rect 327498 130294 327554 130350
rect 327622 130294 327678 130350
rect 327250 130170 327306 130226
rect 327374 130170 327430 130226
rect 327498 130170 327554 130226
rect 327622 130170 327678 130226
rect 327250 130046 327306 130102
rect 327374 130046 327430 130102
rect 327498 130046 327554 130102
rect 327622 130046 327678 130102
rect 327250 129922 327306 129978
rect 327374 129922 327430 129978
rect 327498 129922 327554 129978
rect 327622 129922 327678 129978
rect 276970 118294 277026 118350
rect 277094 118294 277150 118350
rect 277218 118294 277274 118350
rect 277342 118294 277398 118350
rect 276970 118170 277026 118226
rect 277094 118170 277150 118226
rect 277218 118170 277274 118226
rect 277342 118170 277398 118226
rect 276970 118046 277026 118102
rect 277094 118046 277150 118102
rect 277218 118046 277274 118102
rect 277342 118046 277398 118102
rect 276970 117922 277026 117978
rect 277094 117922 277150 117978
rect 277218 117922 277274 117978
rect 277342 117922 277398 117978
rect 273250 112294 273306 112350
rect 273374 112294 273430 112350
rect 273498 112294 273554 112350
rect 273622 112294 273678 112350
rect 273250 112170 273306 112226
rect 273374 112170 273430 112226
rect 273498 112170 273554 112226
rect 273622 112170 273678 112226
rect 273250 112046 273306 112102
rect 273374 112046 273430 112102
rect 273498 112046 273554 112102
rect 273622 112046 273678 112102
rect 273250 111922 273306 111978
rect 273374 111922 273430 111978
rect 273498 111922 273554 111978
rect 273622 111922 273678 111978
rect 294022 118356 294078 118412
rect 294146 118356 294202 118412
rect 294270 118356 294326 118412
rect 294394 118356 294450 118412
rect 294518 118356 294574 118412
rect 294642 118356 294698 118412
rect 294766 118356 294822 118412
rect 294890 118356 294946 118412
rect 295014 118356 295070 118412
rect 295138 118356 295194 118412
rect 294022 118232 294078 118288
rect 294146 118232 294202 118288
rect 294270 118232 294326 118288
rect 294394 118232 294450 118288
rect 294518 118232 294574 118288
rect 294642 118232 294698 118288
rect 294766 118232 294822 118288
rect 294890 118232 294946 118288
rect 295014 118232 295070 118288
rect 295138 118232 295194 118288
rect 294022 118108 294078 118164
rect 294146 118108 294202 118164
rect 294270 118108 294326 118164
rect 294394 118108 294450 118164
rect 294518 118108 294574 118164
rect 294642 118108 294698 118164
rect 294766 118108 294822 118164
rect 294890 118108 294946 118164
rect 295014 118108 295070 118164
rect 295138 118108 295194 118164
rect 294022 117984 294078 118040
rect 294146 117984 294202 118040
rect 294270 117984 294326 118040
rect 294394 117984 294450 118040
rect 294518 117984 294574 118040
rect 294642 117984 294698 118040
rect 294766 117984 294822 118040
rect 294890 117984 294946 118040
rect 295014 117984 295070 118040
rect 295138 117984 295194 118040
rect 294022 117860 294078 117916
rect 294146 117860 294202 117916
rect 294270 117860 294326 117916
rect 294394 117860 294450 117916
rect 294518 117860 294574 117916
rect 294642 117860 294698 117916
rect 294766 117860 294822 117916
rect 294890 117860 294946 117916
rect 295014 117860 295070 117916
rect 295138 117860 295194 117916
rect 314022 118356 314078 118412
rect 314146 118356 314202 118412
rect 314270 118356 314326 118412
rect 314394 118356 314450 118412
rect 314518 118356 314574 118412
rect 314642 118356 314698 118412
rect 314766 118356 314822 118412
rect 314890 118356 314946 118412
rect 315014 118356 315070 118412
rect 315138 118356 315194 118412
rect 314022 118232 314078 118288
rect 314146 118232 314202 118288
rect 314270 118232 314326 118288
rect 314394 118232 314450 118288
rect 314518 118232 314574 118288
rect 314642 118232 314698 118288
rect 314766 118232 314822 118288
rect 314890 118232 314946 118288
rect 315014 118232 315070 118288
rect 315138 118232 315194 118288
rect 314022 118108 314078 118164
rect 314146 118108 314202 118164
rect 314270 118108 314326 118164
rect 314394 118108 314450 118164
rect 314518 118108 314574 118164
rect 314642 118108 314698 118164
rect 314766 118108 314822 118164
rect 314890 118108 314946 118164
rect 315014 118108 315070 118164
rect 315138 118108 315194 118164
rect 314022 117984 314078 118040
rect 314146 117984 314202 118040
rect 314270 117984 314326 118040
rect 314394 117984 314450 118040
rect 314518 117984 314574 118040
rect 314642 117984 314698 118040
rect 314766 117984 314822 118040
rect 314890 117984 314946 118040
rect 315014 117984 315070 118040
rect 315138 117984 315194 118040
rect 314022 117860 314078 117916
rect 314146 117860 314202 117916
rect 314270 117860 314326 117916
rect 314394 117860 314450 117916
rect 314518 117860 314574 117916
rect 314642 117860 314698 117916
rect 314766 117860 314822 117916
rect 314890 117860 314946 117916
rect 315014 117860 315070 117916
rect 315138 117860 315194 117916
rect 284022 112356 284078 112412
rect 284146 112356 284202 112412
rect 284270 112356 284326 112412
rect 284394 112356 284450 112412
rect 284518 112356 284574 112412
rect 284642 112356 284698 112412
rect 284766 112356 284822 112412
rect 284890 112356 284946 112412
rect 285014 112356 285070 112412
rect 285138 112356 285194 112412
rect 284022 112232 284078 112288
rect 284146 112232 284202 112288
rect 284270 112232 284326 112288
rect 284394 112232 284450 112288
rect 284518 112232 284574 112288
rect 284642 112232 284698 112288
rect 284766 112232 284822 112288
rect 284890 112232 284946 112288
rect 285014 112232 285070 112288
rect 285138 112232 285194 112288
rect 284022 112108 284078 112164
rect 284146 112108 284202 112164
rect 284270 112108 284326 112164
rect 284394 112108 284450 112164
rect 284518 112108 284574 112164
rect 284642 112108 284698 112164
rect 284766 112108 284822 112164
rect 284890 112108 284946 112164
rect 285014 112108 285070 112164
rect 285138 112108 285194 112164
rect 284022 111984 284078 112040
rect 284146 111984 284202 112040
rect 284270 111984 284326 112040
rect 284394 111984 284450 112040
rect 284518 111984 284574 112040
rect 284642 111984 284698 112040
rect 284766 111984 284822 112040
rect 284890 111984 284946 112040
rect 285014 111984 285070 112040
rect 285138 111984 285194 112040
rect 284022 111860 284078 111916
rect 284146 111860 284202 111916
rect 284270 111860 284326 111916
rect 284394 111860 284450 111916
rect 284518 111860 284574 111916
rect 284642 111860 284698 111916
rect 284766 111860 284822 111916
rect 284890 111860 284946 111916
rect 285014 111860 285070 111916
rect 285138 111860 285194 111916
rect 304022 112356 304078 112412
rect 304146 112356 304202 112412
rect 304270 112356 304326 112412
rect 304394 112356 304450 112412
rect 304518 112356 304574 112412
rect 304642 112356 304698 112412
rect 304766 112356 304822 112412
rect 304890 112356 304946 112412
rect 305014 112356 305070 112412
rect 305138 112356 305194 112412
rect 304022 112232 304078 112288
rect 304146 112232 304202 112288
rect 304270 112232 304326 112288
rect 304394 112232 304450 112288
rect 304518 112232 304574 112288
rect 304642 112232 304698 112288
rect 304766 112232 304822 112288
rect 304890 112232 304946 112288
rect 305014 112232 305070 112288
rect 305138 112232 305194 112288
rect 304022 112108 304078 112164
rect 304146 112108 304202 112164
rect 304270 112108 304326 112164
rect 304394 112108 304450 112164
rect 304518 112108 304574 112164
rect 304642 112108 304698 112164
rect 304766 112108 304822 112164
rect 304890 112108 304946 112164
rect 305014 112108 305070 112164
rect 305138 112108 305194 112164
rect 304022 111984 304078 112040
rect 304146 111984 304202 112040
rect 304270 111984 304326 112040
rect 304394 111984 304450 112040
rect 304518 111984 304574 112040
rect 304642 111984 304698 112040
rect 304766 111984 304822 112040
rect 304890 111984 304946 112040
rect 305014 111984 305070 112040
rect 305138 111984 305194 112040
rect 304022 111860 304078 111916
rect 304146 111860 304202 111916
rect 304270 111860 304326 111916
rect 304394 111860 304450 111916
rect 304518 111860 304574 111916
rect 304642 111860 304698 111916
rect 304766 111860 304822 111916
rect 304890 111860 304946 111916
rect 305014 111860 305070 111916
rect 305138 111860 305194 111916
rect 327250 112294 327306 112350
rect 327374 112294 327430 112350
rect 327498 112294 327554 112350
rect 327622 112294 327678 112350
rect 327250 112170 327306 112226
rect 327374 112170 327430 112226
rect 327498 112170 327554 112226
rect 327622 112170 327678 112226
rect 327250 112046 327306 112102
rect 327374 112046 327430 112102
rect 327498 112046 327554 112102
rect 327622 112046 327678 112102
rect 327250 111922 327306 111978
rect 327374 111922 327430 111978
rect 327498 111922 327554 111978
rect 327622 111922 327678 111978
rect 276970 100294 277026 100350
rect 277094 100294 277150 100350
rect 277218 100294 277274 100350
rect 277342 100294 277398 100350
rect 276970 100170 277026 100226
rect 277094 100170 277150 100226
rect 277218 100170 277274 100226
rect 277342 100170 277398 100226
rect 276970 100046 277026 100102
rect 277094 100046 277150 100102
rect 277218 100046 277274 100102
rect 277342 100046 277398 100102
rect 276970 99922 277026 99978
rect 277094 99922 277150 99978
rect 277218 99922 277274 99978
rect 277342 99922 277398 99978
rect 273250 94294 273306 94350
rect 273374 94294 273430 94350
rect 273498 94294 273554 94350
rect 273622 94294 273678 94350
rect 273250 94170 273306 94226
rect 273374 94170 273430 94226
rect 273498 94170 273554 94226
rect 273622 94170 273678 94226
rect 273250 94046 273306 94102
rect 273374 94046 273430 94102
rect 273498 94046 273554 94102
rect 273622 94046 273678 94102
rect 273250 93922 273306 93978
rect 273374 93922 273430 93978
rect 273498 93922 273554 93978
rect 273622 93922 273678 93978
rect 273250 76294 273306 76350
rect 273374 76294 273430 76350
rect 273498 76294 273554 76350
rect 273622 76294 273678 76350
rect 273250 76170 273306 76226
rect 273374 76170 273430 76226
rect 273498 76170 273554 76226
rect 273622 76170 273678 76226
rect 273250 76046 273306 76102
rect 273374 76046 273430 76102
rect 273498 76046 273554 76102
rect 273622 76046 273678 76102
rect 273250 75922 273306 75978
rect 273374 75922 273430 75978
rect 273498 75922 273554 75978
rect 273622 75922 273678 75978
rect 294022 100356 294078 100412
rect 294146 100356 294202 100412
rect 294270 100356 294326 100412
rect 294394 100356 294450 100412
rect 294518 100356 294574 100412
rect 294642 100356 294698 100412
rect 294766 100356 294822 100412
rect 294890 100356 294946 100412
rect 295014 100356 295070 100412
rect 295138 100356 295194 100412
rect 294022 100232 294078 100288
rect 294146 100232 294202 100288
rect 294270 100232 294326 100288
rect 294394 100232 294450 100288
rect 294518 100232 294574 100288
rect 294642 100232 294698 100288
rect 294766 100232 294822 100288
rect 294890 100232 294946 100288
rect 295014 100232 295070 100288
rect 295138 100232 295194 100288
rect 294022 100108 294078 100164
rect 294146 100108 294202 100164
rect 294270 100108 294326 100164
rect 294394 100108 294450 100164
rect 294518 100108 294574 100164
rect 294642 100108 294698 100164
rect 294766 100108 294822 100164
rect 294890 100108 294946 100164
rect 295014 100108 295070 100164
rect 295138 100108 295194 100164
rect 294022 99984 294078 100040
rect 294146 99984 294202 100040
rect 294270 99984 294326 100040
rect 294394 99984 294450 100040
rect 294518 99984 294574 100040
rect 294642 99984 294698 100040
rect 294766 99984 294822 100040
rect 294890 99984 294946 100040
rect 295014 99984 295070 100040
rect 295138 99984 295194 100040
rect 294022 99860 294078 99916
rect 294146 99860 294202 99916
rect 294270 99860 294326 99916
rect 294394 99860 294450 99916
rect 294518 99860 294574 99916
rect 294642 99860 294698 99916
rect 294766 99860 294822 99916
rect 294890 99860 294946 99916
rect 295014 99860 295070 99916
rect 295138 99860 295194 99916
rect 314022 100356 314078 100412
rect 314146 100356 314202 100412
rect 314270 100356 314326 100412
rect 314394 100356 314450 100412
rect 314518 100356 314574 100412
rect 314642 100356 314698 100412
rect 314766 100356 314822 100412
rect 314890 100356 314946 100412
rect 315014 100356 315070 100412
rect 315138 100356 315194 100412
rect 314022 100232 314078 100288
rect 314146 100232 314202 100288
rect 314270 100232 314326 100288
rect 314394 100232 314450 100288
rect 314518 100232 314574 100288
rect 314642 100232 314698 100288
rect 314766 100232 314822 100288
rect 314890 100232 314946 100288
rect 315014 100232 315070 100288
rect 315138 100232 315194 100288
rect 314022 100108 314078 100164
rect 314146 100108 314202 100164
rect 314270 100108 314326 100164
rect 314394 100108 314450 100164
rect 314518 100108 314574 100164
rect 314642 100108 314698 100164
rect 314766 100108 314822 100164
rect 314890 100108 314946 100164
rect 315014 100108 315070 100164
rect 315138 100108 315194 100164
rect 314022 99984 314078 100040
rect 314146 99984 314202 100040
rect 314270 99984 314326 100040
rect 314394 99984 314450 100040
rect 314518 99984 314574 100040
rect 314642 99984 314698 100040
rect 314766 99984 314822 100040
rect 314890 99984 314946 100040
rect 315014 99984 315070 100040
rect 315138 99984 315194 100040
rect 314022 99860 314078 99916
rect 314146 99860 314202 99916
rect 314270 99860 314326 99916
rect 314394 99860 314450 99916
rect 314518 99860 314574 99916
rect 314642 99860 314698 99916
rect 314766 99860 314822 99916
rect 314890 99860 314946 99916
rect 315014 99860 315070 99916
rect 315138 99860 315194 99916
rect 284022 94356 284078 94412
rect 284146 94356 284202 94412
rect 284270 94356 284326 94412
rect 284394 94356 284450 94412
rect 284518 94356 284574 94412
rect 284642 94356 284698 94412
rect 284766 94356 284822 94412
rect 284890 94356 284946 94412
rect 285014 94356 285070 94412
rect 285138 94356 285194 94412
rect 284022 94232 284078 94288
rect 284146 94232 284202 94288
rect 284270 94232 284326 94288
rect 284394 94232 284450 94288
rect 284518 94232 284574 94288
rect 284642 94232 284698 94288
rect 284766 94232 284822 94288
rect 284890 94232 284946 94288
rect 285014 94232 285070 94288
rect 285138 94232 285194 94288
rect 284022 94108 284078 94164
rect 284146 94108 284202 94164
rect 284270 94108 284326 94164
rect 284394 94108 284450 94164
rect 284518 94108 284574 94164
rect 284642 94108 284698 94164
rect 284766 94108 284822 94164
rect 284890 94108 284946 94164
rect 285014 94108 285070 94164
rect 285138 94108 285194 94164
rect 284022 93984 284078 94040
rect 284146 93984 284202 94040
rect 284270 93984 284326 94040
rect 284394 93984 284450 94040
rect 284518 93984 284574 94040
rect 284642 93984 284698 94040
rect 284766 93984 284822 94040
rect 284890 93984 284946 94040
rect 285014 93984 285070 94040
rect 285138 93984 285194 94040
rect 284022 93860 284078 93916
rect 284146 93860 284202 93916
rect 284270 93860 284326 93916
rect 284394 93860 284450 93916
rect 284518 93860 284574 93916
rect 284642 93860 284698 93916
rect 284766 93860 284822 93916
rect 284890 93860 284946 93916
rect 285014 93860 285070 93916
rect 285138 93860 285194 93916
rect 304022 94356 304078 94412
rect 304146 94356 304202 94412
rect 304270 94356 304326 94412
rect 304394 94356 304450 94412
rect 304518 94356 304574 94412
rect 304642 94356 304698 94412
rect 304766 94356 304822 94412
rect 304890 94356 304946 94412
rect 305014 94356 305070 94412
rect 305138 94356 305194 94412
rect 304022 94232 304078 94288
rect 304146 94232 304202 94288
rect 304270 94232 304326 94288
rect 304394 94232 304450 94288
rect 304518 94232 304574 94288
rect 304642 94232 304698 94288
rect 304766 94232 304822 94288
rect 304890 94232 304946 94288
rect 305014 94232 305070 94288
rect 305138 94232 305194 94288
rect 304022 94108 304078 94164
rect 304146 94108 304202 94164
rect 304270 94108 304326 94164
rect 304394 94108 304450 94164
rect 304518 94108 304574 94164
rect 304642 94108 304698 94164
rect 304766 94108 304822 94164
rect 304890 94108 304946 94164
rect 305014 94108 305070 94164
rect 305138 94108 305194 94164
rect 304022 93984 304078 94040
rect 304146 93984 304202 94040
rect 304270 93984 304326 94040
rect 304394 93984 304450 94040
rect 304518 93984 304574 94040
rect 304642 93984 304698 94040
rect 304766 93984 304822 94040
rect 304890 93984 304946 94040
rect 305014 93984 305070 94040
rect 305138 93984 305194 94040
rect 304022 93860 304078 93916
rect 304146 93860 304202 93916
rect 304270 93860 304326 93916
rect 304394 93860 304450 93916
rect 304518 93860 304574 93916
rect 304642 93860 304698 93916
rect 304766 93860 304822 93916
rect 304890 93860 304946 93916
rect 305014 93860 305070 93916
rect 305138 93860 305194 93916
rect 327250 94294 327306 94350
rect 327374 94294 327430 94350
rect 327498 94294 327554 94350
rect 327622 94294 327678 94350
rect 327250 94170 327306 94226
rect 327374 94170 327430 94226
rect 327498 94170 327554 94226
rect 327622 94170 327678 94226
rect 327250 94046 327306 94102
rect 327374 94046 327430 94102
rect 327498 94046 327554 94102
rect 327622 94046 327678 94102
rect 327250 93922 327306 93978
rect 327374 93922 327430 93978
rect 327498 93922 327554 93978
rect 327622 93922 327678 93978
rect 276970 82294 277026 82350
rect 277094 82294 277150 82350
rect 277218 82294 277274 82350
rect 277342 82294 277398 82350
rect 276970 82170 277026 82226
rect 277094 82170 277150 82226
rect 277218 82170 277274 82226
rect 277342 82170 277398 82226
rect 276970 82046 277026 82102
rect 277094 82046 277150 82102
rect 277218 82046 277274 82102
rect 277342 82046 277398 82102
rect 276970 81922 277026 81978
rect 277094 81922 277150 81978
rect 277218 81922 277274 81978
rect 277342 81922 277398 81978
rect 294022 82356 294078 82412
rect 294146 82356 294202 82412
rect 294270 82356 294326 82412
rect 294394 82356 294450 82412
rect 294518 82356 294574 82412
rect 294642 82356 294698 82412
rect 294766 82356 294822 82412
rect 294890 82356 294946 82412
rect 295014 82356 295070 82412
rect 295138 82356 295194 82412
rect 294022 82232 294078 82288
rect 294146 82232 294202 82288
rect 294270 82232 294326 82288
rect 294394 82232 294450 82288
rect 294518 82232 294574 82288
rect 294642 82232 294698 82288
rect 294766 82232 294822 82288
rect 294890 82232 294946 82288
rect 295014 82232 295070 82288
rect 295138 82232 295194 82288
rect 294022 82108 294078 82164
rect 294146 82108 294202 82164
rect 294270 82108 294326 82164
rect 294394 82108 294450 82164
rect 294518 82108 294574 82164
rect 294642 82108 294698 82164
rect 294766 82108 294822 82164
rect 294890 82108 294946 82164
rect 295014 82108 295070 82164
rect 295138 82108 295194 82164
rect 294022 81984 294078 82040
rect 294146 81984 294202 82040
rect 294270 81984 294326 82040
rect 294394 81984 294450 82040
rect 294518 81984 294574 82040
rect 294642 81984 294698 82040
rect 294766 81984 294822 82040
rect 294890 81984 294946 82040
rect 295014 81984 295070 82040
rect 295138 81984 295194 82040
rect 294022 81860 294078 81916
rect 294146 81860 294202 81916
rect 294270 81860 294326 81916
rect 294394 81860 294450 81916
rect 294518 81860 294574 81916
rect 294642 81860 294698 81916
rect 294766 81860 294822 81916
rect 294890 81860 294946 81916
rect 295014 81860 295070 81916
rect 295138 81860 295194 81916
rect 314022 82356 314078 82412
rect 314146 82356 314202 82412
rect 314270 82356 314326 82412
rect 314394 82356 314450 82412
rect 314518 82356 314574 82412
rect 314642 82356 314698 82412
rect 314766 82356 314822 82412
rect 314890 82356 314946 82412
rect 315014 82356 315070 82412
rect 315138 82356 315194 82412
rect 314022 82232 314078 82288
rect 314146 82232 314202 82288
rect 314270 82232 314326 82288
rect 314394 82232 314450 82288
rect 314518 82232 314574 82288
rect 314642 82232 314698 82288
rect 314766 82232 314822 82288
rect 314890 82232 314946 82288
rect 315014 82232 315070 82288
rect 315138 82232 315194 82288
rect 314022 82108 314078 82164
rect 314146 82108 314202 82164
rect 314270 82108 314326 82164
rect 314394 82108 314450 82164
rect 314518 82108 314574 82164
rect 314642 82108 314698 82164
rect 314766 82108 314822 82164
rect 314890 82108 314946 82164
rect 315014 82108 315070 82164
rect 315138 82108 315194 82164
rect 314022 81984 314078 82040
rect 314146 81984 314202 82040
rect 314270 81984 314326 82040
rect 314394 81984 314450 82040
rect 314518 81984 314574 82040
rect 314642 81984 314698 82040
rect 314766 81984 314822 82040
rect 314890 81984 314946 82040
rect 315014 81984 315070 82040
rect 315138 81984 315194 82040
rect 314022 81860 314078 81916
rect 314146 81860 314202 81916
rect 314270 81860 314326 81916
rect 314394 81860 314450 81916
rect 314518 81860 314574 81916
rect 314642 81860 314698 81916
rect 314766 81860 314822 81916
rect 314890 81860 314946 81916
rect 315014 81860 315070 81916
rect 315138 81860 315194 81916
rect 284022 76356 284078 76412
rect 284146 76356 284202 76412
rect 284270 76356 284326 76412
rect 284394 76356 284450 76412
rect 284518 76356 284574 76412
rect 284642 76356 284698 76412
rect 284766 76356 284822 76412
rect 284890 76356 284946 76412
rect 285014 76356 285070 76412
rect 285138 76356 285194 76412
rect 284022 76232 284078 76288
rect 284146 76232 284202 76288
rect 284270 76232 284326 76288
rect 284394 76232 284450 76288
rect 284518 76232 284574 76288
rect 284642 76232 284698 76288
rect 284766 76232 284822 76288
rect 284890 76232 284946 76288
rect 285014 76232 285070 76288
rect 285138 76232 285194 76288
rect 284022 76108 284078 76164
rect 284146 76108 284202 76164
rect 284270 76108 284326 76164
rect 284394 76108 284450 76164
rect 284518 76108 284574 76164
rect 284642 76108 284698 76164
rect 284766 76108 284822 76164
rect 284890 76108 284946 76164
rect 285014 76108 285070 76164
rect 285138 76108 285194 76164
rect 284022 75984 284078 76040
rect 284146 75984 284202 76040
rect 284270 75984 284326 76040
rect 284394 75984 284450 76040
rect 284518 75984 284574 76040
rect 284642 75984 284698 76040
rect 284766 75984 284822 76040
rect 284890 75984 284946 76040
rect 285014 75984 285070 76040
rect 285138 75984 285194 76040
rect 284022 75860 284078 75916
rect 284146 75860 284202 75916
rect 284270 75860 284326 75916
rect 284394 75860 284450 75916
rect 284518 75860 284574 75916
rect 284642 75860 284698 75916
rect 284766 75860 284822 75916
rect 284890 75860 284946 75916
rect 285014 75860 285070 75916
rect 285138 75860 285194 75916
rect 291250 76294 291306 76350
rect 291374 76294 291430 76350
rect 291498 76294 291554 76350
rect 291622 76294 291678 76350
rect 291250 76170 291306 76226
rect 291374 76170 291430 76226
rect 291498 76170 291554 76226
rect 291622 76170 291678 76226
rect 291250 76046 291306 76102
rect 291374 76046 291430 76102
rect 291498 76046 291554 76102
rect 291622 76046 291678 76102
rect 291250 75922 291306 75978
rect 291374 75922 291430 75978
rect 291498 75922 291554 75978
rect 291622 75922 291678 75978
rect 276970 64294 277026 64350
rect 277094 64294 277150 64350
rect 277218 64294 277274 64350
rect 277342 64294 277398 64350
rect 276970 64170 277026 64226
rect 277094 64170 277150 64226
rect 277218 64170 277274 64226
rect 277342 64170 277398 64226
rect 276970 64046 277026 64102
rect 277094 64046 277150 64102
rect 277218 64046 277274 64102
rect 277342 64046 277398 64102
rect 276970 63922 277026 63978
rect 277094 63922 277150 63978
rect 277218 63922 277274 63978
rect 277342 63922 277398 63978
rect 273250 58294 273306 58350
rect 273374 58294 273430 58350
rect 273498 58294 273554 58350
rect 273622 58294 273678 58350
rect 273250 58170 273306 58226
rect 273374 58170 273430 58226
rect 273498 58170 273554 58226
rect 273622 58170 273678 58226
rect 273250 58046 273306 58102
rect 273374 58046 273430 58102
rect 273498 58046 273554 58102
rect 273622 58046 273678 58102
rect 273250 57922 273306 57978
rect 273374 57922 273430 57978
rect 273498 57922 273554 57978
rect 273622 57922 273678 57978
rect 273250 40294 273306 40350
rect 273374 40294 273430 40350
rect 273498 40294 273554 40350
rect 273622 40294 273678 40350
rect 273250 40170 273306 40226
rect 273374 40170 273430 40226
rect 273498 40170 273554 40226
rect 273622 40170 273678 40226
rect 273250 40046 273306 40102
rect 273374 40046 273430 40102
rect 273498 40046 273554 40102
rect 273622 40046 273678 40102
rect 273250 39922 273306 39978
rect 273374 39922 273430 39978
rect 273498 39922 273554 39978
rect 273622 39922 273678 39978
rect 273250 22294 273306 22350
rect 273374 22294 273430 22350
rect 273498 22294 273554 22350
rect 273622 22294 273678 22350
rect 273250 22170 273306 22226
rect 273374 22170 273430 22226
rect 273498 22170 273554 22226
rect 273622 22170 273678 22226
rect 273250 22046 273306 22102
rect 273374 22046 273430 22102
rect 273498 22046 273554 22102
rect 273622 22046 273678 22102
rect 273250 21922 273306 21978
rect 273374 21922 273430 21978
rect 273498 21922 273554 21978
rect 273622 21922 273678 21978
rect 273250 4294 273306 4350
rect 273374 4294 273430 4350
rect 273498 4294 273554 4350
rect 273622 4294 273678 4350
rect 273250 4170 273306 4226
rect 273374 4170 273430 4226
rect 273498 4170 273554 4226
rect 273622 4170 273678 4226
rect 273250 4046 273306 4102
rect 273374 4046 273430 4102
rect 273498 4046 273554 4102
rect 273622 4046 273678 4102
rect 273250 3922 273306 3978
rect 273374 3922 273430 3978
rect 273498 3922 273554 3978
rect 273622 3922 273678 3978
rect 273250 -216 273306 -160
rect 273374 -216 273430 -160
rect 273498 -216 273554 -160
rect 273622 -216 273678 -160
rect 273250 -340 273306 -284
rect 273374 -340 273430 -284
rect 273498 -340 273554 -284
rect 273622 -340 273678 -284
rect 273250 -464 273306 -408
rect 273374 -464 273430 -408
rect 273498 -464 273554 -408
rect 273622 -464 273678 -408
rect 273250 -588 273306 -532
rect 273374 -588 273430 -532
rect 273498 -588 273554 -532
rect 273622 -588 273678 -532
rect 276970 46294 277026 46350
rect 277094 46294 277150 46350
rect 277218 46294 277274 46350
rect 277342 46294 277398 46350
rect 276970 46170 277026 46226
rect 277094 46170 277150 46226
rect 277218 46170 277274 46226
rect 277342 46170 277398 46226
rect 276970 46046 277026 46102
rect 277094 46046 277150 46102
rect 277218 46046 277274 46102
rect 277342 46046 277398 46102
rect 276970 45922 277026 45978
rect 277094 45922 277150 45978
rect 277218 45922 277274 45978
rect 277342 45922 277398 45978
rect 276970 28294 277026 28350
rect 277094 28294 277150 28350
rect 277218 28294 277274 28350
rect 277342 28294 277398 28350
rect 276970 28170 277026 28226
rect 277094 28170 277150 28226
rect 277218 28170 277274 28226
rect 277342 28170 277398 28226
rect 276970 28046 277026 28102
rect 277094 28046 277150 28102
rect 277218 28046 277274 28102
rect 277342 28046 277398 28102
rect 276970 27922 277026 27978
rect 277094 27922 277150 27978
rect 277218 27922 277274 27978
rect 277342 27922 277398 27978
rect 276970 10294 277026 10350
rect 277094 10294 277150 10350
rect 277218 10294 277274 10350
rect 277342 10294 277398 10350
rect 276970 10170 277026 10226
rect 277094 10170 277150 10226
rect 277218 10170 277274 10226
rect 277342 10170 277398 10226
rect 276970 10046 277026 10102
rect 277094 10046 277150 10102
rect 277218 10046 277274 10102
rect 277342 10046 277398 10102
rect 276970 9922 277026 9978
rect 277094 9922 277150 9978
rect 277218 9922 277274 9978
rect 277342 9922 277398 9978
rect 276970 -1176 277026 -1120
rect 277094 -1176 277150 -1120
rect 277218 -1176 277274 -1120
rect 277342 -1176 277398 -1120
rect 276970 -1300 277026 -1244
rect 277094 -1300 277150 -1244
rect 277218 -1300 277274 -1244
rect 277342 -1300 277398 -1244
rect 276970 -1424 277026 -1368
rect 277094 -1424 277150 -1368
rect 277218 -1424 277274 -1368
rect 277342 -1424 277398 -1368
rect 276970 -1548 277026 -1492
rect 277094 -1548 277150 -1492
rect 277218 -1548 277274 -1492
rect 277342 -1548 277398 -1492
rect 304022 76356 304078 76412
rect 304146 76356 304202 76412
rect 304270 76356 304326 76412
rect 304394 76356 304450 76412
rect 304518 76356 304574 76412
rect 304642 76356 304698 76412
rect 304766 76356 304822 76412
rect 304890 76356 304946 76412
rect 305014 76356 305070 76412
rect 305138 76356 305194 76412
rect 304022 76232 304078 76288
rect 304146 76232 304202 76288
rect 304270 76232 304326 76288
rect 304394 76232 304450 76288
rect 304518 76232 304574 76288
rect 304642 76232 304698 76288
rect 304766 76232 304822 76288
rect 304890 76232 304946 76288
rect 305014 76232 305070 76288
rect 305138 76232 305194 76288
rect 304022 76108 304078 76164
rect 304146 76108 304202 76164
rect 304270 76108 304326 76164
rect 304394 76108 304450 76164
rect 304518 76108 304574 76164
rect 304642 76108 304698 76164
rect 304766 76108 304822 76164
rect 304890 76108 304946 76164
rect 305014 76108 305070 76164
rect 305138 76108 305194 76164
rect 304022 75984 304078 76040
rect 304146 75984 304202 76040
rect 304270 75984 304326 76040
rect 304394 75984 304450 76040
rect 304518 75984 304574 76040
rect 304642 75984 304698 76040
rect 304766 75984 304822 76040
rect 304890 75984 304946 76040
rect 305014 75984 305070 76040
rect 305138 75984 305194 76040
rect 304022 75860 304078 75916
rect 304146 75860 304202 75916
rect 304270 75860 304326 75916
rect 304394 75860 304450 75916
rect 304518 75860 304574 75916
rect 304642 75860 304698 75916
rect 304766 75860 304822 75916
rect 304890 75860 304946 75916
rect 305014 75860 305070 75916
rect 305138 75860 305194 75916
rect 309250 76294 309306 76350
rect 309374 76294 309430 76350
rect 309498 76294 309554 76350
rect 309622 76294 309678 76350
rect 309250 76170 309306 76226
rect 309374 76170 309430 76226
rect 309498 76170 309554 76226
rect 309622 76170 309678 76226
rect 309250 76046 309306 76102
rect 309374 76046 309430 76102
rect 309498 76046 309554 76102
rect 309622 76046 309678 76102
rect 309250 75922 309306 75978
rect 309374 75922 309430 75978
rect 309498 75922 309554 75978
rect 309622 75922 309678 75978
rect 291250 58294 291306 58350
rect 291374 58294 291430 58350
rect 291498 58294 291554 58350
rect 291622 58294 291678 58350
rect 291250 58170 291306 58226
rect 291374 58170 291430 58226
rect 291498 58170 291554 58226
rect 291622 58170 291678 58226
rect 291250 58046 291306 58102
rect 291374 58046 291430 58102
rect 291498 58046 291554 58102
rect 291622 58046 291678 58102
rect 291250 57922 291306 57978
rect 291374 57922 291430 57978
rect 291498 57922 291554 57978
rect 291622 57922 291678 57978
rect 291250 40294 291306 40350
rect 291374 40294 291430 40350
rect 291498 40294 291554 40350
rect 291622 40294 291678 40350
rect 291250 40170 291306 40226
rect 291374 40170 291430 40226
rect 291498 40170 291554 40226
rect 291622 40170 291678 40226
rect 291250 40046 291306 40102
rect 291374 40046 291430 40102
rect 291498 40046 291554 40102
rect 291622 40046 291678 40102
rect 291250 39922 291306 39978
rect 291374 39922 291430 39978
rect 291498 39922 291554 39978
rect 291622 39922 291678 39978
rect 291250 22294 291306 22350
rect 291374 22294 291430 22350
rect 291498 22294 291554 22350
rect 291622 22294 291678 22350
rect 291250 22170 291306 22226
rect 291374 22170 291430 22226
rect 291498 22170 291554 22226
rect 291622 22170 291678 22226
rect 291250 22046 291306 22102
rect 291374 22046 291430 22102
rect 291498 22046 291554 22102
rect 291622 22046 291678 22102
rect 291250 21922 291306 21978
rect 291374 21922 291430 21978
rect 291498 21922 291554 21978
rect 291622 21922 291678 21978
rect 291250 4294 291306 4350
rect 291374 4294 291430 4350
rect 291498 4294 291554 4350
rect 291622 4294 291678 4350
rect 291250 4170 291306 4226
rect 291374 4170 291430 4226
rect 291498 4170 291554 4226
rect 291622 4170 291678 4226
rect 291250 4046 291306 4102
rect 291374 4046 291430 4102
rect 291498 4046 291554 4102
rect 291622 4046 291678 4102
rect 291250 3922 291306 3978
rect 291374 3922 291430 3978
rect 291498 3922 291554 3978
rect 291622 3922 291678 3978
rect 291250 -216 291306 -160
rect 291374 -216 291430 -160
rect 291498 -216 291554 -160
rect 291622 -216 291678 -160
rect 291250 -340 291306 -284
rect 291374 -340 291430 -284
rect 291498 -340 291554 -284
rect 291622 -340 291678 -284
rect 291250 -464 291306 -408
rect 291374 -464 291430 -408
rect 291498 -464 291554 -408
rect 291622 -464 291678 -408
rect 291250 -588 291306 -532
rect 291374 -588 291430 -532
rect 291498 -588 291554 -532
rect 291622 -588 291678 -532
rect 294970 64294 295026 64350
rect 295094 64294 295150 64350
rect 295218 64294 295274 64350
rect 295342 64294 295398 64350
rect 294970 64170 295026 64226
rect 295094 64170 295150 64226
rect 295218 64170 295274 64226
rect 295342 64170 295398 64226
rect 294970 64046 295026 64102
rect 295094 64046 295150 64102
rect 295218 64046 295274 64102
rect 295342 64046 295398 64102
rect 294970 63922 295026 63978
rect 295094 63922 295150 63978
rect 295218 63922 295274 63978
rect 295342 63922 295398 63978
rect 294970 46294 295026 46350
rect 295094 46294 295150 46350
rect 295218 46294 295274 46350
rect 295342 46294 295398 46350
rect 294970 46170 295026 46226
rect 295094 46170 295150 46226
rect 295218 46170 295274 46226
rect 295342 46170 295398 46226
rect 294970 46046 295026 46102
rect 295094 46046 295150 46102
rect 295218 46046 295274 46102
rect 295342 46046 295398 46102
rect 294970 45922 295026 45978
rect 295094 45922 295150 45978
rect 295218 45922 295274 45978
rect 295342 45922 295398 45978
rect 294970 28294 295026 28350
rect 295094 28294 295150 28350
rect 295218 28294 295274 28350
rect 295342 28294 295398 28350
rect 294970 28170 295026 28226
rect 295094 28170 295150 28226
rect 295218 28170 295274 28226
rect 295342 28170 295398 28226
rect 294970 28046 295026 28102
rect 295094 28046 295150 28102
rect 295218 28046 295274 28102
rect 295342 28046 295398 28102
rect 294970 27922 295026 27978
rect 295094 27922 295150 27978
rect 295218 27922 295274 27978
rect 295342 27922 295398 27978
rect 294970 10294 295026 10350
rect 295094 10294 295150 10350
rect 295218 10294 295274 10350
rect 295342 10294 295398 10350
rect 294970 10170 295026 10226
rect 295094 10170 295150 10226
rect 295218 10170 295274 10226
rect 295342 10170 295398 10226
rect 294970 10046 295026 10102
rect 295094 10046 295150 10102
rect 295218 10046 295274 10102
rect 295342 10046 295398 10102
rect 294970 9922 295026 9978
rect 295094 9922 295150 9978
rect 295218 9922 295274 9978
rect 295342 9922 295398 9978
rect 294970 -1176 295026 -1120
rect 295094 -1176 295150 -1120
rect 295218 -1176 295274 -1120
rect 295342 -1176 295398 -1120
rect 294970 -1300 295026 -1244
rect 295094 -1300 295150 -1244
rect 295218 -1300 295274 -1244
rect 295342 -1300 295398 -1244
rect 294970 -1424 295026 -1368
rect 295094 -1424 295150 -1368
rect 295218 -1424 295274 -1368
rect 295342 -1424 295398 -1368
rect 294970 -1548 295026 -1492
rect 295094 -1548 295150 -1492
rect 295218 -1548 295274 -1492
rect 295342 -1548 295398 -1492
rect 309250 58294 309306 58350
rect 309374 58294 309430 58350
rect 309498 58294 309554 58350
rect 309622 58294 309678 58350
rect 309250 58170 309306 58226
rect 309374 58170 309430 58226
rect 309498 58170 309554 58226
rect 309622 58170 309678 58226
rect 309250 58046 309306 58102
rect 309374 58046 309430 58102
rect 309498 58046 309554 58102
rect 309622 58046 309678 58102
rect 309250 57922 309306 57978
rect 309374 57922 309430 57978
rect 309498 57922 309554 57978
rect 309622 57922 309678 57978
rect 309250 40294 309306 40350
rect 309374 40294 309430 40350
rect 309498 40294 309554 40350
rect 309622 40294 309678 40350
rect 309250 40170 309306 40226
rect 309374 40170 309430 40226
rect 309498 40170 309554 40226
rect 309622 40170 309678 40226
rect 309250 40046 309306 40102
rect 309374 40046 309430 40102
rect 309498 40046 309554 40102
rect 309622 40046 309678 40102
rect 309250 39922 309306 39978
rect 309374 39922 309430 39978
rect 309498 39922 309554 39978
rect 309622 39922 309678 39978
rect 309250 22294 309306 22350
rect 309374 22294 309430 22350
rect 309498 22294 309554 22350
rect 309622 22294 309678 22350
rect 309250 22170 309306 22226
rect 309374 22170 309430 22226
rect 309498 22170 309554 22226
rect 309622 22170 309678 22226
rect 309250 22046 309306 22102
rect 309374 22046 309430 22102
rect 309498 22046 309554 22102
rect 309622 22046 309678 22102
rect 309250 21922 309306 21978
rect 309374 21922 309430 21978
rect 309498 21922 309554 21978
rect 309622 21922 309678 21978
rect 309250 4294 309306 4350
rect 309374 4294 309430 4350
rect 309498 4294 309554 4350
rect 309622 4294 309678 4350
rect 309250 4170 309306 4226
rect 309374 4170 309430 4226
rect 309498 4170 309554 4226
rect 309622 4170 309678 4226
rect 309250 4046 309306 4102
rect 309374 4046 309430 4102
rect 309498 4046 309554 4102
rect 309622 4046 309678 4102
rect 309250 3922 309306 3978
rect 309374 3922 309430 3978
rect 309498 3922 309554 3978
rect 309622 3922 309678 3978
rect 309250 -216 309306 -160
rect 309374 -216 309430 -160
rect 309498 -216 309554 -160
rect 309622 -216 309678 -160
rect 309250 -340 309306 -284
rect 309374 -340 309430 -284
rect 309498 -340 309554 -284
rect 309622 -340 309678 -284
rect 309250 -464 309306 -408
rect 309374 -464 309430 -408
rect 309498 -464 309554 -408
rect 309622 -464 309678 -408
rect 309250 -588 309306 -532
rect 309374 -588 309430 -532
rect 309498 -588 309554 -532
rect 309622 -588 309678 -532
rect 312970 64294 313026 64350
rect 313094 64294 313150 64350
rect 313218 64294 313274 64350
rect 313342 64294 313398 64350
rect 312970 64170 313026 64226
rect 313094 64170 313150 64226
rect 313218 64170 313274 64226
rect 313342 64170 313398 64226
rect 312970 64046 313026 64102
rect 313094 64046 313150 64102
rect 313218 64046 313274 64102
rect 313342 64046 313398 64102
rect 312970 63922 313026 63978
rect 313094 63922 313150 63978
rect 313218 63922 313274 63978
rect 313342 63922 313398 63978
rect 312970 46294 313026 46350
rect 313094 46294 313150 46350
rect 313218 46294 313274 46350
rect 313342 46294 313398 46350
rect 312970 46170 313026 46226
rect 313094 46170 313150 46226
rect 313218 46170 313274 46226
rect 313342 46170 313398 46226
rect 312970 46046 313026 46102
rect 313094 46046 313150 46102
rect 313218 46046 313274 46102
rect 313342 46046 313398 46102
rect 312970 45922 313026 45978
rect 313094 45922 313150 45978
rect 313218 45922 313274 45978
rect 313342 45922 313398 45978
rect 312970 28294 313026 28350
rect 313094 28294 313150 28350
rect 313218 28294 313274 28350
rect 313342 28294 313398 28350
rect 312970 28170 313026 28226
rect 313094 28170 313150 28226
rect 313218 28170 313274 28226
rect 313342 28170 313398 28226
rect 312970 28046 313026 28102
rect 313094 28046 313150 28102
rect 313218 28046 313274 28102
rect 313342 28046 313398 28102
rect 312970 27922 313026 27978
rect 313094 27922 313150 27978
rect 313218 27922 313274 27978
rect 313342 27922 313398 27978
rect 312970 10294 313026 10350
rect 313094 10294 313150 10350
rect 313218 10294 313274 10350
rect 313342 10294 313398 10350
rect 312970 10170 313026 10226
rect 313094 10170 313150 10226
rect 313218 10170 313274 10226
rect 313342 10170 313398 10226
rect 312970 10046 313026 10102
rect 313094 10046 313150 10102
rect 313218 10046 313274 10102
rect 313342 10046 313398 10102
rect 312970 9922 313026 9978
rect 313094 9922 313150 9978
rect 313218 9922 313274 9978
rect 313342 9922 313398 9978
rect 312970 -1176 313026 -1120
rect 313094 -1176 313150 -1120
rect 313218 -1176 313274 -1120
rect 313342 -1176 313398 -1120
rect 312970 -1300 313026 -1244
rect 313094 -1300 313150 -1244
rect 313218 -1300 313274 -1244
rect 313342 -1300 313398 -1244
rect 312970 -1424 313026 -1368
rect 313094 -1424 313150 -1368
rect 313218 -1424 313274 -1368
rect 313342 -1424 313398 -1368
rect 312970 -1548 313026 -1492
rect 313094 -1548 313150 -1492
rect 313218 -1548 313274 -1492
rect 313342 -1548 313398 -1492
rect 327250 76294 327306 76350
rect 327374 76294 327430 76350
rect 327498 76294 327554 76350
rect 327622 76294 327678 76350
rect 327250 76170 327306 76226
rect 327374 76170 327430 76226
rect 327498 76170 327554 76226
rect 327622 76170 327678 76226
rect 327250 76046 327306 76102
rect 327374 76046 327430 76102
rect 327498 76046 327554 76102
rect 327622 76046 327678 76102
rect 327250 75922 327306 75978
rect 327374 75922 327430 75978
rect 327498 75922 327554 75978
rect 327622 75922 327678 75978
rect 327250 58294 327306 58350
rect 327374 58294 327430 58350
rect 327498 58294 327554 58350
rect 327622 58294 327678 58350
rect 327250 58170 327306 58226
rect 327374 58170 327430 58226
rect 327498 58170 327554 58226
rect 327622 58170 327678 58226
rect 327250 58046 327306 58102
rect 327374 58046 327430 58102
rect 327498 58046 327554 58102
rect 327622 58046 327678 58102
rect 327250 57922 327306 57978
rect 327374 57922 327430 57978
rect 327498 57922 327554 57978
rect 327622 57922 327678 57978
rect 327250 40294 327306 40350
rect 327374 40294 327430 40350
rect 327498 40294 327554 40350
rect 327622 40294 327678 40350
rect 327250 40170 327306 40226
rect 327374 40170 327430 40226
rect 327498 40170 327554 40226
rect 327622 40170 327678 40226
rect 327250 40046 327306 40102
rect 327374 40046 327430 40102
rect 327498 40046 327554 40102
rect 327622 40046 327678 40102
rect 327250 39922 327306 39978
rect 327374 39922 327430 39978
rect 327498 39922 327554 39978
rect 327622 39922 327678 39978
rect 327250 22294 327306 22350
rect 327374 22294 327430 22350
rect 327498 22294 327554 22350
rect 327622 22294 327678 22350
rect 327250 22170 327306 22226
rect 327374 22170 327430 22226
rect 327498 22170 327554 22226
rect 327622 22170 327678 22226
rect 327250 22046 327306 22102
rect 327374 22046 327430 22102
rect 327498 22046 327554 22102
rect 327622 22046 327678 22102
rect 327250 21922 327306 21978
rect 327374 21922 327430 21978
rect 327498 21922 327554 21978
rect 327622 21922 327678 21978
rect 327250 4294 327306 4350
rect 327374 4294 327430 4350
rect 327498 4294 327554 4350
rect 327622 4294 327678 4350
rect 327250 4170 327306 4226
rect 327374 4170 327430 4226
rect 327498 4170 327554 4226
rect 327622 4170 327678 4226
rect 327250 4046 327306 4102
rect 327374 4046 327430 4102
rect 327498 4046 327554 4102
rect 327622 4046 327678 4102
rect 327250 3922 327306 3978
rect 327374 3922 327430 3978
rect 327498 3922 327554 3978
rect 327622 3922 327678 3978
rect 327250 -216 327306 -160
rect 327374 -216 327430 -160
rect 327498 -216 327554 -160
rect 327622 -216 327678 -160
rect 327250 -340 327306 -284
rect 327374 -340 327430 -284
rect 327498 -340 327554 -284
rect 327622 -340 327678 -284
rect 327250 -464 327306 -408
rect 327374 -464 327430 -408
rect 327498 -464 327554 -408
rect 327622 -464 327678 -408
rect 327250 -588 327306 -532
rect 327374 -588 327430 -532
rect 327498 -588 327554 -532
rect 327622 -588 327678 -532
rect 330970 598116 331026 598172
rect 331094 598116 331150 598172
rect 331218 598116 331274 598172
rect 331342 598116 331398 598172
rect 330970 597992 331026 598048
rect 331094 597992 331150 598048
rect 331218 597992 331274 598048
rect 331342 597992 331398 598048
rect 330970 597868 331026 597924
rect 331094 597868 331150 597924
rect 331218 597868 331274 597924
rect 331342 597868 331398 597924
rect 330970 597744 331026 597800
rect 331094 597744 331150 597800
rect 331218 597744 331274 597800
rect 331342 597744 331398 597800
rect 330970 586294 331026 586350
rect 331094 586294 331150 586350
rect 331218 586294 331274 586350
rect 331342 586294 331398 586350
rect 330970 586170 331026 586226
rect 331094 586170 331150 586226
rect 331218 586170 331274 586226
rect 331342 586170 331398 586226
rect 330970 586046 331026 586102
rect 331094 586046 331150 586102
rect 331218 586046 331274 586102
rect 331342 586046 331398 586102
rect 330970 585922 331026 585978
rect 331094 585922 331150 585978
rect 331218 585922 331274 585978
rect 331342 585922 331398 585978
rect 330970 568294 331026 568350
rect 331094 568294 331150 568350
rect 331218 568294 331274 568350
rect 331342 568294 331398 568350
rect 330970 568170 331026 568226
rect 331094 568170 331150 568226
rect 331218 568170 331274 568226
rect 331342 568170 331398 568226
rect 330970 568046 331026 568102
rect 331094 568046 331150 568102
rect 331218 568046 331274 568102
rect 331342 568046 331398 568102
rect 330970 567922 331026 567978
rect 331094 567922 331150 567978
rect 331218 567922 331274 567978
rect 331342 567922 331398 567978
rect 330970 550294 331026 550350
rect 331094 550294 331150 550350
rect 331218 550294 331274 550350
rect 331342 550294 331398 550350
rect 330970 550170 331026 550226
rect 331094 550170 331150 550226
rect 331218 550170 331274 550226
rect 331342 550170 331398 550226
rect 330970 550046 331026 550102
rect 331094 550046 331150 550102
rect 331218 550046 331274 550102
rect 331342 550046 331398 550102
rect 330970 549922 331026 549978
rect 331094 549922 331150 549978
rect 331218 549922 331274 549978
rect 331342 549922 331398 549978
rect 330970 532294 331026 532350
rect 331094 532294 331150 532350
rect 331218 532294 331274 532350
rect 331342 532294 331398 532350
rect 330970 532170 331026 532226
rect 331094 532170 331150 532226
rect 331218 532170 331274 532226
rect 331342 532170 331398 532226
rect 330970 532046 331026 532102
rect 331094 532046 331150 532102
rect 331218 532046 331274 532102
rect 331342 532046 331398 532102
rect 330970 531922 331026 531978
rect 331094 531922 331150 531978
rect 331218 531922 331274 531978
rect 331342 531922 331398 531978
rect 330970 514294 331026 514350
rect 331094 514294 331150 514350
rect 331218 514294 331274 514350
rect 331342 514294 331398 514350
rect 330970 514170 331026 514226
rect 331094 514170 331150 514226
rect 331218 514170 331274 514226
rect 331342 514170 331398 514226
rect 330970 514046 331026 514102
rect 331094 514046 331150 514102
rect 331218 514046 331274 514102
rect 331342 514046 331398 514102
rect 330970 513922 331026 513978
rect 331094 513922 331150 513978
rect 331218 513922 331274 513978
rect 331342 513922 331398 513978
rect 330970 496294 331026 496350
rect 331094 496294 331150 496350
rect 331218 496294 331274 496350
rect 331342 496294 331398 496350
rect 330970 496170 331026 496226
rect 331094 496170 331150 496226
rect 331218 496170 331274 496226
rect 331342 496170 331398 496226
rect 330970 496046 331026 496102
rect 331094 496046 331150 496102
rect 331218 496046 331274 496102
rect 331342 496046 331398 496102
rect 330970 495922 331026 495978
rect 331094 495922 331150 495978
rect 331218 495922 331274 495978
rect 331342 495922 331398 495978
rect 330970 478294 331026 478350
rect 331094 478294 331150 478350
rect 331218 478294 331274 478350
rect 331342 478294 331398 478350
rect 330970 478170 331026 478226
rect 331094 478170 331150 478226
rect 331218 478170 331274 478226
rect 331342 478170 331398 478226
rect 330970 478046 331026 478102
rect 331094 478046 331150 478102
rect 331218 478046 331274 478102
rect 331342 478046 331398 478102
rect 330970 477922 331026 477978
rect 331094 477922 331150 477978
rect 331218 477922 331274 477978
rect 331342 477922 331398 477978
rect 330970 460294 331026 460350
rect 331094 460294 331150 460350
rect 331218 460294 331274 460350
rect 331342 460294 331398 460350
rect 330970 460170 331026 460226
rect 331094 460170 331150 460226
rect 331218 460170 331274 460226
rect 331342 460170 331398 460226
rect 330970 460046 331026 460102
rect 331094 460046 331150 460102
rect 331218 460046 331274 460102
rect 331342 460046 331398 460102
rect 330970 459922 331026 459978
rect 331094 459922 331150 459978
rect 331218 459922 331274 459978
rect 331342 459922 331398 459978
rect 330970 442294 331026 442350
rect 331094 442294 331150 442350
rect 331218 442294 331274 442350
rect 331342 442294 331398 442350
rect 330970 442170 331026 442226
rect 331094 442170 331150 442226
rect 331218 442170 331274 442226
rect 331342 442170 331398 442226
rect 330970 442046 331026 442102
rect 331094 442046 331150 442102
rect 331218 442046 331274 442102
rect 331342 442046 331398 442102
rect 330970 441922 331026 441978
rect 331094 441922 331150 441978
rect 331218 441922 331274 441978
rect 331342 441922 331398 441978
rect 330970 424294 331026 424350
rect 331094 424294 331150 424350
rect 331218 424294 331274 424350
rect 331342 424294 331398 424350
rect 330970 424170 331026 424226
rect 331094 424170 331150 424226
rect 331218 424170 331274 424226
rect 331342 424170 331398 424226
rect 330970 424046 331026 424102
rect 331094 424046 331150 424102
rect 331218 424046 331274 424102
rect 331342 424046 331398 424102
rect 330970 423922 331026 423978
rect 331094 423922 331150 423978
rect 331218 423922 331274 423978
rect 331342 423922 331398 423978
rect 330970 406294 331026 406350
rect 331094 406294 331150 406350
rect 331218 406294 331274 406350
rect 331342 406294 331398 406350
rect 330970 406170 331026 406226
rect 331094 406170 331150 406226
rect 331218 406170 331274 406226
rect 331342 406170 331398 406226
rect 330970 406046 331026 406102
rect 331094 406046 331150 406102
rect 331218 406046 331274 406102
rect 331342 406046 331398 406102
rect 330970 405922 331026 405978
rect 331094 405922 331150 405978
rect 331218 405922 331274 405978
rect 331342 405922 331398 405978
rect 330970 388294 331026 388350
rect 331094 388294 331150 388350
rect 331218 388294 331274 388350
rect 331342 388294 331398 388350
rect 330970 388170 331026 388226
rect 331094 388170 331150 388226
rect 331218 388170 331274 388226
rect 331342 388170 331398 388226
rect 330970 388046 331026 388102
rect 331094 388046 331150 388102
rect 331218 388046 331274 388102
rect 331342 388046 331398 388102
rect 330970 387922 331026 387978
rect 331094 387922 331150 387978
rect 331218 387922 331274 387978
rect 331342 387922 331398 387978
rect 330970 370294 331026 370350
rect 331094 370294 331150 370350
rect 331218 370294 331274 370350
rect 331342 370294 331398 370350
rect 330970 370170 331026 370226
rect 331094 370170 331150 370226
rect 331218 370170 331274 370226
rect 331342 370170 331398 370226
rect 330970 370046 331026 370102
rect 331094 370046 331150 370102
rect 331218 370046 331274 370102
rect 331342 370046 331398 370102
rect 330970 369922 331026 369978
rect 331094 369922 331150 369978
rect 331218 369922 331274 369978
rect 331342 369922 331398 369978
rect 330970 352294 331026 352350
rect 331094 352294 331150 352350
rect 331218 352294 331274 352350
rect 331342 352294 331398 352350
rect 330970 352170 331026 352226
rect 331094 352170 331150 352226
rect 331218 352170 331274 352226
rect 331342 352170 331398 352226
rect 330970 352046 331026 352102
rect 331094 352046 331150 352102
rect 331218 352046 331274 352102
rect 331342 352046 331398 352102
rect 330970 351922 331026 351978
rect 331094 351922 331150 351978
rect 331218 351922 331274 351978
rect 331342 351922 331398 351978
rect 330970 334294 331026 334350
rect 331094 334294 331150 334350
rect 331218 334294 331274 334350
rect 331342 334294 331398 334350
rect 330970 334170 331026 334226
rect 331094 334170 331150 334226
rect 331218 334170 331274 334226
rect 331342 334170 331398 334226
rect 330970 334046 331026 334102
rect 331094 334046 331150 334102
rect 331218 334046 331274 334102
rect 331342 334046 331398 334102
rect 330970 333922 331026 333978
rect 331094 333922 331150 333978
rect 331218 333922 331274 333978
rect 331342 333922 331398 333978
rect 330970 316294 331026 316350
rect 331094 316294 331150 316350
rect 331218 316294 331274 316350
rect 331342 316294 331398 316350
rect 330970 316170 331026 316226
rect 331094 316170 331150 316226
rect 331218 316170 331274 316226
rect 331342 316170 331398 316226
rect 330970 316046 331026 316102
rect 331094 316046 331150 316102
rect 331218 316046 331274 316102
rect 331342 316046 331398 316102
rect 330970 315922 331026 315978
rect 331094 315922 331150 315978
rect 331218 315922 331274 315978
rect 331342 315922 331398 315978
rect 330970 298294 331026 298350
rect 331094 298294 331150 298350
rect 331218 298294 331274 298350
rect 331342 298294 331398 298350
rect 330970 298170 331026 298226
rect 331094 298170 331150 298226
rect 331218 298170 331274 298226
rect 331342 298170 331398 298226
rect 330970 298046 331026 298102
rect 331094 298046 331150 298102
rect 331218 298046 331274 298102
rect 331342 298046 331398 298102
rect 330970 297922 331026 297978
rect 331094 297922 331150 297978
rect 331218 297922 331274 297978
rect 331342 297922 331398 297978
rect 330970 280294 331026 280350
rect 331094 280294 331150 280350
rect 331218 280294 331274 280350
rect 331342 280294 331398 280350
rect 330970 280170 331026 280226
rect 331094 280170 331150 280226
rect 331218 280170 331274 280226
rect 331342 280170 331398 280226
rect 330970 280046 331026 280102
rect 331094 280046 331150 280102
rect 331218 280046 331274 280102
rect 331342 280046 331398 280102
rect 330970 279922 331026 279978
rect 331094 279922 331150 279978
rect 331218 279922 331274 279978
rect 331342 279922 331398 279978
rect 330970 262294 331026 262350
rect 331094 262294 331150 262350
rect 331218 262294 331274 262350
rect 331342 262294 331398 262350
rect 330970 262170 331026 262226
rect 331094 262170 331150 262226
rect 331218 262170 331274 262226
rect 331342 262170 331398 262226
rect 330970 262046 331026 262102
rect 331094 262046 331150 262102
rect 331218 262046 331274 262102
rect 331342 262046 331398 262102
rect 330970 261922 331026 261978
rect 331094 261922 331150 261978
rect 331218 261922 331274 261978
rect 331342 261922 331398 261978
rect 330970 244294 331026 244350
rect 331094 244294 331150 244350
rect 331218 244294 331274 244350
rect 331342 244294 331398 244350
rect 330970 244170 331026 244226
rect 331094 244170 331150 244226
rect 331218 244170 331274 244226
rect 331342 244170 331398 244226
rect 330970 244046 331026 244102
rect 331094 244046 331150 244102
rect 331218 244046 331274 244102
rect 331342 244046 331398 244102
rect 330970 243922 331026 243978
rect 331094 243922 331150 243978
rect 331218 243922 331274 243978
rect 331342 243922 331398 243978
rect 348970 598116 349026 598172
rect 349094 598116 349150 598172
rect 349218 598116 349274 598172
rect 349342 598116 349398 598172
rect 348970 597992 349026 598048
rect 349094 597992 349150 598048
rect 349218 597992 349274 598048
rect 349342 597992 349398 598048
rect 348970 597868 349026 597924
rect 349094 597868 349150 597924
rect 349218 597868 349274 597924
rect 349342 597868 349398 597924
rect 348970 597744 349026 597800
rect 349094 597744 349150 597800
rect 349218 597744 349274 597800
rect 349342 597744 349398 597800
rect 348970 586294 349026 586350
rect 349094 586294 349150 586350
rect 349218 586294 349274 586350
rect 349342 586294 349398 586350
rect 348970 586170 349026 586226
rect 349094 586170 349150 586226
rect 349218 586170 349274 586226
rect 349342 586170 349398 586226
rect 348970 586046 349026 586102
rect 349094 586046 349150 586102
rect 349218 586046 349274 586102
rect 349342 586046 349398 586102
rect 348970 585922 349026 585978
rect 349094 585922 349150 585978
rect 349218 585922 349274 585978
rect 349342 585922 349398 585978
rect 348970 568294 349026 568350
rect 349094 568294 349150 568350
rect 349218 568294 349274 568350
rect 349342 568294 349398 568350
rect 348970 568170 349026 568226
rect 349094 568170 349150 568226
rect 349218 568170 349274 568226
rect 349342 568170 349398 568226
rect 348970 568046 349026 568102
rect 349094 568046 349150 568102
rect 349218 568046 349274 568102
rect 349342 568046 349398 568102
rect 348970 567922 349026 567978
rect 349094 567922 349150 567978
rect 349218 567922 349274 567978
rect 349342 567922 349398 567978
rect 348970 550294 349026 550350
rect 349094 550294 349150 550350
rect 349218 550294 349274 550350
rect 349342 550294 349398 550350
rect 348970 550170 349026 550226
rect 349094 550170 349150 550226
rect 349218 550170 349274 550226
rect 349342 550170 349398 550226
rect 348970 550046 349026 550102
rect 349094 550046 349150 550102
rect 349218 550046 349274 550102
rect 349342 550046 349398 550102
rect 348970 549922 349026 549978
rect 349094 549922 349150 549978
rect 349218 549922 349274 549978
rect 349342 549922 349398 549978
rect 348970 532294 349026 532350
rect 349094 532294 349150 532350
rect 349218 532294 349274 532350
rect 349342 532294 349398 532350
rect 348970 532170 349026 532226
rect 349094 532170 349150 532226
rect 349218 532170 349274 532226
rect 349342 532170 349398 532226
rect 348970 532046 349026 532102
rect 349094 532046 349150 532102
rect 349218 532046 349274 532102
rect 349342 532046 349398 532102
rect 348970 531922 349026 531978
rect 349094 531922 349150 531978
rect 349218 531922 349274 531978
rect 349342 531922 349398 531978
rect 348970 514294 349026 514350
rect 349094 514294 349150 514350
rect 349218 514294 349274 514350
rect 349342 514294 349398 514350
rect 348970 514170 349026 514226
rect 349094 514170 349150 514226
rect 349218 514170 349274 514226
rect 349342 514170 349398 514226
rect 348970 514046 349026 514102
rect 349094 514046 349150 514102
rect 349218 514046 349274 514102
rect 349342 514046 349398 514102
rect 348970 513922 349026 513978
rect 349094 513922 349150 513978
rect 349218 513922 349274 513978
rect 349342 513922 349398 513978
rect 348970 496294 349026 496350
rect 349094 496294 349150 496350
rect 349218 496294 349274 496350
rect 349342 496294 349398 496350
rect 348970 496170 349026 496226
rect 349094 496170 349150 496226
rect 349218 496170 349274 496226
rect 349342 496170 349398 496226
rect 348970 496046 349026 496102
rect 349094 496046 349150 496102
rect 349218 496046 349274 496102
rect 349342 496046 349398 496102
rect 348970 495922 349026 495978
rect 349094 495922 349150 495978
rect 349218 495922 349274 495978
rect 349342 495922 349398 495978
rect 348970 478294 349026 478350
rect 349094 478294 349150 478350
rect 349218 478294 349274 478350
rect 349342 478294 349398 478350
rect 348970 478170 349026 478226
rect 349094 478170 349150 478226
rect 349218 478170 349274 478226
rect 349342 478170 349398 478226
rect 348970 478046 349026 478102
rect 349094 478046 349150 478102
rect 349218 478046 349274 478102
rect 349342 478046 349398 478102
rect 348970 477922 349026 477978
rect 349094 477922 349150 477978
rect 349218 477922 349274 477978
rect 349342 477922 349398 477978
rect 348970 460294 349026 460350
rect 349094 460294 349150 460350
rect 349218 460294 349274 460350
rect 349342 460294 349398 460350
rect 348970 460170 349026 460226
rect 349094 460170 349150 460226
rect 349218 460170 349274 460226
rect 349342 460170 349398 460226
rect 348970 460046 349026 460102
rect 349094 460046 349150 460102
rect 349218 460046 349274 460102
rect 349342 460046 349398 460102
rect 348970 459922 349026 459978
rect 349094 459922 349150 459978
rect 349218 459922 349274 459978
rect 349342 459922 349398 459978
rect 348970 442294 349026 442350
rect 349094 442294 349150 442350
rect 349218 442294 349274 442350
rect 349342 442294 349398 442350
rect 348970 442170 349026 442226
rect 349094 442170 349150 442226
rect 349218 442170 349274 442226
rect 349342 442170 349398 442226
rect 348970 442046 349026 442102
rect 349094 442046 349150 442102
rect 349218 442046 349274 442102
rect 349342 442046 349398 442102
rect 348970 441922 349026 441978
rect 349094 441922 349150 441978
rect 349218 441922 349274 441978
rect 349342 441922 349398 441978
rect 348970 424294 349026 424350
rect 349094 424294 349150 424350
rect 349218 424294 349274 424350
rect 349342 424294 349398 424350
rect 348970 424170 349026 424226
rect 349094 424170 349150 424226
rect 349218 424170 349274 424226
rect 349342 424170 349398 424226
rect 348970 424046 349026 424102
rect 349094 424046 349150 424102
rect 349218 424046 349274 424102
rect 349342 424046 349398 424102
rect 348970 423922 349026 423978
rect 349094 423922 349150 423978
rect 349218 423922 349274 423978
rect 349342 423922 349398 423978
rect 348970 406294 349026 406350
rect 349094 406294 349150 406350
rect 349218 406294 349274 406350
rect 349342 406294 349398 406350
rect 348970 406170 349026 406226
rect 349094 406170 349150 406226
rect 349218 406170 349274 406226
rect 349342 406170 349398 406226
rect 348970 406046 349026 406102
rect 349094 406046 349150 406102
rect 349218 406046 349274 406102
rect 349342 406046 349398 406102
rect 348970 405922 349026 405978
rect 349094 405922 349150 405978
rect 349218 405922 349274 405978
rect 349342 405922 349398 405978
rect 348970 388294 349026 388350
rect 349094 388294 349150 388350
rect 349218 388294 349274 388350
rect 349342 388294 349398 388350
rect 348970 388170 349026 388226
rect 349094 388170 349150 388226
rect 349218 388170 349274 388226
rect 349342 388170 349398 388226
rect 348970 388046 349026 388102
rect 349094 388046 349150 388102
rect 349218 388046 349274 388102
rect 349342 388046 349398 388102
rect 348970 387922 349026 387978
rect 349094 387922 349150 387978
rect 349218 387922 349274 387978
rect 349342 387922 349398 387978
rect 348970 370294 349026 370350
rect 349094 370294 349150 370350
rect 349218 370294 349274 370350
rect 349342 370294 349398 370350
rect 348970 370170 349026 370226
rect 349094 370170 349150 370226
rect 349218 370170 349274 370226
rect 349342 370170 349398 370226
rect 348970 370046 349026 370102
rect 349094 370046 349150 370102
rect 349218 370046 349274 370102
rect 349342 370046 349398 370102
rect 348970 369922 349026 369978
rect 349094 369922 349150 369978
rect 349218 369922 349274 369978
rect 349342 369922 349398 369978
rect 348970 352294 349026 352350
rect 349094 352294 349150 352350
rect 349218 352294 349274 352350
rect 349342 352294 349398 352350
rect 348970 352170 349026 352226
rect 349094 352170 349150 352226
rect 349218 352170 349274 352226
rect 349342 352170 349398 352226
rect 348970 352046 349026 352102
rect 349094 352046 349150 352102
rect 349218 352046 349274 352102
rect 349342 352046 349398 352102
rect 348970 351922 349026 351978
rect 349094 351922 349150 351978
rect 349218 351922 349274 351978
rect 349342 351922 349398 351978
rect 348970 334294 349026 334350
rect 349094 334294 349150 334350
rect 349218 334294 349274 334350
rect 349342 334294 349398 334350
rect 348970 334170 349026 334226
rect 349094 334170 349150 334226
rect 349218 334170 349274 334226
rect 349342 334170 349398 334226
rect 348970 334046 349026 334102
rect 349094 334046 349150 334102
rect 349218 334046 349274 334102
rect 349342 334046 349398 334102
rect 348970 333922 349026 333978
rect 349094 333922 349150 333978
rect 349218 333922 349274 333978
rect 349342 333922 349398 333978
rect 348970 316294 349026 316350
rect 349094 316294 349150 316350
rect 349218 316294 349274 316350
rect 349342 316294 349398 316350
rect 348970 316170 349026 316226
rect 349094 316170 349150 316226
rect 349218 316170 349274 316226
rect 349342 316170 349398 316226
rect 348970 316046 349026 316102
rect 349094 316046 349150 316102
rect 349218 316046 349274 316102
rect 349342 316046 349398 316102
rect 348970 315922 349026 315978
rect 349094 315922 349150 315978
rect 349218 315922 349274 315978
rect 349342 315922 349398 315978
rect 348970 298294 349026 298350
rect 349094 298294 349150 298350
rect 349218 298294 349274 298350
rect 349342 298294 349398 298350
rect 348970 298170 349026 298226
rect 349094 298170 349150 298226
rect 349218 298170 349274 298226
rect 349342 298170 349398 298226
rect 348970 298046 349026 298102
rect 349094 298046 349150 298102
rect 349218 298046 349274 298102
rect 349342 298046 349398 298102
rect 348970 297922 349026 297978
rect 349094 297922 349150 297978
rect 349218 297922 349274 297978
rect 349342 297922 349398 297978
rect 348970 280294 349026 280350
rect 349094 280294 349150 280350
rect 349218 280294 349274 280350
rect 349342 280294 349398 280350
rect 348970 280170 349026 280226
rect 349094 280170 349150 280226
rect 349218 280170 349274 280226
rect 349342 280170 349398 280226
rect 348970 280046 349026 280102
rect 349094 280046 349150 280102
rect 349218 280046 349274 280102
rect 349342 280046 349398 280102
rect 348970 279922 349026 279978
rect 349094 279922 349150 279978
rect 349218 279922 349274 279978
rect 349342 279922 349398 279978
rect 348970 262294 349026 262350
rect 349094 262294 349150 262350
rect 349218 262294 349274 262350
rect 349342 262294 349398 262350
rect 348970 262170 349026 262226
rect 349094 262170 349150 262226
rect 349218 262170 349274 262226
rect 349342 262170 349398 262226
rect 348970 262046 349026 262102
rect 349094 262046 349150 262102
rect 349218 262046 349274 262102
rect 349342 262046 349398 262102
rect 348970 261922 349026 261978
rect 349094 261922 349150 261978
rect 349218 261922 349274 261978
rect 349342 261922 349398 261978
rect 348970 244294 349026 244350
rect 349094 244294 349150 244350
rect 349218 244294 349274 244350
rect 349342 244294 349398 244350
rect 348970 244170 349026 244226
rect 349094 244170 349150 244226
rect 349218 244170 349274 244226
rect 349342 244170 349398 244226
rect 348970 244046 349026 244102
rect 349094 244046 349150 244102
rect 349218 244046 349274 244102
rect 349342 244046 349398 244102
rect 348970 243922 349026 243978
rect 349094 243922 349150 243978
rect 349218 243922 349274 243978
rect 349342 243922 349398 243978
rect 330970 226294 331026 226350
rect 331094 226294 331150 226350
rect 331218 226294 331274 226350
rect 331342 226294 331398 226350
rect 330970 226170 331026 226226
rect 331094 226170 331150 226226
rect 331218 226170 331274 226226
rect 331342 226170 331398 226226
rect 330970 226046 331026 226102
rect 331094 226046 331150 226102
rect 331218 226046 331274 226102
rect 331342 226046 331398 226102
rect 330970 225922 331026 225978
rect 331094 225922 331150 225978
rect 331218 225922 331274 225978
rect 331342 225922 331398 225978
rect 330970 208294 331026 208350
rect 331094 208294 331150 208350
rect 331218 208294 331274 208350
rect 331342 208294 331398 208350
rect 330970 208170 331026 208226
rect 331094 208170 331150 208226
rect 331218 208170 331274 208226
rect 331342 208170 331398 208226
rect 330970 208046 331026 208102
rect 331094 208046 331150 208102
rect 331218 208046 331274 208102
rect 331342 208046 331398 208102
rect 330970 207922 331026 207978
rect 331094 207922 331150 207978
rect 331218 207922 331274 207978
rect 331342 207922 331398 207978
rect 330970 190294 331026 190350
rect 331094 190294 331150 190350
rect 331218 190294 331274 190350
rect 331342 190294 331398 190350
rect 330970 190170 331026 190226
rect 331094 190170 331150 190226
rect 331218 190170 331274 190226
rect 331342 190170 331398 190226
rect 330970 190046 331026 190102
rect 331094 190046 331150 190102
rect 331218 190046 331274 190102
rect 331342 190046 331398 190102
rect 330970 189922 331026 189978
rect 331094 189922 331150 189978
rect 331218 189922 331274 189978
rect 331342 189922 331398 189978
rect 330970 172294 331026 172350
rect 331094 172294 331150 172350
rect 331218 172294 331274 172350
rect 331342 172294 331398 172350
rect 330970 172170 331026 172226
rect 331094 172170 331150 172226
rect 331218 172170 331274 172226
rect 331342 172170 331398 172226
rect 330970 172046 331026 172102
rect 331094 172046 331150 172102
rect 331218 172046 331274 172102
rect 331342 172046 331398 172102
rect 330970 171922 331026 171978
rect 331094 171922 331150 171978
rect 331218 171922 331274 171978
rect 331342 171922 331398 171978
rect 330970 154294 331026 154350
rect 331094 154294 331150 154350
rect 331218 154294 331274 154350
rect 331342 154294 331398 154350
rect 330970 154170 331026 154226
rect 331094 154170 331150 154226
rect 331218 154170 331274 154226
rect 331342 154170 331398 154226
rect 330970 154046 331026 154102
rect 331094 154046 331150 154102
rect 331218 154046 331274 154102
rect 331342 154046 331398 154102
rect 330970 153922 331026 153978
rect 331094 153922 331150 153978
rect 331218 153922 331274 153978
rect 331342 153922 331398 153978
rect 330970 136294 331026 136350
rect 331094 136294 331150 136350
rect 331218 136294 331274 136350
rect 331342 136294 331398 136350
rect 330970 136170 331026 136226
rect 331094 136170 331150 136226
rect 331218 136170 331274 136226
rect 331342 136170 331398 136226
rect 330970 136046 331026 136102
rect 331094 136046 331150 136102
rect 331218 136046 331274 136102
rect 331342 136046 331398 136102
rect 330970 135922 331026 135978
rect 331094 135922 331150 135978
rect 331218 135922 331274 135978
rect 331342 135922 331398 135978
rect 330970 118294 331026 118350
rect 331094 118294 331150 118350
rect 331218 118294 331274 118350
rect 331342 118294 331398 118350
rect 330970 118170 331026 118226
rect 331094 118170 331150 118226
rect 331218 118170 331274 118226
rect 331342 118170 331398 118226
rect 330970 118046 331026 118102
rect 331094 118046 331150 118102
rect 331218 118046 331274 118102
rect 331342 118046 331398 118102
rect 330970 117922 331026 117978
rect 331094 117922 331150 117978
rect 331218 117922 331274 117978
rect 331342 117922 331398 117978
rect 330970 100294 331026 100350
rect 331094 100294 331150 100350
rect 331218 100294 331274 100350
rect 331342 100294 331398 100350
rect 330970 100170 331026 100226
rect 331094 100170 331150 100226
rect 331218 100170 331274 100226
rect 331342 100170 331398 100226
rect 330970 100046 331026 100102
rect 331094 100046 331150 100102
rect 331218 100046 331274 100102
rect 331342 100046 331398 100102
rect 330970 99922 331026 99978
rect 331094 99922 331150 99978
rect 331218 99922 331274 99978
rect 331342 99922 331398 99978
rect 330970 82294 331026 82350
rect 331094 82294 331150 82350
rect 331218 82294 331274 82350
rect 331342 82294 331398 82350
rect 330970 82170 331026 82226
rect 331094 82170 331150 82226
rect 331218 82170 331274 82226
rect 331342 82170 331398 82226
rect 330970 82046 331026 82102
rect 331094 82046 331150 82102
rect 331218 82046 331274 82102
rect 331342 82046 331398 82102
rect 330970 81922 331026 81978
rect 331094 81922 331150 81978
rect 331218 81922 331274 81978
rect 331342 81922 331398 81978
rect 330970 64294 331026 64350
rect 331094 64294 331150 64350
rect 331218 64294 331274 64350
rect 331342 64294 331398 64350
rect 330970 64170 331026 64226
rect 331094 64170 331150 64226
rect 331218 64170 331274 64226
rect 331342 64170 331398 64226
rect 330970 64046 331026 64102
rect 331094 64046 331150 64102
rect 331218 64046 331274 64102
rect 331342 64046 331398 64102
rect 330970 63922 331026 63978
rect 331094 63922 331150 63978
rect 331218 63922 331274 63978
rect 331342 63922 331398 63978
rect 345250 238294 345306 238350
rect 345374 238294 345430 238350
rect 345498 238294 345554 238350
rect 345622 238294 345678 238350
rect 345250 238170 345306 238226
rect 345374 238170 345430 238226
rect 345498 238170 345554 238226
rect 345622 238170 345678 238226
rect 345250 238046 345306 238102
rect 345374 238046 345430 238102
rect 345498 238046 345554 238102
rect 345622 238046 345678 238102
rect 345250 237922 345306 237978
rect 345374 237922 345430 237978
rect 345498 237922 345554 237978
rect 345622 237922 345678 237978
rect 345250 220294 345306 220350
rect 345374 220294 345430 220350
rect 345498 220294 345554 220350
rect 345622 220294 345678 220350
rect 345250 220170 345306 220226
rect 345374 220170 345430 220226
rect 345498 220170 345554 220226
rect 345622 220170 345678 220226
rect 345250 220046 345306 220102
rect 345374 220046 345430 220102
rect 345498 220046 345554 220102
rect 345622 220046 345678 220102
rect 345250 219922 345306 219978
rect 345374 219922 345430 219978
rect 345498 219922 345554 219978
rect 345622 219922 345678 219978
rect 345250 202294 345306 202350
rect 345374 202294 345430 202350
rect 345498 202294 345554 202350
rect 345622 202294 345678 202350
rect 345250 202170 345306 202226
rect 345374 202170 345430 202226
rect 345498 202170 345554 202226
rect 345622 202170 345678 202226
rect 345250 202046 345306 202102
rect 345374 202046 345430 202102
rect 345498 202046 345554 202102
rect 345622 202046 345678 202102
rect 345250 201922 345306 201978
rect 345374 201922 345430 201978
rect 345498 201922 345554 201978
rect 345622 201922 345678 201978
rect 345250 184294 345306 184350
rect 345374 184294 345430 184350
rect 345498 184294 345554 184350
rect 345622 184294 345678 184350
rect 345250 184170 345306 184226
rect 345374 184170 345430 184226
rect 345498 184170 345554 184226
rect 345622 184170 345678 184226
rect 345250 184046 345306 184102
rect 345374 184046 345430 184102
rect 345498 184046 345554 184102
rect 345622 184046 345678 184102
rect 345250 183922 345306 183978
rect 345374 183922 345430 183978
rect 345498 183922 345554 183978
rect 345622 183922 345678 183978
rect 348970 226294 349026 226350
rect 349094 226294 349150 226350
rect 349218 226294 349274 226350
rect 349342 226294 349398 226350
rect 348970 226170 349026 226226
rect 349094 226170 349150 226226
rect 349218 226170 349274 226226
rect 349342 226170 349398 226226
rect 348970 226046 349026 226102
rect 349094 226046 349150 226102
rect 349218 226046 349274 226102
rect 349342 226046 349398 226102
rect 348970 225922 349026 225978
rect 349094 225922 349150 225978
rect 349218 225922 349274 225978
rect 349342 225922 349398 225978
rect 363250 597156 363306 597212
rect 363374 597156 363430 597212
rect 363498 597156 363554 597212
rect 363622 597156 363678 597212
rect 363250 597032 363306 597088
rect 363374 597032 363430 597088
rect 363498 597032 363554 597088
rect 363622 597032 363678 597088
rect 363250 596908 363306 596964
rect 363374 596908 363430 596964
rect 363498 596908 363554 596964
rect 363622 596908 363678 596964
rect 363250 596784 363306 596840
rect 363374 596784 363430 596840
rect 363498 596784 363554 596840
rect 363622 596784 363678 596840
rect 363250 580294 363306 580350
rect 363374 580294 363430 580350
rect 363498 580294 363554 580350
rect 363622 580294 363678 580350
rect 363250 580170 363306 580226
rect 363374 580170 363430 580226
rect 363498 580170 363554 580226
rect 363622 580170 363678 580226
rect 363250 580046 363306 580102
rect 363374 580046 363430 580102
rect 363498 580046 363554 580102
rect 363622 580046 363678 580102
rect 363250 579922 363306 579978
rect 363374 579922 363430 579978
rect 363498 579922 363554 579978
rect 363622 579922 363678 579978
rect 363250 562294 363306 562350
rect 363374 562294 363430 562350
rect 363498 562294 363554 562350
rect 363622 562294 363678 562350
rect 363250 562170 363306 562226
rect 363374 562170 363430 562226
rect 363498 562170 363554 562226
rect 363622 562170 363678 562226
rect 363250 562046 363306 562102
rect 363374 562046 363430 562102
rect 363498 562046 363554 562102
rect 363622 562046 363678 562102
rect 363250 561922 363306 561978
rect 363374 561922 363430 561978
rect 363498 561922 363554 561978
rect 363622 561922 363678 561978
rect 363250 544294 363306 544350
rect 363374 544294 363430 544350
rect 363498 544294 363554 544350
rect 363622 544294 363678 544350
rect 363250 544170 363306 544226
rect 363374 544170 363430 544226
rect 363498 544170 363554 544226
rect 363622 544170 363678 544226
rect 363250 544046 363306 544102
rect 363374 544046 363430 544102
rect 363498 544046 363554 544102
rect 363622 544046 363678 544102
rect 363250 543922 363306 543978
rect 363374 543922 363430 543978
rect 363498 543922 363554 543978
rect 363622 543922 363678 543978
rect 363250 526294 363306 526350
rect 363374 526294 363430 526350
rect 363498 526294 363554 526350
rect 363622 526294 363678 526350
rect 363250 526170 363306 526226
rect 363374 526170 363430 526226
rect 363498 526170 363554 526226
rect 363622 526170 363678 526226
rect 363250 526046 363306 526102
rect 363374 526046 363430 526102
rect 363498 526046 363554 526102
rect 363622 526046 363678 526102
rect 363250 525922 363306 525978
rect 363374 525922 363430 525978
rect 363498 525922 363554 525978
rect 363622 525922 363678 525978
rect 363250 508294 363306 508350
rect 363374 508294 363430 508350
rect 363498 508294 363554 508350
rect 363622 508294 363678 508350
rect 363250 508170 363306 508226
rect 363374 508170 363430 508226
rect 363498 508170 363554 508226
rect 363622 508170 363678 508226
rect 363250 508046 363306 508102
rect 363374 508046 363430 508102
rect 363498 508046 363554 508102
rect 363622 508046 363678 508102
rect 363250 507922 363306 507978
rect 363374 507922 363430 507978
rect 363498 507922 363554 507978
rect 363622 507922 363678 507978
rect 363250 490294 363306 490350
rect 363374 490294 363430 490350
rect 363498 490294 363554 490350
rect 363622 490294 363678 490350
rect 363250 490170 363306 490226
rect 363374 490170 363430 490226
rect 363498 490170 363554 490226
rect 363622 490170 363678 490226
rect 363250 490046 363306 490102
rect 363374 490046 363430 490102
rect 363498 490046 363554 490102
rect 363622 490046 363678 490102
rect 363250 489922 363306 489978
rect 363374 489922 363430 489978
rect 363498 489922 363554 489978
rect 363622 489922 363678 489978
rect 363250 472294 363306 472350
rect 363374 472294 363430 472350
rect 363498 472294 363554 472350
rect 363622 472294 363678 472350
rect 363250 472170 363306 472226
rect 363374 472170 363430 472226
rect 363498 472170 363554 472226
rect 363622 472170 363678 472226
rect 363250 472046 363306 472102
rect 363374 472046 363430 472102
rect 363498 472046 363554 472102
rect 363622 472046 363678 472102
rect 363250 471922 363306 471978
rect 363374 471922 363430 471978
rect 363498 471922 363554 471978
rect 363622 471922 363678 471978
rect 363250 454294 363306 454350
rect 363374 454294 363430 454350
rect 363498 454294 363554 454350
rect 363622 454294 363678 454350
rect 363250 454170 363306 454226
rect 363374 454170 363430 454226
rect 363498 454170 363554 454226
rect 363622 454170 363678 454226
rect 363250 454046 363306 454102
rect 363374 454046 363430 454102
rect 363498 454046 363554 454102
rect 363622 454046 363678 454102
rect 363250 453922 363306 453978
rect 363374 453922 363430 453978
rect 363498 453922 363554 453978
rect 363622 453922 363678 453978
rect 363250 436294 363306 436350
rect 363374 436294 363430 436350
rect 363498 436294 363554 436350
rect 363622 436294 363678 436350
rect 363250 436170 363306 436226
rect 363374 436170 363430 436226
rect 363498 436170 363554 436226
rect 363622 436170 363678 436226
rect 363250 436046 363306 436102
rect 363374 436046 363430 436102
rect 363498 436046 363554 436102
rect 363622 436046 363678 436102
rect 363250 435922 363306 435978
rect 363374 435922 363430 435978
rect 363498 435922 363554 435978
rect 363622 435922 363678 435978
rect 363250 418294 363306 418350
rect 363374 418294 363430 418350
rect 363498 418294 363554 418350
rect 363622 418294 363678 418350
rect 363250 418170 363306 418226
rect 363374 418170 363430 418226
rect 363498 418170 363554 418226
rect 363622 418170 363678 418226
rect 363250 418046 363306 418102
rect 363374 418046 363430 418102
rect 363498 418046 363554 418102
rect 363622 418046 363678 418102
rect 363250 417922 363306 417978
rect 363374 417922 363430 417978
rect 363498 417922 363554 417978
rect 363622 417922 363678 417978
rect 363250 400294 363306 400350
rect 363374 400294 363430 400350
rect 363498 400294 363554 400350
rect 363622 400294 363678 400350
rect 363250 400170 363306 400226
rect 363374 400170 363430 400226
rect 363498 400170 363554 400226
rect 363622 400170 363678 400226
rect 363250 400046 363306 400102
rect 363374 400046 363430 400102
rect 363498 400046 363554 400102
rect 363622 400046 363678 400102
rect 363250 399922 363306 399978
rect 363374 399922 363430 399978
rect 363498 399922 363554 399978
rect 363622 399922 363678 399978
rect 363250 382294 363306 382350
rect 363374 382294 363430 382350
rect 363498 382294 363554 382350
rect 363622 382294 363678 382350
rect 363250 382170 363306 382226
rect 363374 382170 363430 382226
rect 363498 382170 363554 382226
rect 363622 382170 363678 382226
rect 363250 382046 363306 382102
rect 363374 382046 363430 382102
rect 363498 382046 363554 382102
rect 363622 382046 363678 382102
rect 363250 381922 363306 381978
rect 363374 381922 363430 381978
rect 363498 381922 363554 381978
rect 363622 381922 363678 381978
rect 363250 364294 363306 364350
rect 363374 364294 363430 364350
rect 363498 364294 363554 364350
rect 363622 364294 363678 364350
rect 363250 364170 363306 364226
rect 363374 364170 363430 364226
rect 363498 364170 363554 364226
rect 363622 364170 363678 364226
rect 363250 364046 363306 364102
rect 363374 364046 363430 364102
rect 363498 364046 363554 364102
rect 363622 364046 363678 364102
rect 363250 363922 363306 363978
rect 363374 363922 363430 363978
rect 363498 363922 363554 363978
rect 363622 363922 363678 363978
rect 363250 346294 363306 346350
rect 363374 346294 363430 346350
rect 363498 346294 363554 346350
rect 363622 346294 363678 346350
rect 363250 346170 363306 346226
rect 363374 346170 363430 346226
rect 363498 346170 363554 346226
rect 363622 346170 363678 346226
rect 363250 346046 363306 346102
rect 363374 346046 363430 346102
rect 363498 346046 363554 346102
rect 363622 346046 363678 346102
rect 363250 345922 363306 345978
rect 363374 345922 363430 345978
rect 363498 345922 363554 345978
rect 363622 345922 363678 345978
rect 363250 328294 363306 328350
rect 363374 328294 363430 328350
rect 363498 328294 363554 328350
rect 363622 328294 363678 328350
rect 363250 328170 363306 328226
rect 363374 328170 363430 328226
rect 363498 328170 363554 328226
rect 363622 328170 363678 328226
rect 363250 328046 363306 328102
rect 363374 328046 363430 328102
rect 363498 328046 363554 328102
rect 363622 328046 363678 328102
rect 363250 327922 363306 327978
rect 363374 327922 363430 327978
rect 363498 327922 363554 327978
rect 363622 327922 363678 327978
rect 363250 310294 363306 310350
rect 363374 310294 363430 310350
rect 363498 310294 363554 310350
rect 363622 310294 363678 310350
rect 363250 310170 363306 310226
rect 363374 310170 363430 310226
rect 363498 310170 363554 310226
rect 363622 310170 363678 310226
rect 363250 310046 363306 310102
rect 363374 310046 363430 310102
rect 363498 310046 363554 310102
rect 363622 310046 363678 310102
rect 363250 309922 363306 309978
rect 363374 309922 363430 309978
rect 363498 309922 363554 309978
rect 363622 309922 363678 309978
rect 363250 292294 363306 292350
rect 363374 292294 363430 292350
rect 363498 292294 363554 292350
rect 363622 292294 363678 292350
rect 363250 292170 363306 292226
rect 363374 292170 363430 292226
rect 363498 292170 363554 292226
rect 363622 292170 363678 292226
rect 363250 292046 363306 292102
rect 363374 292046 363430 292102
rect 363498 292046 363554 292102
rect 363622 292046 363678 292102
rect 363250 291922 363306 291978
rect 363374 291922 363430 291978
rect 363498 291922 363554 291978
rect 363622 291922 363678 291978
rect 363250 274294 363306 274350
rect 363374 274294 363430 274350
rect 363498 274294 363554 274350
rect 363622 274294 363678 274350
rect 363250 274170 363306 274226
rect 363374 274170 363430 274226
rect 363498 274170 363554 274226
rect 363622 274170 363678 274226
rect 363250 274046 363306 274102
rect 363374 274046 363430 274102
rect 363498 274046 363554 274102
rect 363622 274046 363678 274102
rect 363250 273922 363306 273978
rect 363374 273922 363430 273978
rect 363498 273922 363554 273978
rect 363622 273922 363678 273978
rect 363250 256294 363306 256350
rect 363374 256294 363430 256350
rect 363498 256294 363554 256350
rect 363622 256294 363678 256350
rect 363250 256170 363306 256226
rect 363374 256170 363430 256226
rect 363498 256170 363554 256226
rect 363622 256170 363678 256226
rect 363250 256046 363306 256102
rect 363374 256046 363430 256102
rect 363498 256046 363554 256102
rect 363622 256046 363678 256102
rect 363250 255922 363306 255978
rect 363374 255922 363430 255978
rect 363498 255922 363554 255978
rect 363622 255922 363678 255978
rect 363250 238294 363306 238350
rect 363374 238294 363430 238350
rect 363498 238294 363554 238350
rect 363622 238294 363678 238350
rect 363250 238170 363306 238226
rect 363374 238170 363430 238226
rect 363498 238170 363554 238226
rect 363622 238170 363678 238226
rect 363250 238046 363306 238102
rect 363374 238046 363430 238102
rect 363498 238046 363554 238102
rect 363622 238046 363678 238102
rect 363250 237922 363306 237978
rect 363374 237922 363430 237978
rect 363498 237922 363554 237978
rect 363622 237922 363678 237978
rect 363250 220294 363306 220350
rect 363374 220294 363430 220350
rect 363498 220294 363554 220350
rect 363622 220294 363678 220350
rect 363250 220170 363306 220226
rect 363374 220170 363430 220226
rect 363498 220170 363554 220226
rect 363622 220170 363678 220226
rect 363250 220046 363306 220102
rect 363374 220046 363430 220102
rect 363498 220046 363554 220102
rect 363622 220046 363678 220102
rect 363250 219922 363306 219978
rect 363374 219922 363430 219978
rect 363498 219922 363554 219978
rect 363622 219922 363678 219978
rect 366970 598116 367026 598172
rect 367094 598116 367150 598172
rect 367218 598116 367274 598172
rect 367342 598116 367398 598172
rect 366970 597992 367026 598048
rect 367094 597992 367150 598048
rect 367218 597992 367274 598048
rect 367342 597992 367398 598048
rect 366970 597868 367026 597924
rect 367094 597868 367150 597924
rect 367218 597868 367274 597924
rect 367342 597868 367398 597924
rect 366970 597744 367026 597800
rect 367094 597744 367150 597800
rect 367218 597744 367274 597800
rect 367342 597744 367398 597800
rect 366970 586294 367026 586350
rect 367094 586294 367150 586350
rect 367218 586294 367274 586350
rect 367342 586294 367398 586350
rect 366970 586170 367026 586226
rect 367094 586170 367150 586226
rect 367218 586170 367274 586226
rect 367342 586170 367398 586226
rect 366970 586046 367026 586102
rect 367094 586046 367150 586102
rect 367218 586046 367274 586102
rect 367342 586046 367398 586102
rect 366970 585922 367026 585978
rect 367094 585922 367150 585978
rect 367218 585922 367274 585978
rect 367342 585922 367398 585978
rect 366970 568294 367026 568350
rect 367094 568294 367150 568350
rect 367218 568294 367274 568350
rect 367342 568294 367398 568350
rect 366970 568170 367026 568226
rect 367094 568170 367150 568226
rect 367218 568170 367274 568226
rect 367342 568170 367398 568226
rect 366970 568046 367026 568102
rect 367094 568046 367150 568102
rect 367218 568046 367274 568102
rect 367342 568046 367398 568102
rect 366970 567922 367026 567978
rect 367094 567922 367150 567978
rect 367218 567922 367274 567978
rect 367342 567922 367398 567978
rect 366970 550294 367026 550350
rect 367094 550294 367150 550350
rect 367218 550294 367274 550350
rect 367342 550294 367398 550350
rect 366970 550170 367026 550226
rect 367094 550170 367150 550226
rect 367218 550170 367274 550226
rect 367342 550170 367398 550226
rect 366970 550046 367026 550102
rect 367094 550046 367150 550102
rect 367218 550046 367274 550102
rect 367342 550046 367398 550102
rect 366970 549922 367026 549978
rect 367094 549922 367150 549978
rect 367218 549922 367274 549978
rect 367342 549922 367398 549978
rect 366970 532294 367026 532350
rect 367094 532294 367150 532350
rect 367218 532294 367274 532350
rect 367342 532294 367398 532350
rect 366970 532170 367026 532226
rect 367094 532170 367150 532226
rect 367218 532170 367274 532226
rect 367342 532170 367398 532226
rect 366970 532046 367026 532102
rect 367094 532046 367150 532102
rect 367218 532046 367274 532102
rect 367342 532046 367398 532102
rect 366970 531922 367026 531978
rect 367094 531922 367150 531978
rect 367218 531922 367274 531978
rect 367342 531922 367398 531978
rect 366970 514294 367026 514350
rect 367094 514294 367150 514350
rect 367218 514294 367274 514350
rect 367342 514294 367398 514350
rect 366970 514170 367026 514226
rect 367094 514170 367150 514226
rect 367218 514170 367274 514226
rect 367342 514170 367398 514226
rect 366970 514046 367026 514102
rect 367094 514046 367150 514102
rect 367218 514046 367274 514102
rect 367342 514046 367398 514102
rect 366970 513922 367026 513978
rect 367094 513922 367150 513978
rect 367218 513922 367274 513978
rect 367342 513922 367398 513978
rect 366970 496294 367026 496350
rect 367094 496294 367150 496350
rect 367218 496294 367274 496350
rect 367342 496294 367398 496350
rect 366970 496170 367026 496226
rect 367094 496170 367150 496226
rect 367218 496170 367274 496226
rect 367342 496170 367398 496226
rect 366970 496046 367026 496102
rect 367094 496046 367150 496102
rect 367218 496046 367274 496102
rect 367342 496046 367398 496102
rect 366970 495922 367026 495978
rect 367094 495922 367150 495978
rect 367218 495922 367274 495978
rect 367342 495922 367398 495978
rect 366970 478294 367026 478350
rect 367094 478294 367150 478350
rect 367218 478294 367274 478350
rect 367342 478294 367398 478350
rect 366970 478170 367026 478226
rect 367094 478170 367150 478226
rect 367218 478170 367274 478226
rect 367342 478170 367398 478226
rect 366970 478046 367026 478102
rect 367094 478046 367150 478102
rect 367218 478046 367274 478102
rect 367342 478046 367398 478102
rect 366970 477922 367026 477978
rect 367094 477922 367150 477978
rect 367218 477922 367274 477978
rect 367342 477922 367398 477978
rect 366970 460294 367026 460350
rect 367094 460294 367150 460350
rect 367218 460294 367274 460350
rect 367342 460294 367398 460350
rect 366970 460170 367026 460226
rect 367094 460170 367150 460226
rect 367218 460170 367274 460226
rect 367342 460170 367398 460226
rect 366970 460046 367026 460102
rect 367094 460046 367150 460102
rect 367218 460046 367274 460102
rect 367342 460046 367398 460102
rect 366970 459922 367026 459978
rect 367094 459922 367150 459978
rect 367218 459922 367274 459978
rect 367342 459922 367398 459978
rect 366970 442294 367026 442350
rect 367094 442294 367150 442350
rect 367218 442294 367274 442350
rect 367342 442294 367398 442350
rect 366970 442170 367026 442226
rect 367094 442170 367150 442226
rect 367218 442170 367274 442226
rect 367342 442170 367398 442226
rect 366970 442046 367026 442102
rect 367094 442046 367150 442102
rect 367218 442046 367274 442102
rect 367342 442046 367398 442102
rect 366970 441922 367026 441978
rect 367094 441922 367150 441978
rect 367218 441922 367274 441978
rect 367342 441922 367398 441978
rect 366970 424294 367026 424350
rect 367094 424294 367150 424350
rect 367218 424294 367274 424350
rect 367342 424294 367398 424350
rect 366970 424170 367026 424226
rect 367094 424170 367150 424226
rect 367218 424170 367274 424226
rect 367342 424170 367398 424226
rect 366970 424046 367026 424102
rect 367094 424046 367150 424102
rect 367218 424046 367274 424102
rect 367342 424046 367398 424102
rect 366970 423922 367026 423978
rect 367094 423922 367150 423978
rect 367218 423922 367274 423978
rect 367342 423922 367398 423978
rect 366970 406294 367026 406350
rect 367094 406294 367150 406350
rect 367218 406294 367274 406350
rect 367342 406294 367398 406350
rect 366970 406170 367026 406226
rect 367094 406170 367150 406226
rect 367218 406170 367274 406226
rect 367342 406170 367398 406226
rect 366970 406046 367026 406102
rect 367094 406046 367150 406102
rect 367218 406046 367274 406102
rect 367342 406046 367398 406102
rect 366970 405922 367026 405978
rect 367094 405922 367150 405978
rect 367218 405922 367274 405978
rect 367342 405922 367398 405978
rect 366970 388294 367026 388350
rect 367094 388294 367150 388350
rect 367218 388294 367274 388350
rect 367342 388294 367398 388350
rect 366970 388170 367026 388226
rect 367094 388170 367150 388226
rect 367218 388170 367274 388226
rect 367342 388170 367398 388226
rect 366970 388046 367026 388102
rect 367094 388046 367150 388102
rect 367218 388046 367274 388102
rect 367342 388046 367398 388102
rect 366970 387922 367026 387978
rect 367094 387922 367150 387978
rect 367218 387922 367274 387978
rect 367342 387922 367398 387978
rect 366970 370294 367026 370350
rect 367094 370294 367150 370350
rect 367218 370294 367274 370350
rect 367342 370294 367398 370350
rect 366970 370170 367026 370226
rect 367094 370170 367150 370226
rect 367218 370170 367274 370226
rect 367342 370170 367398 370226
rect 366970 370046 367026 370102
rect 367094 370046 367150 370102
rect 367218 370046 367274 370102
rect 367342 370046 367398 370102
rect 366970 369922 367026 369978
rect 367094 369922 367150 369978
rect 367218 369922 367274 369978
rect 367342 369922 367398 369978
rect 366970 352294 367026 352350
rect 367094 352294 367150 352350
rect 367218 352294 367274 352350
rect 367342 352294 367398 352350
rect 366970 352170 367026 352226
rect 367094 352170 367150 352226
rect 367218 352170 367274 352226
rect 367342 352170 367398 352226
rect 366970 352046 367026 352102
rect 367094 352046 367150 352102
rect 367218 352046 367274 352102
rect 367342 352046 367398 352102
rect 366970 351922 367026 351978
rect 367094 351922 367150 351978
rect 367218 351922 367274 351978
rect 367342 351922 367398 351978
rect 366970 334294 367026 334350
rect 367094 334294 367150 334350
rect 367218 334294 367274 334350
rect 367342 334294 367398 334350
rect 366970 334170 367026 334226
rect 367094 334170 367150 334226
rect 367218 334170 367274 334226
rect 367342 334170 367398 334226
rect 366970 334046 367026 334102
rect 367094 334046 367150 334102
rect 367218 334046 367274 334102
rect 367342 334046 367398 334102
rect 366970 333922 367026 333978
rect 367094 333922 367150 333978
rect 367218 333922 367274 333978
rect 367342 333922 367398 333978
rect 366970 316294 367026 316350
rect 367094 316294 367150 316350
rect 367218 316294 367274 316350
rect 367342 316294 367398 316350
rect 366970 316170 367026 316226
rect 367094 316170 367150 316226
rect 367218 316170 367274 316226
rect 367342 316170 367398 316226
rect 366970 316046 367026 316102
rect 367094 316046 367150 316102
rect 367218 316046 367274 316102
rect 367342 316046 367398 316102
rect 366970 315922 367026 315978
rect 367094 315922 367150 315978
rect 367218 315922 367274 315978
rect 367342 315922 367398 315978
rect 366970 298294 367026 298350
rect 367094 298294 367150 298350
rect 367218 298294 367274 298350
rect 367342 298294 367398 298350
rect 366970 298170 367026 298226
rect 367094 298170 367150 298226
rect 367218 298170 367274 298226
rect 367342 298170 367398 298226
rect 366970 298046 367026 298102
rect 367094 298046 367150 298102
rect 367218 298046 367274 298102
rect 367342 298046 367398 298102
rect 366970 297922 367026 297978
rect 367094 297922 367150 297978
rect 367218 297922 367274 297978
rect 367342 297922 367398 297978
rect 366970 280294 367026 280350
rect 367094 280294 367150 280350
rect 367218 280294 367274 280350
rect 367342 280294 367398 280350
rect 366970 280170 367026 280226
rect 367094 280170 367150 280226
rect 367218 280170 367274 280226
rect 367342 280170 367398 280226
rect 366970 280046 367026 280102
rect 367094 280046 367150 280102
rect 367218 280046 367274 280102
rect 367342 280046 367398 280102
rect 366970 279922 367026 279978
rect 367094 279922 367150 279978
rect 367218 279922 367274 279978
rect 367342 279922 367398 279978
rect 366970 262294 367026 262350
rect 367094 262294 367150 262350
rect 367218 262294 367274 262350
rect 367342 262294 367398 262350
rect 366970 262170 367026 262226
rect 367094 262170 367150 262226
rect 367218 262170 367274 262226
rect 367342 262170 367398 262226
rect 366970 262046 367026 262102
rect 367094 262046 367150 262102
rect 367218 262046 367274 262102
rect 367342 262046 367398 262102
rect 366970 261922 367026 261978
rect 367094 261922 367150 261978
rect 367218 261922 367274 261978
rect 367342 261922 367398 261978
rect 366970 244294 367026 244350
rect 367094 244294 367150 244350
rect 367218 244294 367274 244350
rect 367342 244294 367398 244350
rect 366970 244170 367026 244226
rect 367094 244170 367150 244226
rect 367218 244170 367274 244226
rect 367342 244170 367398 244226
rect 366970 244046 367026 244102
rect 367094 244046 367150 244102
rect 367218 244046 367274 244102
rect 367342 244046 367398 244102
rect 366970 243922 367026 243978
rect 367094 243922 367150 243978
rect 367218 243922 367274 243978
rect 367342 243922 367398 243978
rect 366970 226294 367026 226350
rect 367094 226294 367150 226350
rect 367218 226294 367274 226350
rect 367342 226294 367398 226350
rect 366970 226170 367026 226226
rect 367094 226170 367150 226226
rect 367218 226170 367274 226226
rect 367342 226170 367398 226226
rect 366970 226046 367026 226102
rect 367094 226046 367150 226102
rect 367218 226046 367274 226102
rect 367342 226046 367398 226102
rect 366970 225922 367026 225978
rect 367094 225922 367150 225978
rect 367218 225922 367274 225978
rect 367342 225922 367398 225978
rect 381250 597156 381306 597212
rect 381374 597156 381430 597212
rect 381498 597156 381554 597212
rect 381622 597156 381678 597212
rect 381250 597032 381306 597088
rect 381374 597032 381430 597088
rect 381498 597032 381554 597088
rect 381622 597032 381678 597088
rect 381250 596908 381306 596964
rect 381374 596908 381430 596964
rect 381498 596908 381554 596964
rect 381622 596908 381678 596964
rect 381250 596784 381306 596840
rect 381374 596784 381430 596840
rect 381498 596784 381554 596840
rect 381622 596784 381678 596840
rect 381250 580294 381306 580350
rect 381374 580294 381430 580350
rect 381498 580294 381554 580350
rect 381622 580294 381678 580350
rect 381250 580170 381306 580226
rect 381374 580170 381430 580226
rect 381498 580170 381554 580226
rect 381622 580170 381678 580226
rect 381250 580046 381306 580102
rect 381374 580046 381430 580102
rect 381498 580046 381554 580102
rect 381622 580046 381678 580102
rect 381250 579922 381306 579978
rect 381374 579922 381430 579978
rect 381498 579922 381554 579978
rect 381622 579922 381678 579978
rect 381250 562294 381306 562350
rect 381374 562294 381430 562350
rect 381498 562294 381554 562350
rect 381622 562294 381678 562350
rect 381250 562170 381306 562226
rect 381374 562170 381430 562226
rect 381498 562170 381554 562226
rect 381622 562170 381678 562226
rect 381250 562046 381306 562102
rect 381374 562046 381430 562102
rect 381498 562046 381554 562102
rect 381622 562046 381678 562102
rect 381250 561922 381306 561978
rect 381374 561922 381430 561978
rect 381498 561922 381554 561978
rect 381622 561922 381678 561978
rect 381250 544294 381306 544350
rect 381374 544294 381430 544350
rect 381498 544294 381554 544350
rect 381622 544294 381678 544350
rect 381250 544170 381306 544226
rect 381374 544170 381430 544226
rect 381498 544170 381554 544226
rect 381622 544170 381678 544226
rect 381250 544046 381306 544102
rect 381374 544046 381430 544102
rect 381498 544046 381554 544102
rect 381622 544046 381678 544102
rect 381250 543922 381306 543978
rect 381374 543922 381430 543978
rect 381498 543922 381554 543978
rect 381622 543922 381678 543978
rect 381250 526294 381306 526350
rect 381374 526294 381430 526350
rect 381498 526294 381554 526350
rect 381622 526294 381678 526350
rect 381250 526170 381306 526226
rect 381374 526170 381430 526226
rect 381498 526170 381554 526226
rect 381622 526170 381678 526226
rect 381250 526046 381306 526102
rect 381374 526046 381430 526102
rect 381498 526046 381554 526102
rect 381622 526046 381678 526102
rect 381250 525922 381306 525978
rect 381374 525922 381430 525978
rect 381498 525922 381554 525978
rect 381622 525922 381678 525978
rect 381250 508294 381306 508350
rect 381374 508294 381430 508350
rect 381498 508294 381554 508350
rect 381622 508294 381678 508350
rect 381250 508170 381306 508226
rect 381374 508170 381430 508226
rect 381498 508170 381554 508226
rect 381622 508170 381678 508226
rect 381250 508046 381306 508102
rect 381374 508046 381430 508102
rect 381498 508046 381554 508102
rect 381622 508046 381678 508102
rect 381250 507922 381306 507978
rect 381374 507922 381430 507978
rect 381498 507922 381554 507978
rect 381622 507922 381678 507978
rect 381250 490294 381306 490350
rect 381374 490294 381430 490350
rect 381498 490294 381554 490350
rect 381622 490294 381678 490350
rect 381250 490170 381306 490226
rect 381374 490170 381430 490226
rect 381498 490170 381554 490226
rect 381622 490170 381678 490226
rect 381250 490046 381306 490102
rect 381374 490046 381430 490102
rect 381498 490046 381554 490102
rect 381622 490046 381678 490102
rect 381250 489922 381306 489978
rect 381374 489922 381430 489978
rect 381498 489922 381554 489978
rect 381622 489922 381678 489978
rect 381250 472294 381306 472350
rect 381374 472294 381430 472350
rect 381498 472294 381554 472350
rect 381622 472294 381678 472350
rect 381250 472170 381306 472226
rect 381374 472170 381430 472226
rect 381498 472170 381554 472226
rect 381622 472170 381678 472226
rect 381250 472046 381306 472102
rect 381374 472046 381430 472102
rect 381498 472046 381554 472102
rect 381622 472046 381678 472102
rect 381250 471922 381306 471978
rect 381374 471922 381430 471978
rect 381498 471922 381554 471978
rect 381622 471922 381678 471978
rect 381250 454294 381306 454350
rect 381374 454294 381430 454350
rect 381498 454294 381554 454350
rect 381622 454294 381678 454350
rect 381250 454170 381306 454226
rect 381374 454170 381430 454226
rect 381498 454170 381554 454226
rect 381622 454170 381678 454226
rect 381250 454046 381306 454102
rect 381374 454046 381430 454102
rect 381498 454046 381554 454102
rect 381622 454046 381678 454102
rect 381250 453922 381306 453978
rect 381374 453922 381430 453978
rect 381498 453922 381554 453978
rect 381622 453922 381678 453978
rect 381250 436294 381306 436350
rect 381374 436294 381430 436350
rect 381498 436294 381554 436350
rect 381622 436294 381678 436350
rect 381250 436170 381306 436226
rect 381374 436170 381430 436226
rect 381498 436170 381554 436226
rect 381622 436170 381678 436226
rect 381250 436046 381306 436102
rect 381374 436046 381430 436102
rect 381498 436046 381554 436102
rect 381622 436046 381678 436102
rect 381250 435922 381306 435978
rect 381374 435922 381430 435978
rect 381498 435922 381554 435978
rect 381622 435922 381678 435978
rect 381250 418294 381306 418350
rect 381374 418294 381430 418350
rect 381498 418294 381554 418350
rect 381622 418294 381678 418350
rect 381250 418170 381306 418226
rect 381374 418170 381430 418226
rect 381498 418170 381554 418226
rect 381622 418170 381678 418226
rect 381250 418046 381306 418102
rect 381374 418046 381430 418102
rect 381498 418046 381554 418102
rect 381622 418046 381678 418102
rect 381250 417922 381306 417978
rect 381374 417922 381430 417978
rect 381498 417922 381554 417978
rect 381622 417922 381678 417978
rect 381250 400294 381306 400350
rect 381374 400294 381430 400350
rect 381498 400294 381554 400350
rect 381622 400294 381678 400350
rect 381250 400170 381306 400226
rect 381374 400170 381430 400226
rect 381498 400170 381554 400226
rect 381622 400170 381678 400226
rect 381250 400046 381306 400102
rect 381374 400046 381430 400102
rect 381498 400046 381554 400102
rect 381622 400046 381678 400102
rect 381250 399922 381306 399978
rect 381374 399922 381430 399978
rect 381498 399922 381554 399978
rect 381622 399922 381678 399978
rect 381250 382294 381306 382350
rect 381374 382294 381430 382350
rect 381498 382294 381554 382350
rect 381622 382294 381678 382350
rect 381250 382170 381306 382226
rect 381374 382170 381430 382226
rect 381498 382170 381554 382226
rect 381622 382170 381678 382226
rect 381250 382046 381306 382102
rect 381374 382046 381430 382102
rect 381498 382046 381554 382102
rect 381622 382046 381678 382102
rect 381250 381922 381306 381978
rect 381374 381922 381430 381978
rect 381498 381922 381554 381978
rect 381622 381922 381678 381978
rect 381250 364294 381306 364350
rect 381374 364294 381430 364350
rect 381498 364294 381554 364350
rect 381622 364294 381678 364350
rect 381250 364170 381306 364226
rect 381374 364170 381430 364226
rect 381498 364170 381554 364226
rect 381622 364170 381678 364226
rect 381250 364046 381306 364102
rect 381374 364046 381430 364102
rect 381498 364046 381554 364102
rect 381622 364046 381678 364102
rect 381250 363922 381306 363978
rect 381374 363922 381430 363978
rect 381498 363922 381554 363978
rect 381622 363922 381678 363978
rect 381250 346294 381306 346350
rect 381374 346294 381430 346350
rect 381498 346294 381554 346350
rect 381622 346294 381678 346350
rect 381250 346170 381306 346226
rect 381374 346170 381430 346226
rect 381498 346170 381554 346226
rect 381622 346170 381678 346226
rect 381250 346046 381306 346102
rect 381374 346046 381430 346102
rect 381498 346046 381554 346102
rect 381622 346046 381678 346102
rect 381250 345922 381306 345978
rect 381374 345922 381430 345978
rect 381498 345922 381554 345978
rect 381622 345922 381678 345978
rect 381250 328294 381306 328350
rect 381374 328294 381430 328350
rect 381498 328294 381554 328350
rect 381622 328294 381678 328350
rect 381250 328170 381306 328226
rect 381374 328170 381430 328226
rect 381498 328170 381554 328226
rect 381622 328170 381678 328226
rect 381250 328046 381306 328102
rect 381374 328046 381430 328102
rect 381498 328046 381554 328102
rect 381622 328046 381678 328102
rect 381250 327922 381306 327978
rect 381374 327922 381430 327978
rect 381498 327922 381554 327978
rect 381622 327922 381678 327978
rect 381250 310294 381306 310350
rect 381374 310294 381430 310350
rect 381498 310294 381554 310350
rect 381622 310294 381678 310350
rect 381250 310170 381306 310226
rect 381374 310170 381430 310226
rect 381498 310170 381554 310226
rect 381622 310170 381678 310226
rect 381250 310046 381306 310102
rect 381374 310046 381430 310102
rect 381498 310046 381554 310102
rect 381622 310046 381678 310102
rect 381250 309922 381306 309978
rect 381374 309922 381430 309978
rect 381498 309922 381554 309978
rect 381622 309922 381678 309978
rect 381250 292294 381306 292350
rect 381374 292294 381430 292350
rect 381498 292294 381554 292350
rect 381622 292294 381678 292350
rect 381250 292170 381306 292226
rect 381374 292170 381430 292226
rect 381498 292170 381554 292226
rect 381622 292170 381678 292226
rect 381250 292046 381306 292102
rect 381374 292046 381430 292102
rect 381498 292046 381554 292102
rect 381622 292046 381678 292102
rect 381250 291922 381306 291978
rect 381374 291922 381430 291978
rect 381498 291922 381554 291978
rect 381622 291922 381678 291978
rect 381250 274294 381306 274350
rect 381374 274294 381430 274350
rect 381498 274294 381554 274350
rect 381622 274294 381678 274350
rect 381250 274170 381306 274226
rect 381374 274170 381430 274226
rect 381498 274170 381554 274226
rect 381622 274170 381678 274226
rect 381250 274046 381306 274102
rect 381374 274046 381430 274102
rect 381498 274046 381554 274102
rect 381622 274046 381678 274102
rect 381250 273922 381306 273978
rect 381374 273922 381430 273978
rect 381498 273922 381554 273978
rect 381622 273922 381678 273978
rect 381250 256294 381306 256350
rect 381374 256294 381430 256350
rect 381498 256294 381554 256350
rect 381622 256294 381678 256350
rect 381250 256170 381306 256226
rect 381374 256170 381430 256226
rect 381498 256170 381554 256226
rect 381622 256170 381678 256226
rect 381250 256046 381306 256102
rect 381374 256046 381430 256102
rect 381498 256046 381554 256102
rect 381622 256046 381678 256102
rect 381250 255922 381306 255978
rect 381374 255922 381430 255978
rect 381498 255922 381554 255978
rect 381622 255922 381678 255978
rect 381250 238294 381306 238350
rect 381374 238294 381430 238350
rect 381498 238294 381554 238350
rect 381622 238294 381678 238350
rect 381250 238170 381306 238226
rect 381374 238170 381430 238226
rect 381498 238170 381554 238226
rect 381622 238170 381678 238226
rect 381250 238046 381306 238102
rect 381374 238046 381430 238102
rect 381498 238046 381554 238102
rect 381622 238046 381678 238102
rect 381250 237922 381306 237978
rect 381374 237922 381430 237978
rect 381498 237922 381554 237978
rect 381622 237922 381678 237978
rect 381250 220294 381306 220350
rect 381374 220294 381430 220350
rect 381498 220294 381554 220350
rect 381622 220294 381678 220350
rect 381250 220170 381306 220226
rect 381374 220170 381430 220226
rect 381498 220170 381554 220226
rect 381622 220170 381678 220226
rect 381250 220046 381306 220102
rect 381374 220046 381430 220102
rect 381498 220046 381554 220102
rect 381622 220046 381678 220102
rect 381250 219922 381306 219978
rect 381374 219922 381430 219978
rect 381498 219922 381554 219978
rect 381622 219922 381678 219978
rect 399250 597156 399306 597212
rect 399374 597156 399430 597212
rect 399498 597156 399554 597212
rect 399622 597156 399678 597212
rect 399250 597032 399306 597088
rect 399374 597032 399430 597088
rect 399498 597032 399554 597088
rect 399622 597032 399678 597088
rect 399250 596908 399306 596964
rect 399374 596908 399430 596964
rect 399498 596908 399554 596964
rect 399622 596908 399678 596964
rect 399250 596784 399306 596840
rect 399374 596784 399430 596840
rect 399498 596784 399554 596840
rect 399622 596784 399678 596840
rect 399250 580294 399306 580350
rect 399374 580294 399430 580350
rect 399498 580294 399554 580350
rect 399622 580294 399678 580350
rect 399250 580170 399306 580226
rect 399374 580170 399430 580226
rect 399498 580170 399554 580226
rect 399622 580170 399678 580226
rect 399250 580046 399306 580102
rect 399374 580046 399430 580102
rect 399498 580046 399554 580102
rect 399622 580046 399678 580102
rect 399250 579922 399306 579978
rect 399374 579922 399430 579978
rect 399498 579922 399554 579978
rect 399622 579922 399678 579978
rect 399250 562294 399306 562350
rect 399374 562294 399430 562350
rect 399498 562294 399554 562350
rect 399622 562294 399678 562350
rect 399250 562170 399306 562226
rect 399374 562170 399430 562226
rect 399498 562170 399554 562226
rect 399622 562170 399678 562226
rect 399250 562046 399306 562102
rect 399374 562046 399430 562102
rect 399498 562046 399554 562102
rect 399622 562046 399678 562102
rect 399250 561922 399306 561978
rect 399374 561922 399430 561978
rect 399498 561922 399554 561978
rect 399622 561922 399678 561978
rect 399250 544294 399306 544350
rect 399374 544294 399430 544350
rect 399498 544294 399554 544350
rect 399622 544294 399678 544350
rect 399250 544170 399306 544226
rect 399374 544170 399430 544226
rect 399498 544170 399554 544226
rect 399622 544170 399678 544226
rect 399250 544046 399306 544102
rect 399374 544046 399430 544102
rect 399498 544046 399554 544102
rect 399622 544046 399678 544102
rect 399250 543922 399306 543978
rect 399374 543922 399430 543978
rect 399498 543922 399554 543978
rect 399622 543922 399678 543978
rect 399250 526294 399306 526350
rect 399374 526294 399430 526350
rect 399498 526294 399554 526350
rect 399622 526294 399678 526350
rect 399250 526170 399306 526226
rect 399374 526170 399430 526226
rect 399498 526170 399554 526226
rect 399622 526170 399678 526226
rect 399250 526046 399306 526102
rect 399374 526046 399430 526102
rect 399498 526046 399554 526102
rect 399622 526046 399678 526102
rect 399250 525922 399306 525978
rect 399374 525922 399430 525978
rect 399498 525922 399554 525978
rect 399622 525922 399678 525978
rect 399250 508294 399306 508350
rect 399374 508294 399430 508350
rect 399498 508294 399554 508350
rect 399622 508294 399678 508350
rect 399250 508170 399306 508226
rect 399374 508170 399430 508226
rect 399498 508170 399554 508226
rect 399622 508170 399678 508226
rect 399250 508046 399306 508102
rect 399374 508046 399430 508102
rect 399498 508046 399554 508102
rect 399622 508046 399678 508102
rect 399250 507922 399306 507978
rect 399374 507922 399430 507978
rect 399498 507922 399554 507978
rect 399622 507922 399678 507978
rect 399250 490294 399306 490350
rect 399374 490294 399430 490350
rect 399498 490294 399554 490350
rect 399622 490294 399678 490350
rect 399250 490170 399306 490226
rect 399374 490170 399430 490226
rect 399498 490170 399554 490226
rect 399622 490170 399678 490226
rect 399250 490046 399306 490102
rect 399374 490046 399430 490102
rect 399498 490046 399554 490102
rect 399622 490046 399678 490102
rect 399250 489922 399306 489978
rect 399374 489922 399430 489978
rect 399498 489922 399554 489978
rect 399622 489922 399678 489978
rect 399250 472294 399306 472350
rect 399374 472294 399430 472350
rect 399498 472294 399554 472350
rect 399622 472294 399678 472350
rect 399250 472170 399306 472226
rect 399374 472170 399430 472226
rect 399498 472170 399554 472226
rect 399622 472170 399678 472226
rect 399250 472046 399306 472102
rect 399374 472046 399430 472102
rect 399498 472046 399554 472102
rect 399622 472046 399678 472102
rect 399250 471922 399306 471978
rect 399374 471922 399430 471978
rect 399498 471922 399554 471978
rect 399622 471922 399678 471978
rect 399250 454294 399306 454350
rect 399374 454294 399430 454350
rect 399498 454294 399554 454350
rect 399622 454294 399678 454350
rect 399250 454170 399306 454226
rect 399374 454170 399430 454226
rect 399498 454170 399554 454226
rect 399622 454170 399678 454226
rect 399250 454046 399306 454102
rect 399374 454046 399430 454102
rect 399498 454046 399554 454102
rect 399622 454046 399678 454102
rect 399250 453922 399306 453978
rect 399374 453922 399430 453978
rect 399498 453922 399554 453978
rect 399622 453922 399678 453978
rect 399250 436294 399306 436350
rect 399374 436294 399430 436350
rect 399498 436294 399554 436350
rect 399622 436294 399678 436350
rect 399250 436170 399306 436226
rect 399374 436170 399430 436226
rect 399498 436170 399554 436226
rect 399622 436170 399678 436226
rect 399250 436046 399306 436102
rect 399374 436046 399430 436102
rect 399498 436046 399554 436102
rect 399622 436046 399678 436102
rect 399250 435922 399306 435978
rect 399374 435922 399430 435978
rect 399498 435922 399554 435978
rect 399622 435922 399678 435978
rect 399250 418294 399306 418350
rect 399374 418294 399430 418350
rect 399498 418294 399554 418350
rect 399622 418294 399678 418350
rect 399250 418170 399306 418226
rect 399374 418170 399430 418226
rect 399498 418170 399554 418226
rect 399622 418170 399678 418226
rect 399250 418046 399306 418102
rect 399374 418046 399430 418102
rect 399498 418046 399554 418102
rect 399622 418046 399678 418102
rect 399250 417922 399306 417978
rect 399374 417922 399430 417978
rect 399498 417922 399554 417978
rect 399622 417922 399678 417978
rect 399250 400294 399306 400350
rect 399374 400294 399430 400350
rect 399498 400294 399554 400350
rect 399622 400294 399678 400350
rect 399250 400170 399306 400226
rect 399374 400170 399430 400226
rect 399498 400170 399554 400226
rect 399622 400170 399678 400226
rect 399250 400046 399306 400102
rect 399374 400046 399430 400102
rect 399498 400046 399554 400102
rect 399622 400046 399678 400102
rect 399250 399922 399306 399978
rect 399374 399922 399430 399978
rect 399498 399922 399554 399978
rect 399622 399922 399678 399978
rect 399250 382294 399306 382350
rect 399374 382294 399430 382350
rect 399498 382294 399554 382350
rect 399622 382294 399678 382350
rect 399250 382170 399306 382226
rect 399374 382170 399430 382226
rect 399498 382170 399554 382226
rect 399622 382170 399678 382226
rect 399250 382046 399306 382102
rect 399374 382046 399430 382102
rect 399498 382046 399554 382102
rect 399622 382046 399678 382102
rect 399250 381922 399306 381978
rect 399374 381922 399430 381978
rect 399498 381922 399554 381978
rect 399622 381922 399678 381978
rect 399250 364294 399306 364350
rect 399374 364294 399430 364350
rect 399498 364294 399554 364350
rect 399622 364294 399678 364350
rect 399250 364170 399306 364226
rect 399374 364170 399430 364226
rect 399498 364170 399554 364226
rect 399622 364170 399678 364226
rect 399250 364046 399306 364102
rect 399374 364046 399430 364102
rect 399498 364046 399554 364102
rect 399622 364046 399678 364102
rect 399250 363922 399306 363978
rect 399374 363922 399430 363978
rect 399498 363922 399554 363978
rect 399622 363922 399678 363978
rect 399250 346294 399306 346350
rect 399374 346294 399430 346350
rect 399498 346294 399554 346350
rect 399622 346294 399678 346350
rect 399250 346170 399306 346226
rect 399374 346170 399430 346226
rect 399498 346170 399554 346226
rect 399622 346170 399678 346226
rect 399250 346046 399306 346102
rect 399374 346046 399430 346102
rect 399498 346046 399554 346102
rect 399622 346046 399678 346102
rect 399250 345922 399306 345978
rect 399374 345922 399430 345978
rect 399498 345922 399554 345978
rect 399622 345922 399678 345978
rect 399250 328294 399306 328350
rect 399374 328294 399430 328350
rect 399498 328294 399554 328350
rect 399622 328294 399678 328350
rect 399250 328170 399306 328226
rect 399374 328170 399430 328226
rect 399498 328170 399554 328226
rect 399622 328170 399678 328226
rect 399250 328046 399306 328102
rect 399374 328046 399430 328102
rect 399498 328046 399554 328102
rect 399622 328046 399678 328102
rect 399250 327922 399306 327978
rect 399374 327922 399430 327978
rect 399498 327922 399554 327978
rect 399622 327922 399678 327978
rect 399250 310294 399306 310350
rect 399374 310294 399430 310350
rect 399498 310294 399554 310350
rect 399622 310294 399678 310350
rect 399250 310170 399306 310226
rect 399374 310170 399430 310226
rect 399498 310170 399554 310226
rect 399622 310170 399678 310226
rect 399250 310046 399306 310102
rect 399374 310046 399430 310102
rect 399498 310046 399554 310102
rect 399622 310046 399678 310102
rect 399250 309922 399306 309978
rect 399374 309922 399430 309978
rect 399498 309922 399554 309978
rect 399622 309922 399678 309978
rect 399250 292294 399306 292350
rect 399374 292294 399430 292350
rect 399498 292294 399554 292350
rect 399622 292294 399678 292350
rect 399250 292170 399306 292226
rect 399374 292170 399430 292226
rect 399498 292170 399554 292226
rect 399622 292170 399678 292226
rect 399250 292046 399306 292102
rect 399374 292046 399430 292102
rect 399498 292046 399554 292102
rect 399622 292046 399678 292102
rect 399250 291922 399306 291978
rect 399374 291922 399430 291978
rect 399498 291922 399554 291978
rect 399622 291922 399678 291978
rect 399250 274294 399306 274350
rect 399374 274294 399430 274350
rect 399498 274294 399554 274350
rect 399622 274294 399678 274350
rect 399250 274170 399306 274226
rect 399374 274170 399430 274226
rect 399498 274170 399554 274226
rect 399622 274170 399678 274226
rect 399250 274046 399306 274102
rect 399374 274046 399430 274102
rect 399498 274046 399554 274102
rect 399622 274046 399678 274102
rect 399250 273922 399306 273978
rect 399374 273922 399430 273978
rect 399498 273922 399554 273978
rect 399622 273922 399678 273978
rect 399250 256294 399306 256350
rect 399374 256294 399430 256350
rect 399498 256294 399554 256350
rect 399622 256294 399678 256350
rect 399250 256170 399306 256226
rect 399374 256170 399430 256226
rect 399498 256170 399554 256226
rect 399622 256170 399678 256226
rect 399250 256046 399306 256102
rect 399374 256046 399430 256102
rect 399498 256046 399554 256102
rect 399622 256046 399678 256102
rect 399250 255922 399306 255978
rect 399374 255922 399430 255978
rect 399498 255922 399554 255978
rect 399622 255922 399678 255978
rect 399250 238294 399306 238350
rect 399374 238294 399430 238350
rect 399498 238294 399554 238350
rect 399622 238294 399678 238350
rect 399250 238170 399306 238226
rect 399374 238170 399430 238226
rect 399498 238170 399554 238226
rect 399622 238170 399678 238226
rect 399250 238046 399306 238102
rect 399374 238046 399430 238102
rect 399498 238046 399554 238102
rect 399622 238046 399678 238102
rect 399250 237922 399306 237978
rect 399374 237922 399430 237978
rect 399498 237922 399554 237978
rect 399622 237922 399678 237978
rect 399250 220294 399306 220350
rect 399374 220294 399430 220350
rect 399498 220294 399554 220350
rect 399622 220294 399678 220350
rect 399250 220170 399306 220226
rect 399374 220170 399430 220226
rect 399498 220170 399554 220226
rect 399622 220170 399678 220226
rect 399250 220046 399306 220102
rect 399374 220046 399430 220102
rect 399498 220046 399554 220102
rect 399622 220046 399678 220102
rect 399250 219922 399306 219978
rect 399374 219922 399430 219978
rect 399498 219922 399554 219978
rect 399622 219922 399678 219978
rect 402970 598116 403026 598172
rect 403094 598116 403150 598172
rect 403218 598116 403274 598172
rect 403342 598116 403398 598172
rect 402970 597992 403026 598048
rect 403094 597992 403150 598048
rect 403218 597992 403274 598048
rect 403342 597992 403398 598048
rect 402970 597868 403026 597924
rect 403094 597868 403150 597924
rect 403218 597868 403274 597924
rect 403342 597868 403398 597924
rect 402970 597744 403026 597800
rect 403094 597744 403150 597800
rect 403218 597744 403274 597800
rect 403342 597744 403398 597800
rect 417250 597156 417306 597212
rect 417374 597156 417430 597212
rect 417498 597156 417554 597212
rect 417622 597156 417678 597212
rect 417250 597032 417306 597088
rect 417374 597032 417430 597088
rect 417498 597032 417554 597088
rect 417622 597032 417678 597088
rect 417250 596908 417306 596964
rect 417374 596908 417430 596964
rect 417498 596908 417554 596964
rect 417622 596908 417678 596964
rect 417250 596784 417306 596840
rect 417374 596784 417430 596840
rect 417498 596784 417554 596840
rect 417622 596784 417678 596840
rect 402970 586294 403026 586350
rect 403094 586294 403150 586350
rect 403218 586294 403274 586350
rect 403342 586294 403398 586350
rect 402970 586170 403026 586226
rect 403094 586170 403150 586226
rect 403218 586170 403274 586226
rect 403342 586170 403398 586226
rect 402970 586046 403026 586102
rect 403094 586046 403150 586102
rect 403218 586046 403274 586102
rect 403342 586046 403398 586102
rect 402970 585922 403026 585978
rect 403094 585922 403150 585978
rect 403218 585922 403274 585978
rect 403342 585922 403398 585978
rect 402970 568294 403026 568350
rect 403094 568294 403150 568350
rect 403218 568294 403274 568350
rect 403342 568294 403398 568350
rect 402970 568170 403026 568226
rect 403094 568170 403150 568226
rect 403218 568170 403274 568226
rect 403342 568170 403398 568226
rect 402970 568046 403026 568102
rect 403094 568046 403150 568102
rect 403218 568046 403274 568102
rect 403342 568046 403398 568102
rect 402970 567922 403026 567978
rect 403094 567922 403150 567978
rect 403218 567922 403274 567978
rect 403342 567922 403398 567978
rect 402970 550294 403026 550350
rect 403094 550294 403150 550350
rect 403218 550294 403274 550350
rect 403342 550294 403398 550350
rect 402970 550170 403026 550226
rect 403094 550170 403150 550226
rect 403218 550170 403274 550226
rect 403342 550170 403398 550226
rect 402970 550046 403026 550102
rect 403094 550046 403150 550102
rect 403218 550046 403274 550102
rect 403342 550046 403398 550102
rect 402970 549922 403026 549978
rect 403094 549922 403150 549978
rect 403218 549922 403274 549978
rect 403342 549922 403398 549978
rect 402970 532294 403026 532350
rect 403094 532294 403150 532350
rect 403218 532294 403274 532350
rect 403342 532294 403398 532350
rect 402970 532170 403026 532226
rect 403094 532170 403150 532226
rect 403218 532170 403274 532226
rect 403342 532170 403398 532226
rect 402970 532046 403026 532102
rect 403094 532046 403150 532102
rect 403218 532046 403274 532102
rect 403342 532046 403398 532102
rect 402970 531922 403026 531978
rect 403094 531922 403150 531978
rect 403218 531922 403274 531978
rect 403342 531922 403398 531978
rect 402970 514294 403026 514350
rect 403094 514294 403150 514350
rect 403218 514294 403274 514350
rect 403342 514294 403398 514350
rect 402970 514170 403026 514226
rect 403094 514170 403150 514226
rect 403218 514170 403274 514226
rect 403342 514170 403398 514226
rect 402970 514046 403026 514102
rect 403094 514046 403150 514102
rect 403218 514046 403274 514102
rect 403342 514046 403398 514102
rect 402970 513922 403026 513978
rect 403094 513922 403150 513978
rect 403218 513922 403274 513978
rect 403342 513922 403398 513978
rect 402970 496294 403026 496350
rect 403094 496294 403150 496350
rect 403218 496294 403274 496350
rect 403342 496294 403398 496350
rect 402970 496170 403026 496226
rect 403094 496170 403150 496226
rect 403218 496170 403274 496226
rect 403342 496170 403398 496226
rect 402970 496046 403026 496102
rect 403094 496046 403150 496102
rect 403218 496046 403274 496102
rect 403342 496046 403398 496102
rect 402970 495922 403026 495978
rect 403094 495922 403150 495978
rect 403218 495922 403274 495978
rect 403342 495922 403398 495978
rect 402970 478294 403026 478350
rect 403094 478294 403150 478350
rect 403218 478294 403274 478350
rect 403342 478294 403398 478350
rect 402970 478170 403026 478226
rect 403094 478170 403150 478226
rect 403218 478170 403274 478226
rect 403342 478170 403398 478226
rect 402970 478046 403026 478102
rect 403094 478046 403150 478102
rect 403218 478046 403274 478102
rect 403342 478046 403398 478102
rect 402970 477922 403026 477978
rect 403094 477922 403150 477978
rect 403218 477922 403274 477978
rect 403342 477922 403398 477978
rect 402970 460294 403026 460350
rect 403094 460294 403150 460350
rect 403218 460294 403274 460350
rect 403342 460294 403398 460350
rect 402970 460170 403026 460226
rect 403094 460170 403150 460226
rect 403218 460170 403274 460226
rect 403342 460170 403398 460226
rect 402970 460046 403026 460102
rect 403094 460046 403150 460102
rect 403218 460046 403274 460102
rect 403342 460046 403398 460102
rect 402970 459922 403026 459978
rect 403094 459922 403150 459978
rect 403218 459922 403274 459978
rect 403342 459922 403398 459978
rect 402970 442294 403026 442350
rect 403094 442294 403150 442350
rect 403218 442294 403274 442350
rect 403342 442294 403398 442350
rect 402970 442170 403026 442226
rect 403094 442170 403150 442226
rect 403218 442170 403274 442226
rect 403342 442170 403398 442226
rect 402970 442046 403026 442102
rect 403094 442046 403150 442102
rect 403218 442046 403274 442102
rect 403342 442046 403398 442102
rect 402970 441922 403026 441978
rect 403094 441922 403150 441978
rect 403218 441922 403274 441978
rect 403342 441922 403398 441978
rect 402970 424294 403026 424350
rect 403094 424294 403150 424350
rect 403218 424294 403274 424350
rect 403342 424294 403398 424350
rect 402970 424170 403026 424226
rect 403094 424170 403150 424226
rect 403218 424170 403274 424226
rect 403342 424170 403398 424226
rect 402970 424046 403026 424102
rect 403094 424046 403150 424102
rect 403218 424046 403274 424102
rect 403342 424046 403398 424102
rect 402970 423922 403026 423978
rect 403094 423922 403150 423978
rect 403218 423922 403274 423978
rect 403342 423922 403398 423978
rect 402970 406294 403026 406350
rect 403094 406294 403150 406350
rect 403218 406294 403274 406350
rect 403342 406294 403398 406350
rect 402970 406170 403026 406226
rect 403094 406170 403150 406226
rect 403218 406170 403274 406226
rect 403342 406170 403398 406226
rect 402970 406046 403026 406102
rect 403094 406046 403150 406102
rect 403218 406046 403274 406102
rect 403342 406046 403398 406102
rect 402970 405922 403026 405978
rect 403094 405922 403150 405978
rect 403218 405922 403274 405978
rect 403342 405922 403398 405978
rect 402970 388294 403026 388350
rect 403094 388294 403150 388350
rect 403218 388294 403274 388350
rect 403342 388294 403398 388350
rect 402970 388170 403026 388226
rect 403094 388170 403150 388226
rect 403218 388170 403274 388226
rect 403342 388170 403398 388226
rect 402970 388046 403026 388102
rect 403094 388046 403150 388102
rect 403218 388046 403274 388102
rect 403342 388046 403398 388102
rect 402970 387922 403026 387978
rect 403094 387922 403150 387978
rect 403218 387922 403274 387978
rect 403342 387922 403398 387978
rect 402970 370294 403026 370350
rect 403094 370294 403150 370350
rect 403218 370294 403274 370350
rect 403342 370294 403398 370350
rect 402970 370170 403026 370226
rect 403094 370170 403150 370226
rect 403218 370170 403274 370226
rect 403342 370170 403398 370226
rect 402970 370046 403026 370102
rect 403094 370046 403150 370102
rect 403218 370046 403274 370102
rect 403342 370046 403398 370102
rect 402970 369922 403026 369978
rect 403094 369922 403150 369978
rect 403218 369922 403274 369978
rect 403342 369922 403398 369978
rect 402970 352294 403026 352350
rect 403094 352294 403150 352350
rect 403218 352294 403274 352350
rect 403342 352294 403398 352350
rect 402970 352170 403026 352226
rect 403094 352170 403150 352226
rect 403218 352170 403274 352226
rect 403342 352170 403398 352226
rect 402970 352046 403026 352102
rect 403094 352046 403150 352102
rect 403218 352046 403274 352102
rect 403342 352046 403398 352102
rect 402970 351922 403026 351978
rect 403094 351922 403150 351978
rect 403218 351922 403274 351978
rect 403342 351922 403398 351978
rect 402970 334294 403026 334350
rect 403094 334294 403150 334350
rect 403218 334294 403274 334350
rect 403342 334294 403398 334350
rect 402970 334170 403026 334226
rect 403094 334170 403150 334226
rect 403218 334170 403274 334226
rect 403342 334170 403398 334226
rect 402970 334046 403026 334102
rect 403094 334046 403150 334102
rect 403218 334046 403274 334102
rect 403342 334046 403398 334102
rect 402970 333922 403026 333978
rect 403094 333922 403150 333978
rect 403218 333922 403274 333978
rect 403342 333922 403398 333978
rect 402970 316294 403026 316350
rect 403094 316294 403150 316350
rect 403218 316294 403274 316350
rect 403342 316294 403398 316350
rect 402970 316170 403026 316226
rect 403094 316170 403150 316226
rect 403218 316170 403274 316226
rect 403342 316170 403398 316226
rect 402970 316046 403026 316102
rect 403094 316046 403150 316102
rect 403218 316046 403274 316102
rect 403342 316046 403398 316102
rect 402970 315922 403026 315978
rect 403094 315922 403150 315978
rect 403218 315922 403274 315978
rect 403342 315922 403398 315978
rect 402970 298294 403026 298350
rect 403094 298294 403150 298350
rect 403218 298294 403274 298350
rect 403342 298294 403398 298350
rect 402970 298170 403026 298226
rect 403094 298170 403150 298226
rect 403218 298170 403274 298226
rect 403342 298170 403398 298226
rect 402970 298046 403026 298102
rect 403094 298046 403150 298102
rect 403218 298046 403274 298102
rect 403342 298046 403398 298102
rect 402970 297922 403026 297978
rect 403094 297922 403150 297978
rect 403218 297922 403274 297978
rect 403342 297922 403398 297978
rect 402970 280294 403026 280350
rect 403094 280294 403150 280350
rect 403218 280294 403274 280350
rect 403342 280294 403398 280350
rect 402970 280170 403026 280226
rect 403094 280170 403150 280226
rect 403218 280170 403274 280226
rect 403342 280170 403398 280226
rect 402970 280046 403026 280102
rect 403094 280046 403150 280102
rect 403218 280046 403274 280102
rect 403342 280046 403398 280102
rect 402970 279922 403026 279978
rect 403094 279922 403150 279978
rect 403218 279922 403274 279978
rect 403342 279922 403398 279978
rect 402970 262294 403026 262350
rect 403094 262294 403150 262350
rect 403218 262294 403274 262350
rect 403342 262294 403398 262350
rect 402970 262170 403026 262226
rect 403094 262170 403150 262226
rect 403218 262170 403274 262226
rect 403342 262170 403398 262226
rect 402970 262046 403026 262102
rect 403094 262046 403150 262102
rect 403218 262046 403274 262102
rect 403342 262046 403398 262102
rect 402970 261922 403026 261978
rect 403094 261922 403150 261978
rect 403218 261922 403274 261978
rect 403342 261922 403398 261978
rect 402970 244294 403026 244350
rect 403094 244294 403150 244350
rect 403218 244294 403274 244350
rect 403342 244294 403398 244350
rect 402970 244170 403026 244226
rect 403094 244170 403150 244226
rect 403218 244170 403274 244226
rect 403342 244170 403398 244226
rect 402970 244046 403026 244102
rect 403094 244046 403150 244102
rect 403218 244046 403274 244102
rect 403342 244046 403398 244102
rect 402970 243922 403026 243978
rect 403094 243922 403150 243978
rect 403218 243922 403274 243978
rect 403342 243922 403398 243978
rect 402970 226294 403026 226350
rect 403094 226294 403150 226350
rect 403218 226294 403274 226350
rect 403342 226294 403398 226350
rect 402970 226170 403026 226226
rect 403094 226170 403150 226226
rect 403218 226170 403274 226226
rect 403342 226170 403398 226226
rect 402970 226046 403026 226102
rect 403094 226046 403150 226102
rect 403218 226046 403274 226102
rect 403342 226046 403398 226102
rect 402970 225922 403026 225978
rect 403094 225922 403150 225978
rect 403218 225922 403274 225978
rect 403342 225922 403398 225978
rect 417250 580294 417306 580350
rect 417374 580294 417430 580350
rect 417498 580294 417554 580350
rect 417622 580294 417678 580350
rect 417250 580170 417306 580226
rect 417374 580170 417430 580226
rect 417498 580170 417554 580226
rect 417622 580170 417678 580226
rect 417250 580046 417306 580102
rect 417374 580046 417430 580102
rect 417498 580046 417554 580102
rect 417622 580046 417678 580102
rect 417250 579922 417306 579978
rect 417374 579922 417430 579978
rect 417498 579922 417554 579978
rect 417622 579922 417678 579978
rect 417250 562294 417306 562350
rect 417374 562294 417430 562350
rect 417498 562294 417554 562350
rect 417622 562294 417678 562350
rect 417250 562170 417306 562226
rect 417374 562170 417430 562226
rect 417498 562170 417554 562226
rect 417622 562170 417678 562226
rect 417250 562046 417306 562102
rect 417374 562046 417430 562102
rect 417498 562046 417554 562102
rect 417622 562046 417678 562102
rect 417250 561922 417306 561978
rect 417374 561922 417430 561978
rect 417498 561922 417554 561978
rect 417622 561922 417678 561978
rect 417250 544294 417306 544350
rect 417374 544294 417430 544350
rect 417498 544294 417554 544350
rect 417622 544294 417678 544350
rect 417250 544170 417306 544226
rect 417374 544170 417430 544226
rect 417498 544170 417554 544226
rect 417622 544170 417678 544226
rect 417250 544046 417306 544102
rect 417374 544046 417430 544102
rect 417498 544046 417554 544102
rect 417622 544046 417678 544102
rect 417250 543922 417306 543978
rect 417374 543922 417430 543978
rect 417498 543922 417554 543978
rect 417622 543922 417678 543978
rect 417250 526294 417306 526350
rect 417374 526294 417430 526350
rect 417498 526294 417554 526350
rect 417622 526294 417678 526350
rect 417250 526170 417306 526226
rect 417374 526170 417430 526226
rect 417498 526170 417554 526226
rect 417622 526170 417678 526226
rect 417250 526046 417306 526102
rect 417374 526046 417430 526102
rect 417498 526046 417554 526102
rect 417622 526046 417678 526102
rect 417250 525922 417306 525978
rect 417374 525922 417430 525978
rect 417498 525922 417554 525978
rect 417622 525922 417678 525978
rect 417250 508294 417306 508350
rect 417374 508294 417430 508350
rect 417498 508294 417554 508350
rect 417622 508294 417678 508350
rect 417250 508170 417306 508226
rect 417374 508170 417430 508226
rect 417498 508170 417554 508226
rect 417622 508170 417678 508226
rect 417250 508046 417306 508102
rect 417374 508046 417430 508102
rect 417498 508046 417554 508102
rect 417622 508046 417678 508102
rect 417250 507922 417306 507978
rect 417374 507922 417430 507978
rect 417498 507922 417554 507978
rect 417622 507922 417678 507978
rect 417250 490294 417306 490350
rect 417374 490294 417430 490350
rect 417498 490294 417554 490350
rect 417622 490294 417678 490350
rect 417250 490170 417306 490226
rect 417374 490170 417430 490226
rect 417498 490170 417554 490226
rect 417622 490170 417678 490226
rect 417250 490046 417306 490102
rect 417374 490046 417430 490102
rect 417498 490046 417554 490102
rect 417622 490046 417678 490102
rect 417250 489922 417306 489978
rect 417374 489922 417430 489978
rect 417498 489922 417554 489978
rect 417622 489922 417678 489978
rect 417250 472294 417306 472350
rect 417374 472294 417430 472350
rect 417498 472294 417554 472350
rect 417622 472294 417678 472350
rect 417250 472170 417306 472226
rect 417374 472170 417430 472226
rect 417498 472170 417554 472226
rect 417622 472170 417678 472226
rect 417250 472046 417306 472102
rect 417374 472046 417430 472102
rect 417498 472046 417554 472102
rect 417622 472046 417678 472102
rect 417250 471922 417306 471978
rect 417374 471922 417430 471978
rect 417498 471922 417554 471978
rect 417622 471922 417678 471978
rect 417250 454294 417306 454350
rect 417374 454294 417430 454350
rect 417498 454294 417554 454350
rect 417622 454294 417678 454350
rect 417250 454170 417306 454226
rect 417374 454170 417430 454226
rect 417498 454170 417554 454226
rect 417622 454170 417678 454226
rect 417250 454046 417306 454102
rect 417374 454046 417430 454102
rect 417498 454046 417554 454102
rect 417622 454046 417678 454102
rect 417250 453922 417306 453978
rect 417374 453922 417430 453978
rect 417498 453922 417554 453978
rect 417622 453922 417678 453978
rect 417250 436294 417306 436350
rect 417374 436294 417430 436350
rect 417498 436294 417554 436350
rect 417622 436294 417678 436350
rect 417250 436170 417306 436226
rect 417374 436170 417430 436226
rect 417498 436170 417554 436226
rect 417622 436170 417678 436226
rect 417250 436046 417306 436102
rect 417374 436046 417430 436102
rect 417498 436046 417554 436102
rect 417622 436046 417678 436102
rect 417250 435922 417306 435978
rect 417374 435922 417430 435978
rect 417498 435922 417554 435978
rect 417622 435922 417678 435978
rect 417250 418294 417306 418350
rect 417374 418294 417430 418350
rect 417498 418294 417554 418350
rect 417622 418294 417678 418350
rect 417250 418170 417306 418226
rect 417374 418170 417430 418226
rect 417498 418170 417554 418226
rect 417622 418170 417678 418226
rect 417250 418046 417306 418102
rect 417374 418046 417430 418102
rect 417498 418046 417554 418102
rect 417622 418046 417678 418102
rect 417250 417922 417306 417978
rect 417374 417922 417430 417978
rect 417498 417922 417554 417978
rect 417622 417922 417678 417978
rect 417250 400294 417306 400350
rect 417374 400294 417430 400350
rect 417498 400294 417554 400350
rect 417622 400294 417678 400350
rect 417250 400170 417306 400226
rect 417374 400170 417430 400226
rect 417498 400170 417554 400226
rect 417622 400170 417678 400226
rect 417250 400046 417306 400102
rect 417374 400046 417430 400102
rect 417498 400046 417554 400102
rect 417622 400046 417678 400102
rect 417250 399922 417306 399978
rect 417374 399922 417430 399978
rect 417498 399922 417554 399978
rect 417622 399922 417678 399978
rect 417250 382294 417306 382350
rect 417374 382294 417430 382350
rect 417498 382294 417554 382350
rect 417622 382294 417678 382350
rect 417250 382170 417306 382226
rect 417374 382170 417430 382226
rect 417498 382170 417554 382226
rect 417622 382170 417678 382226
rect 417250 382046 417306 382102
rect 417374 382046 417430 382102
rect 417498 382046 417554 382102
rect 417622 382046 417678 382102
rect 417250 381922 417306 381978
rect 417374 381922 417430 381978
rect 417498 381922 417554 381978
rect 417622 381922 417678 381978
rect 417250 364294 417306 364350
rect 417374 364294 417430 364350
rect 417498 364294 417554 364350
rect 417622 364294 417678 364350
rect 417250 364170 417306 364226
rect 417374 364170 417430 364226
rect 417498 364170 417554 364226
rect 417622 364170 417678 364226
rect 417250 364046 417306 364102
rect 417374 364046 417430 364102
rect 417498 364046 417554 364102
rect 417622 364046 417678 364102
rect 417250 363922 417306 363978
rect 417374 363922 417430 363978
rect 417498 363922 417554 363978
rect 417622 363922 417678 363978
rect 417250 346294 417306 346350
rect 417374 346294 417430 346350
rect 417498 346294 417554 346350
rect 417622 346294 417678 346350
rect 417250 346170 417306 346226
rect 417374 346170 417430 346226
rect 417498 346170 417554 346226
rect 417622 346170 417678 346226
rect 417250 346046 417306 346102
rect 417374 346046 417430 346102
rect 417498 346046 417554 346102
rect 417622 346046 417678 346102
rect 417250 345922 417306 345978
rect 417374 345922 417430 345978
rect 417498 345922 417554 345978
rect 417622 345922 417678 345978
rect 417250 328294 417306 328350
rect 417374 328294 417430 328350
rect 417498 328294 417554 328350
rect 417622 328294 417678 328350
rect 417250 328170 417306 328226
rect 417374 328170 417430 328226
rect 417498 328170 417554 328226
rect 417622 328170 417678 328226
rect 417250 328046 417306 328102
rect 417374 328046 417430 328102
rect 417498 328046 417554 328102
rect 417622 328046 417678 328102
rect 417250 327922 417306 327978
rect 417374 327922 417430 327978
rect 417498 327922 417554 327978
rect 417622 327922 417678 327978
rect 417250 310294 417306 310350
rect 417374 310294 417430 310350
rect 417498 310294 417554 310350
rect 417622 310294 417678 310350
rect 417250 310170 417306 310226
rect 417374 310170 417430 310226
rect 417498 310170 417554 310226
rect 417622 310170 417678 310226
rect 417250 310046 417306 310102
rect 417374 310046 417430 310102
rect 417498 310046 417554 310102
rect 417622 310046 417678 310102
rect 417250 309922 417306 309978
rect 417374 309922 417430 309978
rect 417498 309922 417554 309978
rect 417622 309922 417678 309978
rect 417250 292294 417306 292350
rect 417374 292294 417430 292350
rect 417498 292294 417554 292350
rect 417622 292294 417678 292350
rect 417250 292170 417306 292226
rect 417374 292170 417430 292226
rect 417498 292170 417554 292226
rect 417622 292170 417678 292226
rect 417250 292046 417306 292102
rect 417374 292046 417430 292102
rect 417498 292046 417554 292102
rect 417622 292046 417678 292102
rect 417250 291922 417306 291978
rect 417374 291922 417430 291978
rect 417498 291922 417554 291978
rect 417622 291922 417678 291978
rect 417250 274294 417306 274350
rect 417374 274294 417430 274350
rect 417498 274294 417554 274350
rect 417622 274294 417678 274350
rect 417250 274170 417306 274226
rect 417374 274170 417430 274226
rect 417498 274170 417554 274226
rect 417622 274170 417678 274226
rect 417250 274046 417306 274102
rect 417374 274046 417430 274102
rect 417498 274046 417554 274102
rect 417622 274046 417678 274102
rect 417250 273922 417306 273978
rect 417374 273922 417430 273978
rect 417498 273922 417554 273978
rect 417622 273922 417678 273978
rect 417250 256294 417306 256350
rect 417374 256294 417430 256350
rect 417498 256294 417554 256350
rect 417622 256294 417678 256350
rect 417250 256170 417306 256226
rect 417374 256170 417430 256226
rect 417498 256170 417554 256226
rect 417622 256170 417678 256226
rect 417250 256046 417306 256102
rect 417374 256046 417430 256102
rect 417498 256046 417554 256102
rect 417622 256046 417678 256102
rect 417250 255922 417306 255978
rect 417374 255922 417430 255978
rect 417498 255922 417554 255978
rect 417622 255922 417678 255978
rect 417250 238294 417306 238350
rect 417374 238294 417430 238350
rect 417498 238294 417554 238350
rect 417622 238294 417678 238350
rect 417250 238170 417306 238226
rect 417374 238170 417430 238226
rect 417498 238170 417554 238226
rect 417622 238170 417678 238226
rect 417250 238046 417306 238102
rect 417374 238046 417430 238102
rect 417498 238046 417554 238102
rect 417622 238046 417678 238102
rect 417250 237922 417306 237978
rect 417374 237922 417430 237978
rect 417498 237922 417554 237978
rect 417622 237922 417678 237978
rect 417250 220294 417306 220350
rect 417374 220294 417430 220350
rect 417498 220294 417554 220350
rect 417622 220294 417678 220350
rect 417250 220170 417306 220226
rect 417374 220170 417430 220226
rect 417498 220170 417554 220226
rect 417622 220170 417678 220226
rect 417250 220046 417306 220102
rect 417374 220046 417430 220102
rect 417498 220046 417554 220102
rect 417622 220046 417678 220102
rect 417250 219922 417306 219978
rect 417374 219922 417430 219978
rect 417498 219922 417554 219978
rect 417622 219922 417678 219978
rect 420970 598116 421026 598172
rect 421094 598116 421150 598172
rect 421218 598116 421274 598172
rect 421342 598116 421398 598172
rect 420970 597992 421026 598048
rect 421094 597992 421150 598048
rect 421218 597992 421274 598048
rect 421342 597992 421398 598048
rect 420970 597868 421026 597924
rect 421094 597868 421150 597924
rect 421218 597868 421274 597924
rect 421342 597868 421398 597924
rect 420970 597744 421026 597800
rect 421094 597744 421150 597800
rect 421218 597744 421274 597800
rect 421342 597744 421398 597800
rect 420970 586294 421026 586350
rect 421094 586294 421150 586350
rect 421218 586294 421274 586350
rect 421342 586294 421398 586350
rect 420970 586170 421026 586226
rect 421094 586170 421150 586226
rect 421218 586170 421274 586226
rect 421342 586170 421398 586226
rect 420970 586046 421026 586102
rect 421094 586046 421150 586102
rect 421218 586046 421274 586102
rect 421342 586046 421398 586102
rect 420970 585922 421026 585978
rect 421094 585922 421150 585978
rect 421218 585922 421274 585978
rect 421342 585922 421398 585978
rect 420970 568294 421026 568350
rect 421094 568294 421150 568350
rect 421218 568294 421274 568350
rect 421342 568294 421398 568350
rect 420970 568170 421026 568226
rect 421094 568170 421150 568226
rect 421218 568170 421274 568226
rect 421342 568170 421398 568226
rect 420970 568046 421026 568102
rect 421094 568046 421150 568102
rect 421218 568046 421274 568102
rect 421342 568046 421398 568102
rect 420970 567922 421026 567978
rect 421094 567922 421150 567978
rect 421218 567922 421274 567978
rect 421342 567922 421398 567978
rect 420970 550294 421026 550350
rect 421094 550294 421150 550350
rect 421218 550294 421274 550350
rect 421342 550294 421398 550350
rect 420970 550170 421026 550226
rect 421094 550170 421150 550226
rect 421218 550170 421274 550226
rect 421342 550170 421398 550226
rect 420970 550046 421026 550102
rect 421094 550046 421150 550102
rect 421218 550046 421274 550102
rect 421342 550046 421398 550102
rect 420970 549922 421026 549978
rect 421094 549922 421150 549978
rect 421218 549922 421274 549978
rect 421342 549922 421398 549978
rect 420970 532294 421026 532350
rect 421094 532294 421150 532350
rect 421218 532294 421274 532350
rect 421342 532294 421398 532350
rect 420970 532170 421026 532226
rect 421094 532170 421150 532226
rect 421218 532170 421274 532226
rect 421342 532170 421398 532226
rect 420970 532046 421026 532102
rect 421094 532046 421150 532102
rect 421218 532046 421274 532102
rect 421342 532046 421398 532102
rect 420970 531922 421026 531978
rect 421094 531922 421150 531978
rect 421218 531922 421274 531978
rect 421342 531922 421398 531978
rect 420970 514294 421026 514350
rect 421094 514294 421150 514350
rect 421218 514294 421274 514350
rect 421342 514294 421398 514350
rect 420970 514170 421026 514226
rect 421094 514170 421150 514226
rect 421218 514170 421274 514226
rect 421342 514170 421398 514226
rect 420970 514046 421026 514102
rect 421094 514046 421150 514102
rect 421218 514046 421274 514102
rect 421342 514046 421398 514102
rect 420970 513922 421026 513978
rect 421094 513922 421150 513978
rect 421218 513922 421274 513978
rect 421342 513922 421398 513978
rect 420970 496294 421026 496350
rect 421094 496294 421150 496350
rect 421218 496294 421274 496350
rect 421342 496294 421398 496350
rect 420970 496170 421026 496226
rect 421094 496170 421150 496226
rect 421218 496170 421274 496226
rect 421342 496170 421398 496226
rect 420970 496046 421026 496102
rect 421094 496046 421150 496102
rect 421218 496046 421274 496102
rect 421342 496046 421398 496102
rect 420970 495922 421026 495978
rect 421094 495922 421150 495978
rect 421218 495922 421274 495978
rect 421342 495922 421398 495978
rect 420970 478294 421026 478350
rect 421094 478294 421150 478350
rect 421218 478294 421274 478350
rect 421342 478294 421398 478350
rect 420970 478170 421026 478226
rect 421094 478170 421150 478226
rect 421218 478170 421274 478226
rect 421342 478170 421398 478226
rect 420970 478046 421026 478102
rect 421094 478046 421150 478102
rect 421218 478046 421274 478102
rect 421342 478046 421398 478102
rect 420970 477922 421026 477978
rect 421094 477922 421150 477978
rect 421218 477922 421274 477978
rect 421342 477922 421398 477978
rect 420970 460294 421026 460350
rect 421094 460294 421150 460350
rect 421218 460294 421274 460350
rect 421342 460294 421398 460350
rect 420970 460170 421026 460226
rect 421094 460170 421150 460226
rect 421218 460170 421274 460226
rect 421342 460170 421398 460226
rect 420970 460046 421026 460102
rect 421094 460046 421150 460102
rect 421218 460046 421274 460102
rect 421342 460046 421398 460102
rect 420970 459922 421026 459978
rect 421094 459922 421150 459978
rect 421218 459922 421274 459978
rect 421342 459922 421398 459978
rect 420970 442294 421026 442350
rect 421094 442294 421150 442350
rect 421218 442294 421274 442350
rect 421342 442294 421398 442350
rect 420970 442170 421026 442226
rect 421094 442170 421150 442226
rect 421218 442170 421274 442226
rect 421342 442170 421398 442226
rect 420970 442046 421026 442102
rect 421094 442046 421150 442102
rect 421218 442046 421274 442102
rect 421342 442046 421398 442102
rect 420970 441922 421026 441978
rect 421094 441922 421150 441978
rect 421218 441922 421274 441978
rect 421342 441922 421398 441978
rect 420970 424294 421026 424350
rect 421094 424294 421150 424350
rect 421218 424294 421274 424350
rect 421342 424294 421398 424350
rect 420970 424170 421026 424226
rect 421094 424170 421150 424226
rect 421218 424170 421274 424226
rect 421342 424170 421398 424226
rect 420970 424046 421026 424102
rect 421094 424046 421150 424102
rect 421218 424046 421274 424102
rect 421342 424046 421398 424102
rect 420970 423922 421026 423978
rect 421094 423922 421150 423978
rect 421218 423922 421274 423978
rect 421342 423922 421398 423978
rect 420970 406294 421026 406350
rect 421094 406294 421150 406350
rect 421218 406294 421274 406350
rect 421342 406294 421398 406350
rect 420970 406170 421026 406226
rect 421094 406170 421150 406226
rect 421218 406170 421274 406226
rect 421342 406170 421398 406226
rect 420970 406046 421026 406102
rect 421094 406046 421150 406102
rect 421218 406046 421274 406102
rect 421342 406046 421398 406102
rect 420970 405922 421026 405978
rect 421094 405922 421150 405978
rect 421218 405922 421274 405978
rect 421342 405922 421398 405978
rect 420970 388294 421026 388350
rect 421094 388294 421150 388350
rect 421218 388294 421274 388350
rect 421342 388294 421398 388350
rect 420970 388170 421026 388226
rect 421094 388170 421150 388226
rect 421218 388170 421274 388226
rect 421342 388170 421398 388226
rect 420970 388046 421026 388102
rect 421094 388046 421150 388102
rect 421218 388046 421274 388102
rect 421342 388046 421398 388102
rect 420970 387922 421026 387978
rect 421094 387922 421150 387978
rect 421218 387922 421274 387978
rect 421342 387922 421398 387978
rect 420970 370294 421026 370350
rect 421094 370294 421150 370350
rect 421218 370294 421274 370350
rect 421342 370294 421398 370350
rect 420970 370170 421026 370226
rect 421094 370170 421150 370226
rect 421218 370170 421274 370226
rect 421342 370170 421398 370226
rect 420970 370046 421026 370102
rect 421094 370046 421150 370102
rect 421218 370046 421274 370102
rect 421342 370046 421398 370102
rect 420970 369922 421026 369978
rect 421094 369922 421150 369978
rect 421218 369922 421274 369978
rect 421342 369922 421398 369978
rect 420970 352294 421026 352350
rect 421094 352294 421150 352350
rect 421218 352294 421274 352350
rect 421342 352294 421398 352350
rect 420970 352170 421026 352226
rect 421094 352170 421150 352226
rect 421218 352170 421274 352226
rect 421342 352170 421398 352226
rect 420970 352046 421026 352102
rect 421094 352046 421150 352102
rect 421218 352046 421274 352102
rect 421342 352046 421398 352102
rect 420970 351922 421026 351978
rect 421094 351922 421150 351978
rect 421218 351922 421274 351978
rect 421342 351922 421398 351978
rect 420970 334294 421026 334350
rect 421094 334294 421150 334350
rect 421218 334294 421274 334350
rect 421342 334294 421398 334350
rect 420970 334170 421026 334226
rect 421094 334170 421150 334226
rect 421218 334170 421274 334226
rect 421342 334170 421398 334226
rect 420970 334046 421026 334102
rect 421094 334046 421150 334102
rect 421218 334046 421274 334102
rect 421342 334046 421398 334102
rect 420970 333922 421026 333978
rect 421094 333922 421150 333978
rect 421218 333922 421274 333978
rect 421342 333922 421398 333978
rect 420970 316294 421026 316350
rect 421094 316294 421150 316350
rect 421218 316294 421274 316350
rect 421342 316294 421398 316350
rect 420970 316170 421026 316226
rect 421094 316170 421150 316226
rect 421218 316170 421274 316226
rect 421342 316170 421398 316226
rect 420970 316046 421026 316102
rect 421094 316046 421150 316102
rect 421218 316046 421274 316102
rect 421342 316046 421398 316102
rect 420970 315922 421026 315978
rect 421094 315922 421150 315978
rect 421218 315922 421274 315978
rect 421342 315922 421398 315978
rect 420970 298294 421026 298350
rect 421094 298294 421150 298350
rect 421218 298294 421274 298350
rect 421342 298294 421398 298350
rect 420970 298170 421026 298226
rect 421094 298170 421150 298226
rect 421218 298170 421274 298226
rect 421342 298170 421398 298226
rect 420970 298046 421026 298102
rect 421094 298046 421150 298102
rect 421218 298046 421274 298102
rect 421342 298046 421398 298102
rect 420970 297922 421026 297978
rect 421094 297922 421150 297978
rect 421218 297922 421274 297978
rect 421342 297922 421398 297978
rect 420970 280294 421026 280350
rect 421094 280294 421150 280350
rect 421218 280294 421274 280350
rect 421342 280294 421398 280350
rect 420970 280170 421026 280226
rect 421094 280170 421150 280226
rect 421218 280170 421274 280226
rect 421342 280170 421398 280226
rect 420970 280046 421026 280102
rect 421094 280046 421150 280102
rect 421218 280046 421274 280102
rect 421342 280046 421398 280102
rect 420970 279922 421026 279978
rect 421094 279922 421150 279978
rect 421218 279922 421274 279978
rect 421342 279922 421398 279978
rect 420970 262294 421026 262350
rect 421094 262294 421150 262350
rect 421218 262294 421274 262350
rect 421342 262294 421398 262350
rect 420970 262170 421026 262226
rect 421094 262170 421150 262226
rect 421218 262170 421274 262226
rect 421342 262170 421398 262226
rect 420970 262046 421026 262102
rect 421094 262046 421150 262102
rect 421218 262046 421274 262102
rect 421342 262046 421398 262102
rect 420970 261922 421026 261978
rect 421094 261922 421150 261978
rect 421218 261922 421274 261978
rect 421342 261922 421398 261978
rect 420970 244294 421026 244350
rect 421094 244294 421150 244350
rect 421218 244294 421274 244350
rect 421342 244294 421398 244350
rect 420970 244170 421026 244226
rect 421094 244170 421150 244226
rect 421218 244170 421274 244226
rect 421342 244170 421398 244226
rect 420970 244046 421026 244102
rect 421094 244046 421150 244102
rect 421218 244046 421274 244102
rect 421342 244046 421398 244102
rect 420970 243922 421026 243978
rect 421094 243922 421150 243978
rect 421218 243922 421274 243978
rect 421342 243922 421398 243978
rect 438970 598116 439026 598172
rect 439094 598116 439150 598172
rect 439218 598116 439274 598172
rect 439342 598116 439398 598172
rect 438970 597992 439026 598048
rect 439094 597992 439150 598048
rect 439218 597992 439274 598048
rect 439342 597992 439398 598048
rect 438970 597868 439026 597924
rect 439094 597868 439150 597924
rect 439218 597868 439274 597924
rect 439342 597868 439398 597924
rect 438970 597744 439026 597800
rect 439094 597744 439150 597800
rect 439218 597744 439274 597800
rect 439342 597744 439398 597800
rect 438970 586294 439026 586350
rect 439094 586294 439150 586350
rect 439218 586294 439274 586350
rect 439342 586294 439398 586350
rect 438970 586170 439026 586226
rect 439094 586170 439150 586226
rect 439218 586170 439274 586226
rect 439342 586170 439398 586226
rect 438970 586046 439026 586102
rect 439094 586046 439150 586102
rect 439218 586046 439274 586102
rect 439342 586046 439398 586102
rect 438970 585922 439026 585978
rect 439094 585922 439150 585978
rect 439218 585922 439274 585978
rect 439342 585922 439398 585978
rect 438970 568294 439026 568350
rect 439094 568294 439150 568350
rect 439218 568294 439274 568350
rect 439342 568294 439398 568350
rect 438970 568170 439026 568226
rect 439094 568170 439150 568226
rect 439218 568170 439274 568226
rect 439342 568170 439398 568226
rect 438970 568046 439026 568102
rect 439094 568046 439150 568102
rect 439218 568046 439274 568102
rect 439342 568046 439398 568102
rect 438970 567922 439026 567978
rect 439094 567922 439150 567978
rect 439218 567922 439274 567978
rect 439342 567922 439398 567978
rect 438970 550294 439026 550350
rect 439094 550294 439150 550350
rect 439218 550294 439274 550350
rect 439342 550294 439398 550350
rect 438970 550170 439026 550226
rect 439094 550170 439150 550226
rect 439218 550170 439274 550226
rect 439342 550170 439398 550226
rect 438970 550046 439026 550102
rect 439094 550046 439150 550102
rect 439218 550046 439274 550102
rect 439342 550046 439398 550102
rect 438970 549922 439026 549978
rect 439094 549922 439150 549978
rect 439218 549922 439274 549978
rect 439342 549922 439398 549978
rect 438970 532294 439026 532350
rect 439094 532294 439150 532350
rect 439218 532294 439274 532350
rect 439342 532294 439398 532350
rect 438970 532170 439026 532226
rect 439094 532170 439150 532226
rect 439218 532170 439274 532226
rect 439342 532170 439398 532226
rect 438970 532046 439026 532102
rect 439094 532046 439150 532102
rect 439218 532046 439274 532102
rect 439342 532046 439398 532102
rect 438970 531922 439026 531978
rect 439094 531922 439150 531978
rect 439218 531922 439274 531978
rect 439342 531922 439398 531978
rect 438970 514294 439026 514350
rect 439094 514294 439150 514350
rect 439218 514294 439274 514350
rect 439342 514294 439398 514350
rect 438970 514170 439026 514226
rect 439094 514170 439150 514226
rect 439218 514170 439274 514226
rect 439342 514170 439398 514226
rect 438970 514046 439026 514102
rect 439094 514046 439150 514102
rect 439218 514046 439274 514102
rect 439342 514046 439398 514102
rect 438970 513922 439026 513978
rect 439094 513922 439150 513978
rect 439218 513922 439274 513978
rect 439342 513922 439398 513978
rect 438970 496294 439026 496350
rect 439094 496294 439150 496350
rect 439218 496294 439274 496350
rect 439342 496294 439398 496350
rect 438970 496170 439026 496226
rect 439094 496170 439150 496226
rect 439218 496170 439274 496226
rect 439342 496170 439398 496226
rect 438970 496046 439026 496102
rect 439094 496046 439150 496102
rect 439218 496046 439274 496102
rect 439342 496046 439398 496102
rect 438970 495922 439026 495978
rect 439094 495922 439150 495978
rect 439218 495922 439274 495978
rect 439342 495922 439398 495978
rect 438970 478294 439026 478350
rect 439094 478294 439150 478350
rect 439218 478294 439274 478350
rect 439342 478294 439398 478350
rect 438970 478170 439026 478226
rect 439094 478170 439150 478226
rect 439218 478170 439274 478226
rect 439342 478170 439398 478226
rect 438970 478046 439026 478102
rect 439094 478046 439150 478102
rect 439218 478046 439274 478102
rect 439342 478046 439398 478102
rect 438970 477922 439026 477978
rect 439094 477922 439150 477978
rect 439218 477922 439274 477978
rect 439342 477922 439398 477978
rect 438970 460294 439026 460350
rect 439094 460294 439150 460350
rect 439218 460294 439274 460350
rect 439342 460294 439398 460350
rect 438970 460170 439026 460226
rect 439094 460170 439150 460226
rect 439218 460170 439274 460226
rect 439342 460170 439398 460226
rect 438970 460046 439026 460102
rect 439094 460046 439150 460102
rect 439218 460046 439274 460102
rect 439342 460046 439398 460102
rect 438970 459922 439026 459978
rect 439094 459922 439150 459978
rect 439218 459922 439274 459978
rect 439342 459922 439398 459978
rect 438970 442294 439026 442350
rect 439094 442294 439150 442350
rect 439218 442294 439274 442350
rect 439342 442294 439398 442350
rect 438970 442170 439026 442226
rect 439094 442170 439150 442226
rect 439218 442170 439274 442226
rect 439342 442170 439398 442226
rect 438970 442046 439026 442102
rect 439094 442046 439150 442102
rect 439218 442046 439274 442102
rect 439342 442046 439398 442102
rect 438970 441922 439026 441978
rect 439094 441922 439150 441978
rect 439218 441922 439274 441978
rect 439342 441922 439398 441978
rect 438970 424294 439026 424350
rect 439094 424294 439150 424350
rect 439218 424294 439274 424350
rect 439342 424294 439398 424350
rect 438970 424170 439026 424226
rect 439094 424170 439150 424226
rect 439218 424170 439274 424226
rect 439342 424170 439398 424226
rect 438970 424046 439026 424102
rect 439094 424046 439150 424102
rect 439218 424046 439274 424102
rect 439342 424046 439398 424102
rect 438970 423922 439026 423978
rect 439094 423922 439150 423978
rect 439218 423922 439274 423978
rect 439342 423922 439398 423978
rect 438970 406294 439026 406350
rect 439094 406294 439150 406350
rect 439218 406294 439274 406350
rect 439342 406294 439398 406350
rect 438970 406170 439026 406226
rect 439094 406170 439150 406226
rect 439218 406170 439274 406226
rect 439342 406170 439398 406226
rect 438970 406046 439026 406102
rect 439094 406046 439150 406102
rect 439218 406046 439274 406102
rect 439342 406046 439398 406102
rect 438970 405922 439026 405978
rect 439094 405922 439150 405978
rect 439218 405922 439274 405978
rect 439342 405922 439398 405978
rect 438970 388294 439026 388350
rect 439094 388294 439150 388350
rect 439218 388294 439274 388350
rect 439342 388294 439398 388350
rect 438970 388170 439026 388226
rect 439094 388170 439150 388226
rect 439218 388170 439274 388226
rect 439342 388170 439398 388226
rect 438970 388046 439026 388102
rect 439094 388046 439150 388102
rect 439218 388046 439274 388102
rect 439342 388046 439398 388102
rect 438970 387922 439026 387978
rect 439094 387922 439150 387978
rect 439218 387922 439274 387978
rect 439342 387922 439398 387978
rect 438970 370294 439026 370350
rect 439094 370294 439150 370350
rect 439218 370294 439274 370350
rect 439342 370294 439398 370350
rect 438970 370170 439026 370226
rect 439094 370170 439150 370226
rect 439218 370170 439274 370226
rect 439342 370170 439398 370226
rect 438970 370046 439026 370102
rect 439094 370046 439150 370102
rect 439218 370046 439274 370102
rect 439342 370046 439398 370102
rect 438970 369922 439026 369978
rect 439094 369922 439150 369978
rect 439218 369922 439274 369978
rect 439342 369922 439398 369978
rect 438970 352294 439026 352350
rect 439094 352294 439150 352350
rect 439218 352294 439274 352350
rect 439342 352294 439398 352350
rect 438970 352170 439026 352226
rect 439094 352170 439150 352226
rect 439218 352170 439274 352226
rect 439342 352170 439398 352226
rect 438970 352046 439026 352102
rect 439094 352046 439150 352102
rect 439218 352046 439274 352102
rect 439342 352046 439398 352102
rect 438970 351922 439026 351978
rect 439094 351922 439150 351978
rect 439218 351922 439274 351978
rect 439342 351922 439398 351978
rect 438970 334294 439026 334350
rect 439094 334294 439150 334350
rect 439218 334294 439274 334350
rect 439342 334294 439398 334350
rect 438970 334170 439026 334226
rect 439094 334170 439150 334226
rect 439218 334170 439274 334226
rect 439342 334170 439398 334226
rect 438970 334046 439026 334102
rect 439094 334046 439150 334102
rect 439218 334046 439274 334102
rect 439342 334046 439398 334102
rect 438970 333922 439026 333978
rect 439094 333922 439150 333978
rect 439218 333922 439274 333978
rect 439342 333922 439398 333978
rect 438970 316294 439026 316350
rect 439094 316294 439150 316350
rect 439218 316294 439274 316350
rect 439342 316294 439398 316350
rect 438970 316170 439026 316226
rect 439094 316170 439150 316226
rect 439218 316170 439274 316226
rect 439342 316170 439398 316226
rect 438970 316046 439026 316102
rect 439094 316046 439150 316102
rect 439218 316046 439274 316102
rect 439342 316046 439398 316102
rect 438970 315922 439026 315978
rect 439094 315922 439150 315978
rect 439218 315922 439274 315978
rect 439342 315922 439398 315978
rect 438970 298294 439026 298350
rect 439094 298294 439150 298350
rect 439218 298294 439274 298350
rect 439342 298294 439398 298350
rect 438970 298170 439026 298226
rect 439094 298170 439150 298226
rect 439218 298170 439274 298226
rect 439342 298170 439398 298226
rect 438970 298046 439026 298102
rect 439094 298046 439150 298102
rect 439218 298046 439274 298102
rect 439342 298046 439398 298102
rect 438970 297922 439026 297978
rect 439094 297922 439150 297978
rect 439218 297922 439274 297978
rect 439342 297922 439398 297978
rect 438970 280294 439026 280350
rect 439094 280294 439150 280350
rect 439218 280294 439274 280350
rect 439342 280294 439398 280350
rect 438970 280170 439026 280226
rect 439094 280170 439150 280226
rect 439218 280170 439274 280226
rect 439342 280170 439398 280226
rect 438970 280046 439026 280102
rect 439094 280046 439150 280102
rect 439218 280046 439274 280102
rect 439342 280046 439398 280102
rect 438970 279922 439026 279978
rect 439094 279922 439150 279978
rect 439218 279922 439274 279978
rect 439342 279922 439398 279978
rect 438970 262294 439026 262350
rect 439094 262294 439150 262350
rect 439218 262294 439274 262350
rect 439342 262294 439398 262350
rect 438970 262170 439026 262226
rect 439094 262170 439150 262226
rect 439218 262170 439274 262226
rect 439342 262170 439398 262226
rect 438970 262046 439026 262102
rect 439094 262046 439150 262102
rect 439218 262046 439274 262102
rect 439342 262046 439398 262102
rect 438970 261922 439026 261978
rect 439094 261922 439150 261978
rect 439218 261922 439274 261978
rect 439342 261922 439398 261978
rect 438970 244294 439026 244350
rect 439094 244294 439150 244350
rect 439218 244294 439274 244350
rect 439342 244294 439398 244350
rect 438970 244170 439026 244226
rect 439094 244170 439150 244226
rect 439218 244170 439274 244226
rect 439342 244170 439398 244226
rect 438970 244046 439026 244102
rect 439094 244046 439150 244102
rect 439218 244046 439274 244102
rect 439342 244046 439398 244102
rect 438970 243922 439026 243978
rect 439094 243922 439150 243978
rect 439218 243922 439274 243978
rect 439342 243922 439398 243978
rect 420970 226294 421026 226350
rect 421094 226294 421150 226350
rect 421218 226294 421274 226350
rect 421342 226294 421398 226350
rect 420970 226170 421026 226226
rect 421094 226170 421150 226226
rect 421218 226170 421274 226226
rect 421342 226170 421398 226226
rect 420970 226046 421026 226102
rect 421094 226046 421150 226102
rect 421218 226046 421274 226102
rect 421342 226046 421398 226102
rect 420970 225922 421026 225978
rect 421094 225922 421150 225978
rect 421218 225922 421274 225978
rect 421342 225922 421398 225978
rect 435250 238294 435306 238350
rect 435374 238294 435430 238350
rect 435498 238294 435554 238350
rect 435622 238294 435678 238350
rect 435250 238170 435306 238226
rect 435374 238170 435430 238226
rect 435498 238170 435554 238226
rect 435622 238170 435678 238226
rect 435250 238046 435306 238102
rect 435374 238046 435430 238102
rect 435498 238046 435554 238102
rect 435622 238046 435678 238102
rect 435250 237922 435306 237978
rect 435374 237922 435430 237978
rect 435498 237922 435554 237978
rect 435622 237922 435678 237978
rect 435250 220294 435306 220350
rect 435374 220294 435430 220350
rect 435498 220294 435554 220350
rect 435622 220294 435678 220350
rect 435250 220170 435306 220226
rect 435374 220170 435430 220226
rect 435498 220170 435554 220226
rect 435622 220170 435678 220226
rect 435250 220046 435306 220102
rect 435374 220046 435430 220102
rect 435498 220046 435554 220102
rect 435622 220046 435678 220102
rect 435250 219922 435306 219978
rect 435374 219922 435430 219978
rect 435498 219922 435554 219978
rect 435622 219922 435678 219978
rect 438970 226294 439026 226350
rect 439094 226294 439150 226350
rect 439218 226294 439274 226350
rect 439342 226294 439398 226350
rect 438970 226170 439026 226226
rect 439094 226170 439150 226226
rect 439218 226170 439274 226226
rect 439342 226170 439398 226226
rect 438970 226046 439026 226102
rect 439094 226046 439150 226102
rect 439218 226046 439274 226102
rect 439342 226046 439398 226102
rect 438970 225922 439026 225978
rect 439094 225922 439150 225978
rect 439218 225922 439274 225978
rect 439342 225922 439398 225978
rect 453250 597156 453306 597212
rect 453374 597156 453430 597212
rect 453498 597156 453554 597212
rect 453622 597156 453678 597212
rect 453250 597032 453306 597088
rect 453374 597032 453430 597088
rect 453498 597032 453554 597088
rect 453622 597032 453678 597088
rect 453250 596908 453306 596964
rect 453374 596908 453430 596964
rect 453498 596908 453554 596964
rect 453622 596908 453678 596964
rect 453250 596784 453306 596840
rect 453374 596784 453430 596840
rect 453498 596784 453554 596840
rect 453622 596784 453678 596840
rect 453250 580294 453306 580350
rect 453374 580294 453430 580350
rect 453498 580294 453554 580350
rect 453622 580294 453678 580350
rect 453250 580170 453306 580226
rect 453374 580170 453430 580226
rect 453498 580170 453554 580226
rect 453622 580170 453678 580226
rect 453250 580046 453306 580102
rect 453374 580046 453430 580102
rect 453498 580046 453554 580102
rect 453622 580046 453678 580102
rect 453250 579922 453306 579978
rect 453374 579922 453430 579978
rect 453498 579922 453554 579978
rect 453622 579922 453678 579978
rect 453250 562294 453306 562350
rect 453374 562294 453430 562350
rect 453498 562294 453554 562350
rect 453622 562294 453678 562350
rect 453250 562170 453306 562226
rect 453374 562170 453430 562226
rect 453498 562170 453554 562226
rect 453622 562170 453678 562226
rect 453250 562046 453306 562102
rect 453374 562046 453430 562102
rect 453498 562046 453554 562102
rect 453622 562046 453678 562102
rect 453250 561922 453306 561978
rect 453374 561922 453430 561978
rect 453498 561922 453554 561978
rect 453622 561922 453678 561978
rect 453250 544294 453306 544350
rect 453374 544294 453430 544350
rect 453498 544294 453554 544350
rect 453622 544294 453678 544350
rect 453250 544170 453306 544226
rect 453374 544170 453430 544226
rect 453498 544170 453554 544226
rect 453622 544170 453678 544226
rect 453250 544046 453306 544102
rect 453374 544046 453430 544102
rect 453498 544046 453554 544102
rect 453622 544046 453678 544102
rect 453250 543922 453306 543978
rect 453374 543922 453430 543978
rect 453498 543922 453554 543978
rect 453622 543922 453678 543978
rect 453250 526294 453306 526350
rect 453374 526294 453430 526350
rect 453498 526294 453554 526350
rect 453622 526294 453678 526350
rect 453250 526170 453306 526226
rect 453374 526170 453430 526226
rect 453498 526170 453554 526226
rect 453622 526170 453678 526226
rect 453250 526046 453306 526102
rect 453374 526046 453430 526102
rect 453498 526046 453554 526102
rect 453622 526046 453678 526102
rect 453250 525922 453306 525978
rect 453374 525922 453430 525978
rect 453498 525922 453554 525978
rect 453622 525922 453678 525978
rect 453250 508294 453306 508350
rect 453374 508294 453430 508350
rect 453498 508294 453554 508350
rect 453622 508294 453678 508350
rect 453250 508170 453306 508226
rect 453374 508170 453430 508226
rect 453498 508170 453554 508226
rect 453622 508170 453678 508226
rect 453250 508046 453306 508102
rect 453374 508046 453430 508102
rect 453498 508046 453554 508102
rect 453622 508046 453678 508102
rect 453250 507922 453306 507978
rect 453374 507922 453430 507978
rect 453498 507922 453554 507978
rect 453622 507922 453678 507978
rect 453250 490294 453306 490350
rect 453374 490294 453430 490350
rect 453498 490294 453554 490350
rect 453622 490294 453678 490350
rect 453250 490170 453306 490226
rect 453374 490170 453430 490226
rect 453498 490170 453554 490226
rect 453622 490170 453678 490226
rect 453250 490046 453306 490102
rect 453374 490046 453430 490102
rect 453498 490046 453554 490102
rect 453622 490046 453678 490102
rect 453250 489922 453306 489978
rect 453374 489922 453430 489978
rect 453498 489922 453554 489978
rect 453622 489922 453678 489978
rect 453250 472294 453306 472350
rect 453374 472294 453430 472350
rect 453498 472294 453554 472350
rect 453622 472294 453678 472350
rect 453250 472170 453306 472226
rect 453374 472170 453430 472226
rect 453498 472170 453554 472226
rect 453622 472170 453678 472226
rect 453250 472046 453306 472102
rect 453374 472046 453430 472102
rect 453498 472046 453554 472102
rect 453622 472046 453678 472102
rect 453250 471922 453306 471978
rect 453374 471922 453430 471978
rect 453498 471922 453554 471978
rect 453622 471922 453678 471978
rect 453250 454294 453306 454350
rect 453374 454294 453430 454350
rect 453498 454294 453554 454350
rect 453622 454294 453678 454350
rect 453250 454170 453306 454226
rect 453374 454170 453430 454226
rect 453498 454170 453554 454226
rect 453622 454170 453678 454226
rect 453250 454046 453306 454102
rect 453374 454046 453430 454102
rect 453498 454046 453554 454102
rect 453622 454046 453678 454102
rect 453250 453922 453306 453978
rect 453374 453922 453430 453978
rect 453498 453922 453554 453978
rect 453622 453922 453678 453978
rect 453250 436294 453306 436350
rect 453374 436294 453430 436350
rect 453498 436294 453554 436350
rect 453622 436294 453678 436350
rect 453250 436170 453306 436226
rect 453374 436170 453430 436226
rect 453498 436170 453554 436226
rect 453622 436170 453678 436226
rect 453250 436046 453306 436102
rect 453374 436046 453430 436102
rect 453498 436046 453554 436102
rect 453622 436046 453678 436102
rect 453250 435922 453306 435978
rect 453374 435922 453430 435978
rect 453498 435922 453554 435978
rect 453622 435922 453678 435978
rect 453250 418294 453306 418350
rect 453374 418294 453430 418350
rect 453498 418294 453554 418350
rect 453622 418294 453678 418350
rect 453250 418170 453306 418226
rect 453374 418170 453430 418226
rect 453498 418170 453554 418226
rect 453622 418170 453678 418226
rect 453250 418046 453306 418102
rect 453374 418046 453430 418102
rect 453498 418046 453554 418102
rect 453622 418046 453678 418102
rect 453250 417922 453306 417978
rect 453374 417922 453430 417978
rect 453498 417922 453554 417978
rect 453622 417922 453678 417978
rect 453250 400294 453306 400350
rect 453374 400294 453430 400350
rect 453498 400294 453554 400350
rect 453622 400294 453678 400350
rect 453250 400170 453306 400226
rect 453374 400170 453430 400226
rect 453498 400170 453554 400226
rect 453622 400170 453678 400226
rect 453250 400046 453306 400102
rect 453374 400046 453430 400102
rect 453498 400046 453554 400102
rect 453622 400046 453678 400102
rect 453250 399922 453306 399978
rect 453374 399922 453430 399978
rect 453498 399922 453554 399978
rect 453622 399922 453678 399978
rect 453250 382294 453306 382350
rect 453374 382294 453430 382350
rect 453498 382294 453554 382350
rect 453622 382294 453678 382350
rect 453250 382170 453306 382226
rect 453374 382170 453430 382226
rect 453498 382170 453554 382226
rect 453622 382170 453678 382226
rect 453250 382046 453306 382102
rect 453374 382046 453430 382102
rect 453498 382046 453554 382102
rect 453622 382046 453678 382102
rect 453250 381922 453306 381978
rect 453374 381922 453430 381978
rect 453498 381922 453554 381978
rect 453622 381922 453678 381978
rect 453250 364294 453306 364350
rect 453374 364294 453430 364350
rect 453498 364294 453554 364350
rect 453622 364294 453678 364350
rect 453250 364170 453306 364226
rect 453374 364170 453430 364226
rect 453498 364170 453554 364226
rect 453622 364170 453678 364226
rect 453250 364046 453306 364102
rect 453374 364046 453430 364102
rect 453498 364046 453554 364102
rect 453622 364046 453678 364102
rect 453250 363922 453306 363978
rect 453374 363922 453430 363978
rect 453498 363922 453554 363978
rect 453622 363922 453678 363978
rect 453250 346294 453306 346350
rect 453374 346294 453430 346350
rect 453498 346294 453554 346350
rect 453622 346294 453678 346350
rect 453250 346170 453306 346226
rect 453374 346170 453430 346226
rect 453498 346170 453554 346226
rect 453622 346170 453678 346226
rect 453250 346046 453306 346102
rect 453374 346046 453430 346102
rect 453498 346046 453554 346102
rect 453622 346046 453678 346102
rect 453250 345922 453306 345978
rect 453374 345922 453430 345978
rect 453498 345922 453554 345978
rect 453622 345922 453678 345978
rect 453250 328294 453306 328350
rect 453374 328294 453430 328350
rect 453498 328294 453554 328350
rect 453622 328294 453678 328350
rect 453250 328170 453306 328226
rect 453374 328170 453430 328226
rect 453498 328170 453554 328226
rect 453622 328170 453678 328226
rect 453250 328046 453306 328102
rect 453374 328046 453430 328102
rect 453498 328046 453554 328102
rect 453622 328046 453678 328102
rect 453250 327922 453306 327978
rect 453374 327922 453430 327978
rect 453498 327922 453554 327978
rect 453622 327922 453678 327978
rect 453250 310294 453306 310350
rect 453374 310294 453430 310350
rect 453498 310294 453554 310350
rect 453622 310294 453678 310350
rect 453250 310170 453306 310226
rect 453374 310170 453430 310226
rect 453498 310170 453554 310226
rect 453622 310170 453678 310226
rect 453250 310046 453306 310102
rect 453374 310046 453430 310102
rect 453498 310046 453554 310102
rect 453622 310046 453678 310102
rect 453250 309922 453306 309978
rect 453374 309922 453430 309978
rect 453498 309922 453554 309978
rect 453622 309922 453678 309978
rect 453250 292294 453306 292350
rect 453374 292294 453430 292350
rect 453498 292294 453554 292350
rect 453622 292294 453678 292350
rect 453250 292170 453306 292226
rect 453374 292170 453430 292226
rect 453498 292170 453554 292226
rect 453622 292170 453678 292226
rect 453250 292046 453306 292102
rect 453374 292046 453430 292102
rect 453498 292046 453554 292102
rect 453622 292046 453678 292102
rect 453250 291922 453306 291978
rect 453374 291922 453430 291978
rect 453498 291922 453554 291978
rect 453622 291922 453678 291978
rect 453250 274294 453306 274350
rect 453374 274294 453430 274350
rect 453498 274294 453554 274350
rect 453622 274294 453678 274350
rect 453250 274170 453306 274226
rect 453374 274170 453430 274226
rect 453498 274170 453554 274226
rect 453622 274170 453678 274226
rect 453250 274046 453306 274102
rect 453374 274046 453430 274102
rect 453498 274046 453554 274102
rect 453622 274046 453678 274102
rect 453250 273922 453306 273978
rect 453374 273922 453430 273978
rect 453498 273922 453554 273978
rect 453622 273922 453678 273978
rect 453250 256294 453306 256350
rect 453374 256294 453430 256350
rect 453498 256294 453554 256350
rect 453622 256294 453678 256350
rect 453250 256170 453306 256226
rect 453374 256170 453430 256226
rect 453498 256170 453554 256226
rect 453622 256170 453678 256226
rect 453250 256046 453306 256102
rect 453374 256046 453430 256102
rect 453498 256046 453554 256102
rect 453622 256046 453678 256102
rect 453250 255922 453306 255978
rect 453374 255922 453430 255978
rect 453498 255922 453554 255978
rect 453622 255922 453678 255978
rect 453250 238294 453306 238350
rect 453374 238294 453430 238350
rect 453498 238294 453554 238350
rect 453622 238294 453678 238350
rect 453250 238170 453306 238226
rect 453374 238170 453430 238226
rect 453498 238170 453554 238226
rect 453622 238170 453678 238226
rect 453250 238046 453306 238102
rect 453374 238046 453430 238102
rect 453498 238046 453554 238102
rect 453622 238046 453678 238102
rect 453250 237922 453306 237978
rect 453374 237922 453430 237978
rect 453498 237922 453554 237978
rect 453622 237922 453678 237978
rect 453250 220294 453306 220350
rect 453374 220294 453430 220350
rect 453498 220294 453554 220350
rect 453622 220294 453678 220350
rect 453250 220170 453306 220226
rect 453374 220170 453430 220226
rect 453498 220170 453554 220226
rect 453622 220170 453678 220226
rect 453250 220046 453306 220102
rect 453374 220046 453430 220102
rect 453498 220046 453554 220102
rect 453622 220046 453678 220102
rect 453250 219922 453306 219978
rect 453374 219922 453430 219978
rect 453498 219922 453554 219978
rect 453622 219922 453678 219978
rect 456970 598116 457026 598172
rect 457094 598116 457150 598172
rect 457218 598116 457274 598172
rect 457342 598116 457398 598172
rect 456970 597992 457026 598048
rect 457094 597992 457150 598048
rect 457218 597992 457274 598048
rect 457342 597992 457398 598048
rect 456970 597868 457026 597924
rect 457094 597868 457150 597924
rect 457218 597868 457274 597924
rect 457342 597868 457398 597924
rect 456970 597744 457026 597800
rect 457094 597744 457150 597800
rect 457218 597744 457274 597800
rect 457342 597744 457398 597800
rect 456970 586294 457026 586350
rect 457094 586294 457150 586350
rect 457218 586294 457274 586350
rect 457342 586294 457398 586350
rect 456970 586170 457026 586226
rect 457094 586170 457150 586226
rect 457218 586170 457274 586226
rect 457342 586170 457398 586226
rect 456970 586046 457026 586102
rect 457094 586046 457150 586102
rect 457218 586046 457274 586102
rect 457342 586046 457398 586102
rect 456970 585922 457026 585978
rect 457094 585922 457150 585978
rect 457218 585922 457274 585978
rect 457342 585922 457398 585978
rect 456970 568294 457026 568350
rect 457094 568294 457150 568350
rect 457218 568294 457274 568350
rect 457342 568294 457398 568350
rect 456970 568170 457026 568226
rect 457094 568170 457150 568226
rect 457218 568170 457274 568226
rect 457342 568170 457398 568226
rect 456970 568046 457026 568102
rect 457094 568046 457150 568102
rect 457218 568046 457274 568102
rect 457342 568046 457398 568102
rect 456970 567922 457026 567978
rect 457094 567922 457150 567978
rect 457218 567922 457274 567978
rect 457342 567922 457398 567978
rect 456970 550294 457026 550350
rect 457094 550294 457150 550350
rect 457218 550294 457274 550350
rect 457342 550294 457398 550350
rect 456970 550170 457026 550226
rect 457094 550170 457150 550226
rect 457218 550170 457274 550226
rect 457342 550170 457398 550226
rect 456970 550046 457026 550102
rect 457094 550046 457150 550102
rect 457218 550046 457274 550102
rect 457342 550046 457398 550102
rect 456970 549922 457026 549978
rect 457094 549922 457150 549978
rect 457218 549922 457274 549978
rect 457342 549922 457398 549978
rect 456970 532294 457026 532350
rect 457094 532294 457150 532350
rect 457218 532294 457274 532350
rect 457342 532294 457398 532350
rect 456970 532170 457026 532226
rect 457094 532170 457150 532226
rect 457218 532170 457274 532226
rect 457342 532170 457398 532226
rect 456970 532046 457026 532102
rect 457094 532046 457150 532102
rect 457218 532046 457274 532102
rect 457342 532046 457398 532102
rect 456970 531922 457026 531978
rect 457094 531922 457150 531978
rect 457218 531922 457274 531978
rect 457342 531922 457398 531978
rect 456970 514294 457026 514350
rect 457094 514294 457150 514350
rect 457218 514294 457274 514350
rect 457342 514294 457398 514350
rect 456970 514170 457026 514226
rect 457094 514170 457150 514226
rect 457218 514170 457274 514226
rect 457342 514170 457398 514226
rect 456970 514046 457026 514102
rect 457094 514046 457150 514102
rect 457218 514046 457274 514102
rect 457342 514046 457398 514102
rect 456970 513922 457026 513978
rect 457094 513922 457150 513978
rect 457218 513922 457274 513978
rect 457342 513922 457398 513978
rect 456970 496294 457026 496350
rect 457094 496294 457150 496350
rect 457218 496294 457274 496350
rect 457342 496294 457398 496350
rect 456970 496170 457026 496226
rect 457094 496170 457150 496226
rect 457218 496170 457274 496226
rect 457342 496170 457398 496226
rect 456970 496046 457026 496102
rect 457094 496046 457150 496102
rect 457218 496046 457274 496102
rect 457342 496046 457398 496102
rect 456970 495922 457026 495978
rect 457094 495922 457150 495978
rect 457218 495922 457274 495978
rect 457342 495922 457398 495978
rect 456970 478294 457026 478350
rect 457094 478294 457150 478350
rect 457218 478294 457274 478350
rect 457342 478294 457398 478350
rect 456970 478170 457026 478226
rect 457094 478170 457150 478226
rect 457218 478170 457274 478226
rect 457342 478170 457398 478226
rect 456970 478046 457026 478102
rect 457094 478046 457150 478102
rect 457218 478046 457274 478102
rect 457342 478046 457398 478102
rect 456970 477922 457026 477978
rect 457094 477922 457150 477978
rect 457218 477922 457274 477978
rect 457342 477922 457398 477978
rect 456970 460294 457026 460350
rect 457094 460294 457150 460350
rect 457218 460294 457274 460350
rect 457342 460294 457398 460350
rect 456970 460170 457026 460226
rect 457094 460170 457150 460226
rect 457218 460170 457274 460226
rect 457342 460170 457398 460226
rect 456970 460046 457026 460102
rect 457094 460046 457150 460102
rect 457218 460046 457274 460102
rect 457342 460046 457398 460102
rect 456970 459922 457026 459978
rect 457094 459922 457150 459978
rect 457218 459922 457274 459978
rect 457342 459922 457398 459978
rect 456970 442294 457026 442350
rect 457094 442294 457150 442350
rect 457218 442294 457274 442350
rect 457342 442294 457398 442350
rect 456970 442170 457026 442226
rect 457094 442170 457150 442226
rect 457218 442170 457274 442226
rect 457342 442170 457398 442226
rect 456970 442046 457026 442102
rect 457094 442046 457150 442102
rect 457218 442046 457274 442102
rect 457342 442046 457398 442102
rect 456970 441922 457026 441978
rect 457094 441922 457150 441978
rect 457218 441922 457274 441978
rect 457342 441922 457398 441978
rect 456970 424294 457026 424350
rect 457094 424294 457150 424350
rect 457218 424294 457274 424350
rect 457342 424294 457398 424350
rect 456970 424170 457026 424226
rect 457094 424170 457150 424226
rect 457218 424170 457274 424226
rect 457342 424170 457398 424226
rect 456970 424046 457026 424102
rect 457094 424046 457150 424102
rect 457218 424046 457274 424102
rect 457342 424046 457398 424102
rect 456970 423922 457026 423978
rect 457094 423922 457150 423978
rect 457218 423922 457274 423978
rect 457342 423922 457398 423978
rect 456970 406294 457026 406350
rect 457094 406294 457150 406350
rect 457218 406294 457274 406350
rect 457342 406294 457398 406350
rect 456970 406170 457026 406226
rect 457094 406170 457150 406226
rect 457218 406170 457274 406226
rect 457342 406170 457398 406226
rect 456970 406046 457026 406102
rect 457094 406046 457150 406102
rect 457218 406046 457274 406102
rect 457342 406046 457398 406102
rect 456970 405922 457026 405978
rect 457094 405922 457150 405978
rect 457218 405922 457274 405978
rect 457342 405922 457398 405978
rect 456970 388294 457026 388350
rect 457094 388294 457150 388350
rect 457218 388294 457274 388350
rect 457342 388294 457398 388350
rect 456970 388170 457026 388226
rect 457094 388170 457150 388226
rect 457218 388170 457274 388226
rect 457342 388170 457398 388226
rect 456970 388046 457026 388102
rect 457094 388046 457150 388102
rect 457218 388046 457274 388102
rect 457342 388046 457398 388102
rect 456970 387922 457026 387978
rect 457094 387922 457150 387978
rect 457218 387922 457274 387978
rect 457342 387922 457398 387978
rect 456970 370294 457026 370350
rect 457094 370294 457150 370350
rect 457218 370294 457274 370350
rect 457342 370294 457398 370350
rect 456970 370170 457026 370226
rect 457094 370170 457150 370226
rect 457218 370170 457274 370226
rect 457342 370170 457398 370226
rect 456970 370046 457026 370102
rect 457094 370046 457150 370102
rect 457218 370046 457274 370102
rect 457342 370046 457398 370102
rect 456970 369922 457026 369978
rect 457094 369922 457150 369978
rect 457218 369922 457274 369978
rect 457342 369922 457398 369978
rect 456970 352294 457026 352350
rect 457094 352294 457150 352350
rect 457218 352294 457274 352350
rect 457342 352294 457398 352350
rect 456970 352170 457026 352226
rect 457094 352170 457150 352226
rect 457218 352170 457274 352226
rect 457342 352170 457398 352226
rect 456970 352046 457026 352102
rect 457094 352046 457150 352102
rect 457218 352046 457274 352102
rect 457342 352046 457398 352102
rect 456970 351922 457026 351978
rect 457094 351922 457150 351978
rect 457218 351922 457274 351978
rect 457342 351922 457398 351978
rect 456970 334294 457026 334350
rect 457094 334294 457150 334350
rect 457218 334294 457274 334350
rect 457342 334294 457398 334350
rect 456970 334170 457026 334226
rect 457094 334170 457150 334226
rect 457218 334170 457274 334226
rect 457342 334170 457398 334226
rect 456970 334046 457026 334102
rect 457094 334046 457150 334102
rect 457218 334046 457274 334102
rect 457342 334046 457398 334102
rect 456970 333922 457026 333978
rect 457094 333922 457150 333978
rect 457218 333922 457274 333978
rect 457342 333922 457398 333978
rect 456970 316294 457026 316350
rect 457094 316294 457150 316350
rect 457218 316294 457274 316350
rect 457342 316294 457398 316350
rect 456970 316170 457026 316226
rect 457094 316170 457150 316226
rect 457218 316170 457274 316226
rect 457342 316170 457398 316226
rect 456970 316046 457026 316102
rect 457094 316046 457150 316102
rect 457218 316046 457274 316102
rect 457342 316046 457398 316102
rect 456970 315922 457026 315978
rect 457094 315922 457150 315978
rect 457218 315922 457274 315978
rect 457342 315922 457398 315978
rect 456970 298294 457026 298350
rect 457094 298294 457150 298350
rect 457218 298294 457274 298350
rect 457342 298294 457398 298350
rect 456970 298170 457026 298226
rect 457094 298170 457150 298226
rect 457218 298170 457274 298226
rect 457342 298170 457398 298226
rect 456970 298046 457026 298102
rect 457094 298046 457150 298102
rect 457218 298046 457274 298102
rect 457342 298046 457398 298102
rect 456970 297922 457026 297978
rect 457094 297922 457150 297978
rect 457218 297922 457274 297978
rect 457342 297922 457398 297978
rect 456970 280294 457026 280350
rect 457094 280294 457150 280350
rect 457218 280294 457274 280350
rect 457342 280294 457398 280350
rect 456970 280170 457026 280226
rect 457094 280170 457150 280226
rect 457218 280170 457274 280226
rect 457342 280170 457398 280226
rect 456970 280046 457026 280102
rect 457094 280046 457150 280102
rect 457218 280046 457274 280102
rect 457342 280046 457398 280102
rect 456970 279922 457026 279978
rect 457094 279922 457150 279978
rect 457218 279922 457274 279978
rect 457342 279922 457398 279978
rect 456970 262294 457026 262350
rect 457094 262294 457150 262350
rect 457218 262294 457274 262350
rect 457342 262294 457398 262350
rect 456970 262170 457026 262226
rect 457094 262170 457150 262226
rect 457218 262170 457274 262226
rect 457342 262170 457398 262226
rect 456970 262046 457026 262102
rect 457094 262046 457150 262102
rect 457218 262046 457274 262102
rect 457342 262046 457398 262102
rect 456970 261922 457026 261978
rect 457094 261922 457150 261978
rect 457218 261922 457274 261978
rect 457342 261922 457398 261978
rect 456970 244294 457026 244350
rect 457094 244294 457150 244350
rect 457218 244294 457274 244350
rect 457342 244294 457398 244350
rect 456970 244170 457026 244226
rect 457094 244170 457150 244226
rect 457218 244170 457274 244226
rect 457342 244170 457398 244226
rect 456970 244046 457026 244102
rect 457094 244046 457150 244102
rect 457218 244046 457274 244102
rect 457342 244046 457398 244102
rect 456970 243922 457026 243978
rect 457094 243922 457150 243978
rect 457218 243922 457274 243978
rect 457342 243922 457398 243978
rect 456970 226294 457026 226350
rect 457094 226294 457150 226350
rect 457218 226294 457274 226350
rect 457342 226294 457398 226350
rect 456970 226170 457026 226226
rect 457094 226170 457150 226226
rect 457218 226170 457274 226226
rect 457342 226170 457398 226226
rect 456970 226046 457026 226102
rect 457094 226046 457150 226102
rect 457218 226046 457274 226102
rect 457342 226046 457398 226102
rect 456970 225922 457026 225978
rect 457094 225922 457150 225978
rect 457218 225922 457274 225978
rect 457342 225922 457398 225978
rect 471250 597156 471306 597212
rect 471374 597156 471430 597212
rect 471498 597156 471554 597212
rect 471622 597156 471678 597212
rect 471250 597032 471306 597088
rect 471374 597032 471430 597088
rect 471498 597032 471554 597088
rect 471622 597032 471678 597088
rect 471250 596908 471306 596964
rect 471374 596908 471430 596964
rect 471498 596908 471554 596964
rect 471622 596908 471678 596964
rect 471250 596784 471306 596840
rect 471374 596784 471430 596840
rect 471498 596784 471554 596840
rect 471622 596784 471678 596840
rect 489250 597156 489306 597212
rect 489374 597156 489430 597212
rect 489498 597156 489554 597212
rect 489622 597156 489678 597212
rect 489250 597032 489306 597088
rect 489374 597032 489430 597088
rect 489498 597032 489554 597088
rect 489622 597032 489678 597088
rect 489250 596908 489306 596964
rect 489374 596908 489430 596964
rect 489498 596908 489554 596964
rect 489622 596908 489678 596964
rect 489250 596784 489306 596840
rect 489374 596784 489430 596840
rect 489498 596784 489554 596840
rect 489622 596784 489678 596840
rect 471250 580294 471306 580350
rect 471374 580294 471430 580350
rect 471498 580294 471554 580350
rect 471622 580294 471678 580350
rect 471250 580170 471306 580226
rect 471374 580170 471430 580226
rect 471498 580170 471554 580226
rect 471622 580170 471678 580226
rect 471250 580046 471306 580102
rect 471374 580046 471430 580102
rect 471498 580046 471554 580102
rect 471622 580046 471678 580102
rect 471250 579922 471306 579978
rect 471374 579922 471430 579978
rect 471498 579922 471554 579978
rect 471622 579922 471678 579978
rect 471250 562294 471306 562350
rect 471374 562294 471430 562350
rect 471498 562294 471554 562350
rect 471622 562294 471678 562350
rect 471250 562170 471306 562226
rect 471374 562170 471430 562226
rect 471498 562170 471554 562226
rect 471622 562170 471678 562226
rect 471250 562046 471306 562102
rect 471374 562046 471430 562102
rect 471498 562046 471554 562102
rect 471622 562046 471678 562102
rect 471250 561922 471306 561978
rect 471374 561922 471430 561978
rect 471498 561922 471554 561978
rect 471622 561922 471678 561978
rect 471250 544294 471306 544350
rect 471374 544294 471430 544350
rect 471498 544294 471554 544350
rect 471622 544294 471678 544350
rect 471250 544170 471306 544226
rect 471374 544170 471430 544226
rect 471498 544170 471554 544226
rect 471622 544170 471678 544226
rect 471250 544046 471306 544102
rect 471374 544046 471430 544102
rect 471498 544046 471554 544102
rect 471622 544046 471678 544102
rect 471250 543922 471306 543978
rect 471374 543922 471430 543978
rect 471498 543922 471554 543978
rect 471622 543922 471678 543978
rect 471250 526294 471306 526350
rect 471374 526294 471430 526350
rect 471498 526294 471554 526350
rect 471622 526294 471678 526350
rect 471250 526170 471306 526226
rect 471374 526170 471430 526226
rect 471498 526170 471554 526226
rect 471622 526170 471678 526226
rect 471250 526046 471306 526102
rect 471374 526046 471430 526102
rect 471498 526046 471554 526102
rect 471622 526046 471678 526102
rect 471250 525922 471306 525978
rect 471374 525922 471430 525978
rect 471498 525922 471554 525978
rect 471622 525922 471678 525978
rect 471250 508294 471306 508350
rect 471374 508294 471430 508350
rect 471498 508294 471554 508350
rect 471622 508294 471678 508350
rect 471250 508170 471306 508226
rect 471374 508170 471430 508226
rect 471498 508170 471554 508226
rect 471622 508170 471678 508226
rect 471250 508046 471306 508102
rect 471374 508046 471430 508102
rect 471498 508046 471554 508102
rect 471622 508046 471678 508102
rect 471250 507922 471306 507978
rect 471374 507922 471430 507978
rect 471498 507922 471554 507978
rect 471622 507922 471678 507978
rect 471250 490294 471306 490350
rect 471374 490294 471430 490350
rect 471498 490294 471554 490350
rect 471622 490294 471678 490350
rect 471250 490170 471306 490226
rect 471374 490170 471430 490226
rect 471498 490170 471554 490226
rect 471622 490170 471678 490226
rect 471250 490046 471306 490102
rect 471374 490046 471430 490102
rect 471498 490046 471554 490102
rect 471622 490046 471678 490102
rect 471250 489922 471306 489978
rect 471374 489922 471430 489978
rect 471498 489922 471554 489978
rect 471622 489922 471678 489978
rect 471250 472294 471306 472350
rect 471374 472294 471430 472350
rect 471498 472294 471554 472350
rect 471622 472294 471678 472350
rect 471250 472170 471306 472226
rect 471374 472170 471430 472226
rect 471498 472170 471554 472226
rect 471622 472170 471678 472226
rect 471250 472046 471306 472102
rect 471374 472046 471430 472102
rect 471498 472046 471554 472102
rect 471622 472046 471678 472102
rect 471250 471922 471306 471978
rect 471374 471922 471430 471978
rect 471498 471922 471554 471978
rect 471622 471922 471678 471978
rect 471250 454294 471306 454350
rect 471374 454294 471430 454350
rect 471498 454294 471554 454350
rect 471622 454294 471678 454350
rect 471250 454170 471306 454226
rect 471374 454170 471430 454226
rect 471498 454170 471554 454226
rect 471622 454170 471678 454226
rect 471250 454046 471306 454102
rect 471374 454046 471430 454102
rect 471498 454046 471554 454102
rect 471622 454046 471678 454102
rect 471250 453922 471306 453978
rect 471374 453922 471430 453978
rect 471498 453922 471554 453978
rect 471622 453922 471678 453978
rect 471250 436294 471306 436350
rect 471374 436294 471430 436350
rect 471498 436294 471554 436350
rect 471622 436294 471678 436350
rect 471250 436170 471306 436226
rect 471374 436170 471430 436226
rect 471498 436170 471554 436226
rect 471622 436170 471678 436226
rect 471250 436046 471306 436102
rect 471374 436046 471430 436102
rect 471498 436046 471554 436102
rect 471622 436046 471678 436102
rect 471250 435922 471306 435978
rect 471374 435922 471430 435978
rect 471498 435922 471554 435978
rect 471622 435922 471678 435978
rect 471250 418294 471306 418350
rect 471374 418294 471430 418350
rect 471498 418294 471554 418350
rect 471622 418294 471678 418350
rect 471250 418170 471306 418226
rect 471374 418170 471430 418226
rect 471498 418170 471554 418226
rect 471622 418170 471678 418226
rect 471250 418046 471306 418102
rect 471374 418046 471430 418102
rect 471498 418046 471554 418102
rect 471622 418046 471678 418102
rect 471250 417922 471306 417978
rect 471374 417922 471430 417978
rect 471498 417922 471554 417978
rect 471622 417922 471678 417978
rect 471250 400294 471306 400350
rect 471374 400294 471430 400350
rect 471498 400294 471554 400350
rect 471622 400294 471678 400350
rect 471250 400170 471306 400226
rect 471374 400170 471430 400226
rect 471498 400170 471554 400226
rect 471622 400170 471678 400226
rect 471250 400046 471306 400102
rect 471374 400046 471430 400102
rect 471498 400046 471554 400102
rect 471622 400046 471678 400102
rect 471250 399922 471306 399978
rect 471374 399922 471430 399978
rect 471498 399922 471554 399978
rect 471622 399922 471678 399978
rect 471250 382294 471306 382350
rect 471374 382294 471430 382350
rect 471498 382294 471554 382350
rect 471622 382294 471678 382350
rect 471250 382170 471306 382226
rect 471374 382170 471430 382226
rect 471498 382170 471554 382226
rect 471622 382170 471678 382226
rect 471250 382046 471306 382102
rect 471374 382046 471430 382102
rect 471498 382046 471554 382102
rect 471622 382046 471678 382102
rect 471250 381922 471306 381978
rect 471374 381922 471430 381978
rect 471498 381922 471554 381978
rect 471622 381922 471678 381978
rect 471250 364294 471306 364350
rect 471374 364294 471430 364350
rect 471498 364294 471554 364350
rect 471622 364294 471678 364350
rect 471250 364170 471306 364226
rect 471374 364170 471430 364226
rect 471498 364170 471554 364226
rect 471622 364170 471678 364226
rect 471250 364046 471306 364102
rect 471374 364046 471430 364102
rect 471498 364046 471554 364102
rect 471622 364046 471678 364102
rect 471250 363922 471306 363978
rect 471374 363922 471430 363978
rect 471498 363922 471554 363978
rect 471622 363922 471678 363978
rect 471250 346294 471306 346350
rect 471374 346294 471430 346350
rect 471498 346294 471554 346350
rect 471622 346294 471678 346350
rect 471250 346170 471306 346226
rect 471374 346170 471430 346226
rect 471498 346170 471554 346226
rect 471622 346170 471678 346226
rect 471250 346046 471306 346102
rect 471374 346046 471430 346102
rect 471498 346046 471554 346102
rect 471622 346046 471678 346102
rect 471250 345922 471306 345978
rect 471374 345922 471430 345978
rect 471498 345922 471554 345978
rect 471622 345922 471678 345978
rect 471250 328294 471306 328350
rect 471374 328294 471430 328350
rect 471498 328294 471554 328350
rect 471622 328294 471678 328350
rect 471250 328170 471306 328226
rect 471374 328170 471430 328226
rect 471498 328170 471554 328226
rect 471622 328170 471678 328226
rect 471250 328046 471306 328102
rect 471374 328046 471430 328102
rect 471498 328046 471554 328102
rect 471622 328046 471678 328102
rect 471250 327922 471306 327978
rect 471374 327922 471430 327978
rect 471498 327922 471554 327978
rect 471622 327922 471678 327978
rect 471250 310294 471306 310350
rect 471374 310294 471430 310350
rect 471498 310294 471554 310350
rect 471622 310294 471678 310350
rect 471250 310170 471306 310226
rect 471374 310170 471430 310226
rect 471498 310170 471554 310226
rect 471622 310170 471678 310226
rect 471250 310046 471306 310102
rect 471374 310046 471430 310102
rect 471498 310046 471554 310102
rect 471622 310046 471678 310102
rect 471250 309922 471306 309978
rect 471374 309922 471430 309978
rect 471498 309922 471554 309978
rect 471622 309922 471678 309978
rect 471250 292294 471306 292350
rect 471374 292294 471430 292350
rect 471498 292294 471554 292350
rect 471622 292294 471678 292350
rect 471250 292170 471306 292226
rect 471374 292170 471430 292226
rect 471498 292170 471554 292226
rect 471622 292170 471678 292226
rect 471250 292046 471306 292102
rect 471374 292046 471430 292102
rect 471498 292046 471554 292102
rect 471622 292046 471678 292102
rect 471250 291922 471306 291978
rect 471374 291922 471430 291978
rect 471498 291922 471554 291978
rect 471622 291922 471678 291978
rect 471250 274294 471306 274350
rect 471374 274294 471430 274350
rect 471498 274294 471554 274350
rect 471622 274294 471678 274350
rect 471250 274170 471306 274226
rect 471374 274170 471430 274226
rect 471498 274170 471554 274226
rect 471622 274170 471678 274226
rect 471250 274046 471306 274102
rect 471374 274046 471430 274102
rect 471498 274046 471554 274102
rect 471622 274046 471678 274102
rect 471250 273922 471306 273978
rect 471374 273922 471430 273978
rect 471498 273922 471554 273978
rect 471622 273922 471678 273978
rect 471250 256294 471306 256350
rect 471374 256294 471430 256350
rect 471498 256294 471554 256350
rect 471622 256294 471678 256350
rect 471250 256170 471306 256226
rect 471374 256170 471430 256226
rect 471498 256170 471554 256226
rect 471622 256170 471678 256226
rect 471250 256046 471306 256102
rect 471374 256046 471430 256102
rect 471498 256046 471554 256102
rect 471622 256046 471678 256102
rect 471250 255922 471306 255978
rect 471374 255922 471430 255978
rect 471498 255922 471554 255978
rect 471622 255922 471678 255978
rect 471250 238294 471306 238350
rect 471374 238294 471430 238350
rect 471498 238294 471554 238350
rect 471622 238294 471678 238350
rect 471250 238170 471306 238226
rect 471374 238170 471430 238226
rect 471498 238170 471554 238226
rect 471622 238170 471678 238226
rect 471250 238046 471306 238102
rect 471374 238046 471430 238102
rect 471498 238046 471554 238102
rect 471622 238046 471678 238102
rect 471250 237922 471306 237978
rect 471374 237922 471430 237978
rect 471498 237922 471554 237978
rect 471622 237922 471678 237978
rect 471250 220294 471306 220350
rect 471374 220294 471430 220350
rect 471498 220294 471554 220350
rect 471622 220294 471678 220350
rect 471250 220170 471306 220226
rect 471374 220170 471430 220226
rect 471498 220170 471554 220226
rect 471622 220170 471678 220226
rect 471250 220046 471306 220102
rect 471374 220046 471430 220102
rect 471498 220046 471554 220102
rect 471622 220046 471678 220102
rect 471250 219922 471306 219978
rect 471374 219922 471430 219978
rect 471498 219922 471554 219978
rect 471622 219922 471678 219978
rect 489250 580294 489306 580350
rect 489374 580294 489430 580350
rect 489498 580294 489554 580350
rect 489622 580294 489678 580350
rect 489250 580170 489306 580226
rect 489374 580170 489430 580226
rect 489498 580170 489554 580226
rect 489622 580170 489678 580226
rect 489250 580046 489306 580102
rect 489374 580046 489430 580102
rect 489498 580046 489554 580102
rect 489622 580046 489678 580102
rect 489250 579922 489306 579978
rect 489374 579922 489430 579978
rect 489498 579922 489554 579978
rect 489622 579922 489678 579978
rect 489250 562294 489306 562350
rect 489374 562294 489430 562350
rect 489498 562294 489554 562350
rect 489622 562294 489678 562350
rect 489250 562170 489306 562226
rect 489374 562170 489430 562226
rect 489498 562170 489554 562226
rect 489622 562170 489678 562226
rect 489250 562046 489306 562102
rect 489374 562046 489430 562102
rect 489498 562046 489554 562102
rect 489622 562046 489678 562102
rect 489250 561922 489306 561978
rect 489374 561922 489430 561978
rect 489498 561922 489554 561978
rect 489622 561922 489678 561978
rect 489250 544294 489306 544350
rect 489374 544294 489430 544350
rect 489498 544294 489554 544350
rect 489622 544294 489678 544350
rect 489250 544170 489306 544226
rect 489374 544170 489430 544226
rect 489498 544170 489554 544226
rect 489622 544170 489678 544226
rect 489250 544046 489306 544102
rect 489374 544046 489430 544102
rect 489498 544046 489554 544102
rect 489622 544046 489678 544102
rect 489250 543922 489306 543978
rect 489374 543922 489430 543978
rect 489498 543922 489554 543978
rect 489622 543922 489678 543978
rect 489250 526294 489306 526350
rect 489374 526294 489430 526350
rect 489498 526294 489554 526350
rect 489622 526294 489678 526350
rect 489250 526170 489306 526226
rect 489374 526170 489430 526226
rect 489498 526170 489554 526226
rect 489622 526170 489678 526226
rect 489250 526046 489306 526102
rect 489374 526046 489430 526102
rect 489498 526046 489554 526102
rect 489622 526046 489678 526102
rect 489250 525922 489306 525978
rect 489374 525922 489430 525978
rect 489498 525922 489554 525978
rect 489622 525922 489678 525978
rect 489250 508294 489306 508350
rect 489374 508294 489430 508350
rect 489498 508294 489554 508350
rect 489622 508294 489678 508350
rect 489250 508170 489306 508226
rect 489374 508170 489430 508226
rect 489498 508170 489554 508226
rect 489622 508170 489678 508226
rect 489250 508046 489306 508102
rect 489374 508046 489430 508102
rect 489498 508046 489554 508102
rect 489622 508046 489678 508102
rect 489250 507922 489306 507978
rect 489374 507922 489430 507978
rect 489498 507922 489554 507978
rect 489622 507922 489678 507978
rect 489250 490294 489306 490350
rect 489374 490294 489430 490350
rect 489498 490294 489554 490350
rect 489622 490294 489678 490350
rect 489250 490170 489306 490226
rect 489374 490170 489430 490226
rect 489498 490170 489554 490226
rect 489622 490170 489678 490226
rect 489250 490046 489306 490102
rect 489374 490046 489430 490102
rect 489498 490046 489554 490102
rect 489622 490046 489678 490102
rect 489250 489922 489306 489978
rect 489374 489922 489430 489978
rect 489498 489922 489554 489978
rect 489622 489922 489678 489978
rect 489250 472294 489306 472350
rect 489374 472294 489430 472350
rect 489498 472294 489554 472350
rect 489622 472294 489678 472350
rect 489250 472170 489306 472226
rect 489374 472170 489430 472226
rect 489498 472170 489554 472226
rect 489622 472170 489678 472226
rect 489250 472046 489306 472102
rect 489374 472046 489430 472102
rect 489498 472046 489554 472102
rect 489622 472046 489678 472102
rect 489250 471922 489306 471978
rect 489374 471922 489430 471978
rect 489498 471922 489554 471978
rect 489622 471922 489678 471978
rect 489250 454294 489306 454350
rect 489374 454294 489430 454350
rect 489498 454294 489554 454350
rect 489622 454294 489678 454350
rect 489250 454170 489306 454226
rect 489374 454170 489430 454226
rect 489498 454170 489554 454226
rect 489622 454170 489678 454226
rect 489250 454046 489306 454102
rect 489374 454046 489430 454102
rect 489498 454046 489554 454102
rect 489622 454046 489678 454102
rect 489250 453922 489306 453978
rect 489374 453922 489430 453978
rect 489498 453922 489554 453978
rect 489622 453922 489678 453978
rect 489250 436294 489306 436350
rect 489374 436294 489430 436350
rect 489498 436294 489554 436350
rect 489622 436294 489678 436350
rect 489250 436170 489306 436226
rect 489374 436170 489430 436226
rect 489498 436170 489554 436226
rect 489622 436170 489678 436226
rect 489250 436046 489306 436102
rect 489374 436046 489430 436102
rect 489498 436046 489554 436102
rect 489622 436046 489678 436102
rect 489250 435922 489306 435978
rect 489374 435922 489430 435978
rect 489498 435922 489554 435978
rect 489622 435922 489678 435978
rect 489250 418294 489306 418350
rect 489374 418294 489430 418350
rect 489498 418294 489554 418350
rect 489622 418294 489678 418350
rect 489250 418170 489306 418226
rect 489374 418170 489430 418226
rect 489498 418170 489554 418226
rect 489622 418170 489678 418226
rect 489250 418046 489306 418102
rect 489374 418046 489430 418102
rect 489498 418046 489554 418102
rect 489622 418046 489678 418102
rect 489250 417922 489306 417978
rect 489374 417922 489430 417978
rect 489498 417922 489554 417978
rect 489622 417922 489678 417978
rect 489250 400294 489306 400350
rect 489374 400294 489430 400350
rect 489498 400294 489554 400350
rect 489622 400294 489678 400350
rect 489250 400170 489306 400226
rect 489374 400170 489430 400226
rect 489498 400170 489554 400226
rect 489622 400170 489678 400226
rect 489250 400046 489306 400102
rect 489374 400046 489430 400102
rect 489498 400046 489554 400102
rect 489622 400046 489678 400102
rect 489250 399922 489306 399978
rect 489374 399922 489430 399978
rect 489498 399922 489554 399978
rect 489622 399922 489678 399978
rect 489250 382294 489306 382350
rect 489374 382294 489430 382350
rect 489498 382294 489554 382350
rect 489622 382294 489678 382350
rect 489250 382170 489306 382226
rect 489374 382170 489430 382226
rect 489498 382170 489554 382226
rect 489622 382170 489678 382226
rect 489250 382046 489306 382102
rect 489374 382046 489430 382102
rect 489498 382046 489554 382102
rect 489622 382046 489678 382102
rect 489250 381922 489306 381978
rect 489374 381922 489430 381978
rect 489498 381922 489554 381978
rect 489622 381922 489678 381978
rect 489250 364294 489306 364350
rect 489374 364294 489430 364350
rect 489498 364294 489554 364350
rect 489622 364294 489678 364350
rect 489250 364170 489306 364226
rect 489374 364170 489430 364226
rect 489498 364170 489554 364226
rect 489622 364170 489678 364226
rect 489250 364046 489306 364102
rect 489374 364046 489430 364102
rect 489498 364046 489554 364102
rect 489622 364046 489678 364102
rect 489250 363922 489306 363978
rect 489374 363922 489430 363978
rect 489498 363922 489554 363978
rect 489622 363922 489678 363978
rect 489250 346294 489306 346350
rect 489374 346294 489430 346350
rect 489498 346294 489554 346350
rect 489622 346294 489678 346350
rect 489250 346170 489306 346226
rect 489374 346170 489430 346226
rect 489498 346170 489554 346226
rect 489622 346170 489678 346226
rect 489250 346046 489306 346102
rect 489374 346046 489430 346102
rect 489498 346046 489554 346102
rect 489622 346046 489678 346102
rect 489250 345922 489306 345978
rect 489374 345922 489430 345978
rect 489498 345922 489554 345978
rect 489622 345922 489678 345978
rect 489250 328294 489306 328350
rect 489374 328294 489430 328350
rect 489498 328294 489554 328350
rect 489622 328294 489678 328350
rect 489250 328170 489306 328226
rect 489374 328170 489430 328226
rect 489498 328170 489554 328226
rect 489622 328170 489678 328226
rect 489250 328046 489306 328102
rect 489374 328046 489430 328102
rect 489498 328046 489554 328102
rect 489622 328046 489678 328102
rect 489250 327922 489306 327978
rect 489374 327922 489430 327978
rect 489498 327922 489554 327978
rect 489622 327922 489678 327978
rect 489250 310294 489306 310350
rect 489374 310294 489430 310350
rect 489498 310294 489554 310350
rect 489622 310294 489678 310350
rect 489250 310170 489306 310226
rect 489374 310170 489430 310226
rect 489498 310170 489554 310226
rect 489622 310170 489678 310226
rect 489250 310046 489306 310102
rect 489374 310046 489430 310102
rect 489498 310046 489554 310102
rect 489622 310046 489678 310102
rect 489250 309922 489306 309978
rect 489374 309922 489430 309978
rect 489498 309922 489554 309978
rect 489622 309922 489678 309978
rect 489250 292294 489306 292350
rect 489374 292294 489430 292350
rect 489498 292294 489554 292350
rect 489622 292294 489678 292350
rect 489250 292170 489306 292226
rect 489374 292170 489430 292226
rect 489498 292170 489554 292226
rect 489622 292170 489678 292226
rect 489250 292046 489306 292102
rect 489374 292046 489430 292102
rect 489498 292046 489554 292102
rect 489622 292046 489678 292102
rect 489250 291922 489306 291978
rect 489374 291922 489430 291978
rect 489498 291922 489554 291978
rect 489622 291922 489678 291978
rect 489250 274294 489306 274350
rect 489374 274294 489430 274350
rect 489498 274294 489554 274350
rect 489622 274294 489678 274350
rect 489250 274170 489306 274226
rect 489374 274170 489430 274226
rect 489498 274170 489554 274226
rect 489622 274170 489678 274226
rect 489250 274046 489306 274102
rect 489374 274046 489430 274102
rect 489498 274046 489554 274102
rect 489622 274046 489678 274102
rect 489250 273922 489306 273978
rect 489374 273922 489430 273978
rect 489498 273922 489554 273978
rect 489622 273922 489678 273978
rect 489250 256294 489306 256350
rect 489374 256294 489430 256350
rect 489498 256294 489554 256350
rect 489622 256294 489678 256350
rect 489250 256170 489306 256226
rect 489374 256170 489430 256226
rect 489498 256170 489554 256226
rect 489622 256170 489678 256226
rect 489250 256046 489306 256102
rect 489374 256046 489430 256102
rect 489498 256046 489554 256102
rect 489622 256046 489678 256102
rect 489250 255922 489306 255978
rect 489374 255922 489430 255978
rect 489498 255922 489554 255978
rect 489622 255922 489678 255978
rect 489250 238294 489306 238350
rect 489374 238294 489430 238350
rect 489498 238294 489554 238350
rect 489622 238294 489678 238350
rect 489250 238170 489306 238226
rect 489374 238170 489430 238226
rect 489498 238170 489554 238226
rect 489622 238170 489678 238226
rect 489250 238046 489306 238102
rect 489374 238046 489430 238102
rect 489498 238046 489554 238102
rect 489622 238046 489678 238102
rect 489250 237922 489306 237978
rect 489374 237922 489430 237978
rect 489498 237922 489554 237978
rect 489622 237922 489678 237978
rect 489250 220294 489306 220350
rect 489374 220294 489430 220350
rect 489498 220294 489554 220350
rect 489622 220294 489678 220350
rect 489250 220170 489306 220226
rect 489374 220170 489430 220226
rect 489498 220170 489554 220226
rect 489622 220170 489678 220226
rect 489250 220046 489306 220102
rect 489374 220046 489430 220102
rect 489498 220046 489554 220102
rect 489622 220046 489678 220102
rect 489250 219922 489306 219978
rect 489374 219922 489430 219978
rect 489498 219922 489554 219978
rect 489622 219922 489678 219978
rect 492970 598116 493026 598172
rect 493094 598116 493150 598172
rect 493218 598116 493274 598172
rect 493342 598116 493398 598172
rect 492970 597992 493026 598048
rect 493094 597992 493150 598048
rect 493218 597992 493274 598048
rect 493342 597992 493398 598048
rect 492970 597868 493026 597924
rect 493094 597868 493150 597924
rect 493218 597868 493274 597924
rect 493342 597868 493398 597924
rect 492970 597744 493026 597800
rect 493094 597744 493150 597800
rect 493218 597744 493274 597800
rect 493342 597744 493398 597800
rect 492970 586294 493026 586350
rect 493094 586294 493150 586350
rect 493218 586294 493274 586350
rect 493342 586294 493398 586350
rect 492970 586170 493026 586226
rect 493094 586170 493150 586226
rect 493218 586170 493274 586226
rect 493342 586170 493398 586226
rect 492970 586046 493026 586102
rect 493094 586046 493150 586102
rect 493218 586046 493274 586102
rect 493342 586046 493398 586102
rect 492970 585922 493026 585978
rect 493094 585922 493150 585978
rect 493218 585922 493274 585978
rect 493342 585922 493398 585978
rect 492970 568294 493026 568350
rect 493094 568294 493150 568350
rect 493218 568294 493274 568350
rect 493342 568294 493398 568350
rect 492970 568170 493026 568226
rect 493094 568170 493150 568226
rect 493218 568170 493274 568226
rect 493342 568170 493398 568226
rect 492970 568046 493026 568102
rect 493094 568046 493150 568102
rect 493218 568046 493274 568102
rect 493342 568046 493398 568102
rect 492970 567922 493026 567978
rect 493094 567922 493150 567978
rect 493218 567922 493274 567978
rect 493342 567922 493398 567978
rect 492970 550294 493026 550350
rect 493094 550294 493150 550350
rect 493218 550294 493274 550350
rect 493342 550294 493398 550350
rect 492970 550170 493026 550226
rect 493094 550170 493150 550226
rect 493218 550170 493274 550226
rect 493342 550170 493398 550226
rect 492970 550046 493026 550102
rect 493094 550046 493150 550102
rect 493218 550046 493274 550102
rect 493342 550046 493398 550102
rect 492970 549922 493026 549978
rect 493094 549922 493150 549978
rect 493218 549922 493274 549978
rect 493342 549922 493398 549978
rect 492970 532294 493026 532350
rect 493094 532294 493150 532350
rect 493218 532294 493274 532350
rect 493342 532294 493398 532350
rect 492970 532170 493026 532226
rect 493094 532170 493150 532226
rect 493218 532170 493274 532226
rect 493342 532170 493398 532226
rect 492970 532046 493026 532102
rect 493094 532046 493150 532102
rect 493218 532046 493274 532102
rect 493342 532046 493398 532102
rect 492970 531922 493026 531978
rect 493094 531922 493150 531978
rect 493218 531922 493274 531978
rect 493342 531922 493398 531978
rect 492970 514294 493026 514350
rect 493094 514294 493150 514350
rect 493218 514294 493274 514350
rect 493342 514294 493398 514350
rect 492970 514170 493026 514226
rect 493094 514170 493150 514226
rect 493218 514170 493274 514226
rect 493342 514170 493398 514226
rect 492970 514046 493026 514102
rect 493094 514046 493150 514102
rect 493218 514046 493274 514102
rect 493342 514046 493398 514102
rect 492970 513922 493026 513978
rect 493094 513922 493150 513978
rect 493218 513922 493274 513978
rect 493342 513922 493398 513978
rect 492970 496294 493026 496350
rect 493094 496294 493150 496350
rect 493218 496294 493274 496350
rect 493342 496294 493398 496350
rect 492970 496170 493026 496226
rect 493094 496170 493150 496226
rect 493218 496170 493274 496226
rect 493342 496170 493398 496226
rect 492970 496046 493026 496102
rect 493094 496046 493150 496102
rect 493218 496046 493274 496102
rect 493342 496046 493398 496102
rect 492970 495922 493026 495978
rect 493094 495922 493150 495978
rect 493218 495922 493274 495978
rect 493342 495922 493398 495978
rect 492970 478294 493026 478350
rect 493094 478294 493150 478350
rect 493218 478294 493274 478350
rect 493342 478294 493398 478350
rect 492970 478170 493026 478226
rect 493094 478170 493150 478226
rect 493218 478170 493274 478226
rect 493342 478170 493398 478226
rect 492970 478046 493026 478102
rect 493094 478046 493150 478102
rect 493218 478046 493274 478102
rect 493342 478046 493398 478102
rect 492970 477922 493026 477978
rect 493094 477922 493150 477978
rect 493218 477922 493274 477978
rect 493342 477922 493398 477978
rect 492970 460294 493026 460350
rect 493094 460294 493150 460350
rect 493218 460294 493274 460350
rect 493342 460294 493398 460350
rect 492970 460170 493026 460226
rect 493094 460170 493150 460226
rect 493218 460170 493274 460226
rect 493342 460170 493398 460226
rect 492970 460046 493026 460102
rect 493094 460046 493150 460102
rect 493218 460046 493274 460102
rect 493342 460046 493398 460102
rect 492970 459922 493026 459978
rect 493094 459922 493150 459978
rect 493218 459922 493274 459978
rect 493342 459922 493398 459978
rect 492970 442294 493026 442350
rect 493094 442294 493150 442350
rect 493218 442294 493274 442350
rect 493342 442294 493398 442350
rect 492970 442170 493026 442226
rect 493094 442170 493150 442226
rect 493218 442170 493274 442226
rect 493342 442170 493398 442226
rect 492970 442046 493026 442102
rect 493094 442046 493150 442102
rect 493218 442046 493274 442102
rect 493342 442046 493398 442102
rect 492970 441922 493026 441978
rect 493094 441922 493150 441978
rect 493218 441922 493274 441978
rect 493342 441922 493398 441978
rect 492970 424294 493026 424350
rect 493094 424294 493150 424350
rect 493218 424294 493274 424350
rect 493342 424294 493398 424350
rect 492970 424170 493026 424226
rect 493094 424170 493150 424226
rect 493218 424170 493274 424226
rect 493342 424170 493398 424226
rect 492970 424046 493026 424102
rect 493094 424046 493150 424102
rect 493218 424046 493274 424102
rect 493342 424046 493398 424102
rect 492970 423922 493026 423978
rect 493094 423922 493150 423978
rect 493218 423922 493274 423978
rect 493342 423922 493398 423978
rect 492970 406294 493026 406350
rect 493094 406294 493150 406350
rect 493218 406294 493274 406350
rect 493342 406294 493398 406350
rect 492970 406170 493026 406226
rect 493094 406170 493150 406226
rect 493218 406170 493274 406226
rect 493342 406170 493398 406226
rect 492970 406046 493026 406102
rect 493094 406046 493150 406102
rect 493218 406046 493274 406102
rect 493342 406046 493398 406102
rect 492970 405922 493026 405978
rect 493094 405922 493150 405978
rect 493218 405922 493274 405978
rect 493342 405922 493398 405978
rect 492970 388294 493026 388350
rect 493094 388294 493150 388350
rect 493218 388294 493274 388350
rect 493342 388294 493398 388350
rect 492970 388170 493026 388226
rect 493094 388170 493150 388226
rect 493218 388170 493274 388226
rect 493342 388170 493398 388226
rect 492970 388046 493026 388102
rect 493094 388046 493150 388102
rect 493218 388046 493274 388102
rect 493342 388046 493398 388102
rect 492970 387922 493026 387978
rect 493094 387922 493150 387978
rect 493218 387922 493274 387978
rect 493342 387922 493398 387978
rect 492970 370294 493026 370350
rect 493094 370294 493150 370350
rect 493218 370294 493274 370350
rect 493342 370294 493398 370350
rect 492970 370170 493026 370226
rect 493094 370170 493150 370226
rect 493218 370170 493274 370226
rect 493342 370170 493398 370226
rect 492970 370046 493026 370102
rect 493094 370046 493150 370102
rect 493218 370046 493274 370102
rect 493342 370046 493398 370102
rect 492970 369922 493026 369978
rect 493094 369922 493150 369978
rect 493218 369922 493274 369978
rect 493342 369922 493398 369978
rect 492970 352294 493026 352350
rect 493094 352294 493150 352350
rect 493218 352294 493274 352350
rect 493342 352294 493398 352350
rect 492970 352170 493026 352226
rect 493094 352170 493150 352226
rect 493218 352170 493274 352226
rect 493342 352170 493398 352226
rect 492970 352046 493026 352102
rect 493094 352046 493150 352102
rect 493218 352046 493274 352102
rect 493342 352046 493398 352102
rect 492970 351922 493026 351978
rect 493094 351922 493150 351978
rect 493218 351922 493274 351978
rect 493342 351922 493398 351978
rect 492970 334294 493026 334350
rect 493094 334294 493150 334350
rect 493218 334294 493274 334350
rect 493342 334294 493398 334350
rect 492970 334170 493026 334226
rect 493094 334170 493150 334226
rect 493218 334170 493274 334226
rect 493342 334170 493398 334226
rect 492970 334046 493026 334102
rect 493094 334046 493150 334102
rect 493218 334046 493274 334102
rect 493342 334046 493398 334102
rect 492970 333922 493026 333978
rect 493094 333922 493150 333978
rect 493218 333922 493274 333978
rect 493342 333922 493398 333978
rect 492970 316294 493026 316350
rect 493094 316294 493150 316350
rect 493218 316294 493274 316350
rect 493342 316294 493398 316350
rect 492970 316170 493026 316226
rect 493094 316170 493150 316226
rect 493218 316170 493274 316226
rect 493342 316170 493398 316226
rect 492970 316046 493026 316102
rect 493094 316046 493150 316102
rect 493218 316046 493274 316102
rect 493342 316046 493398 316102
rect 492970 315922 493026 315978
rect 493094 315922 493150 315978
rect 493218 315922 493274 315978
rect 493342 315922 493398 315978
rect 492970 298294 493026 298350
rect 493094 298294 493150 298350
rect 493218 298294 493274 298350
rect 493342 298294 493398 298350
rect 492970 298170 493026 298226
rect 493094 298170 493150 298226
rect 493218 298170 493274 298226
rect 493342 298170 493398 298226
rect 492970 298046 493026 298102
rect 493094 298046 493150 298102
rect 493218 298046 493274 298102
rect 493342 298046 493398 298102
rect 492970 297922 493026 297978
rect 493094 297922 493150 297978
rect 493218 297922 493274 297978
rect 493342 297922 493398 297978
rect 492970 280294 493026 280350
rect 493094 280294 493150 280350
rect 493218 280294 493274 280350
rect 493342 280294 493398 280350
rect 492970 280170 493026 280226
rect 493094 280170 493150 280226
rect 493218 280170 493274 280226
rect 493342 280170 493398 280226
rect 492970 280046 493026 280102
rect 493094 280046 493150 280102
rect 493218 280046 493274 280102
rect 493342 280046 493398 280102
rect 492970 279922 493026 279978
rect 493094 279922 493150 279978
rect 493218 279922 493274 279978
rect 493342 279922 493398 279978
rect 492970 262294 493026 262350
rect 493094 262294 493150 262350
rect 493218 262294 493274 262350
rect 493342 262294 493398 262350
rect 492970 262170 493026 262226
rect 493094 262170 493150 262226
rect 493218 262170 493274 262226
rect 493342 262170 493398 262226
rect 492970 262046 493026 262102
rect 493094 262046 493150 262102
rect 493218 262046 493274 262102
rect 493342 262046 493398 262102
rect 492970 261922 493026 261978
rect 493094 261922 493150 261978
rect 493218 261922 493274 261978
rect 493342 261922 493398 261978
rect 492970 244294 493026 244350
rect 493094 244294 493150 244350
rect 493218 244294 493274 244350
rect 493342 244294 493398 244350
rect 492970 244170 493026 244226
rect 493094 244170 493150 244226
rect 493218 244170 493274 244226
rect 493342 244170 493398 244226
rect 492970 244046 493026 244102
rect 493094 244046 493150 244102
rect 493218 244046 493274 244102
rect 493342 244046 493398 244102
rect 492970 243922 493026 243978
rect 493094 243922 493150 243978
rect 493218 243922 493274 243978
rect 493342 243922 493398 243978
rect 492970 226294 493026 226350
rect 493094 226294 493150 226350
rect 493218 226294 493274 226350
rect 493342 226294 493398 226350
rect 492970 226170 493026 226226
rect 493094 226170 493150 226226
rect 493218 226170 493274 226226
rect 493342 226170 493398 226226
rect 492970 226046 493026 226102
rect 493094 226046 493150 226102
rect 493218 226046 493274 226102
rect 493342 226046 493398 226102
rect 492970 225922 493026 225978
rect 493094 225922 493150 225978
rect 493218 225922 493274 225978
rect 493342 225922 493398 225978
rect 507250 597156 507306 597212
rect 507374 597156 507430 597212
rect 507498 597156 507554 597212
rect 507622 597156 507678 597212
rect 507250 597032 507306 597088
rect 507374 597032 507430 597088
rect 507498 597032 507554 597088
rect 507622 597032 507678 597088
rect 507250 596908 507306 596964
rect 507374 596908 507430 596964
rect 507498 596908 507554 596964
rect 507622 596908 507678 596964
rect 507250 596784 507306 596840
rect 507374 596784 507430 596840
rect 507498 596784 507554 596840
rect 507622 596784 507678 596840
rect 507250 580294 507306 580350
rect 507374 580294 507430 580350
rect 507498 580294 507554 580350
rect 507622 580294 507678 580350
rect 507250 580170 507306 580226
rect 507374 580170 507430 580226
rect 507498 580170 507554 580226
rect 507622 580170 507678 580226
rect 507250 580046 507306 580102
rect 507374 580046 507430 580102
rect 507498 580046 507554 580102
rect 507622 580046 507678 580102
rect 507250 579922 507306 579978
rect 507374 579922 507430 579978
rect 507498 579922 507554 579978
rect 507622 579922 507678 579978
rect 507250 562294 507306 562350
rect 507374 562294 507430 562350
rect 507498 562294 507554 562350
rect 507622 562294 507678 562350
rect 507250 562170 507306 562226
rect 507374 562170 507430 562226
rect 507498 562170 507554 562226
rect 507622 562170 507678 562226
rect 507250 562046 507306 562102
rect 507374 562046 507430 562102
rect 507498 562046 507554 562102
rect 507622 562046 507678 562102
rect 507250 561922 507306 561978
rect 507374 561922 507430 561978
rect 507498 561922 507554 561978
rect 507622 561922 507678 561978
rect 507250 544294 507306 544350
rect 507374 544294 507430 544350
rect 507498 544294 507554 544350
rect 507622 544294 507678 544350
rect 507250 544170 507306 544226
rect 507374 544170 507430 544226
rect 507498 544170 507554 544226
rect 507622 544170 507678 544226
rect 507250 544046 507306 544102
rect 507374 544046 507430 544102
rect 507498 544046 507554 544102
rect 507622 544046 507678 544102
rect 507250 543922 507306 543978
rect 507374 543922 507430 543978
rect 507498 543922 507554 543978
rect 507622 543922 507678 543978
rect 507250 526294 507306 526350
rect 507374 526294 507430 526350
rect 507498 526294 507554 526350
rect 507622 526294 507678 526350
rect 507250 526170 507306 526226
rect 507374 526170 507430 526226
rect 507498 526170 507554 526226
rect 507622 526170 507678 526226
rect 507250 526046 507306 526102
rect 507374 526046 507430 526102
rect 507498 526046 507554 526102
rect 507622 526046 507678 526102
rect 507250 525922 507306 525978
rect 507374 525922 507430 525978
rect 507498 525922 507554 525978
rect 507622 525922 507678 525978
rect 507250 508294 507306 508350
rect 507374 508294 507430 508350
rect 507498 508294 507554 508350
rect 507622 508294 507678 508350
rect 507250 508170 507306 508226
rect 507374 508170 507430 508226
rect 507498 508170 507554 508226
rect 507622 508170 507678 508226
rect 507250 508046 507306 508102
rect 507374 508046 507430 508102
rect 507498 508046 507554 508102
rect 507622 508046 507678 508102
rect 507250 507922 507306 507978
rect 507374 507922 507430 507978
rect 507498 507922 507554 507978
rect 507622 507922 507678 507978
rect 507250 490294 507306 490350
rect 507374 490294 507430 490350
rect 507498 490294 507554 490350
rect 507622 490294 507678 490350
rect 507250 490170 507306 490226
rect 507374 490170 507430 490226
rect 507498 490170 507554 490226
rect 507622 490170 507678 490226
rect 507250 490046 507306 490102
rect 507374 490046 507430 490102
rect 507498 490046 507554 490102
rect 507622 490046 507678 490102
rect 507250 489922 507306 489978
rect 507374 489922 507430 489978
rect 507498 489922 507554 489978
rect 507622 489922 507678 489978
rect 507250 472294 507306 472350
rect 507374 472294 507430 472350
rect 507498 472294 507554 472350
rect 507622 472294 507678 472350
rect 507250 472170 507306 472226
rect 507374 472170 507430 472226
rect 507498 472170 507554 472226
rect 507622 472170 507678 472226
rect 507250 472046 507306 472102
rect 507374 472046 507430 472102
rect 507498 472046 507554 472102
rect 507622 472046 507678 472102
rect 507250 471922 507306 471978
rect 507374 471922 507430 471978
rect 507498 471922 507554 471978
rect 507622 471922 507678 471978
rect 507250 454294 507306 454350
rect 507374 454294 507430 454350
rect 507498 454294 507554 454350
rect 507622 454294 507678 454350
rect 507250 454170 507306 454226
rect 507374 454170 507430 454226
rect 507498 454170 507554 454226
rect 507622 454170 507678 454226
rect 507250 454046 507306 454102
rect 507374 454046 507430 454102
rect 507498 454046 507554 454102
rect 507622 454046 507678 454102
rect 507250 453922 507306 453978
rect 507374 453922 507430 453978
rect 507498 453922 507554 453978
rect 507622 453922 507678 453978
rect 507250 436294 507306 436350
rect 507374 436294 507430 436350
rect 507498 436294 507554 436350
rect 507622 436294 507678 436350
rect 507250 436170 507306 436226
rect 507374 436170 507430 436226
rect 507498 436170 507554 436226
rect 507622 436170 507678 436226
rect 507250 436046 507306 436102
rect 507374 436046 507430 436102
rect 507498 436046 507554 436102
rect 507622 436046 507678 436102
rect 507250 435922 507306 435978
rect 507374 435922 507430 435978
rect 507498 435922 507554 435978
rect 507622 435922 507678 435978
rect 507250 418294 507306 418350
rect 507374 418294 507430 418350
rect 507498 418294 507554 418350
rect 507622 418294 507678 418350
rect 507250 418170 507306 418226
rect 507374 418170 507430 418226
rect 507498 418170 507554 418226
rect 507622 418170 507678 418226
rect 507250 418046 507306 418102
rect 507374 418046 507430 418102
rect 507498 418046 507554 418102
rect 507622 418046 507678 418102
rect 507250 417922 507306 417978
rect 507374 417922 507430 417978
rect 507498 417922 507554 417978
rect 507622 417922 507678 417978
rect 507250 400294 507306 400350
rect 507374 400294 507430 400350
rect 507498 400294 507554 400350
rect 507622 400294 507678 400350
rect 507250 400170 507306 400226
rect 507374 400170 507430 400226
rect 507498 400170 507554 400226
rect 507622 400170 507678 400226
rect 507250 400046 507306 400102
rect 507374 400046 507430 400102
rect 507498 400046 507554 400102
rect 507622 400046 507678 400102
rect 507250 399922 507306 399978
rect 507374 399922 507430 399978
rect 507498 399922 507554 399978
rect 507622 399922 507678 399978
rect 507250 382294 507306 382350
rect 507374 382294 507430 382350
rect 507498 382294 507554 382350
rect 507622 382294 507678 382350
rect 507250 382170 507306 382226
rect 507374 382170 507430 382226
rect 507498 382170 507554 382226
rect 507622 382170 507678 382226
rect 507250 382046 507306 382102
rect 507374 382046 507430 382102
rect 507498 382046 507554 382102
rect 507622 382046 507678 382102
rect 507250 381922 507306 381978
rect 507374 381922 507430 381978
rect 507498 381922 507554 381978
rect 507622 381922 507678 381978
rect 507250 364294 507306 364350
rect 507374 364294 507430 364350
rect 507498 364294 507554 364350
rect 507622 364294 507678 364350
rect 507250 364170 507306 364226
rect 507374 364170 507430 364226
rect 507498 364170 507554 364226
rect 507622 364170 507678 364226
rect 507250 364046 507306 364102
rect 507374 364046 507430 364102
rect 507498 364046 507554 364102
rect 507622 364046 507678 364102
rect 507250 363922 507306 363978
rect 507374 363922 507430 363978
rect 507498 363922 507554 363978
rect 507622 363922 507678 363978
rect 507250 346294 507306 346350
rect 507374 346294 507430 346350
rect 507498 346294 507554 346350
rect 507622 346294 507678 346350
rect 507250 346170 507306 346226
rect 507374 346170 507430 346226
rect 507498 346170 507554 346226
rect 507622 346170 507678 346226
rect 507250 346046 507306 346102
rect 507374 346046 507430 346102
rect 507498 346046 507554 346102
rect 507622 346046 507678 346102
rect 507250 345922 507306 345978
rect 507374 345922 507430 345978
rect 507498 345922 507554 345978
rect 507622 345922 507678 345978
rect 507250 328294 507306 328350
rect 507374 328294 507430 328350
rect 507498 328294 507554 328350
rect 507622 328294 507678 328350
rect 507250 328170 507306 328226
rect 507374 328170 507430 328226
rect 507498 328170 507554 328226
rect 507622 328170 507678 328226
rect 507250 328046 507306 328102
rect 507374 328046 507430 328102
rect 507498 328046 507554 328102
rect 507622 328046 507678 328102
rect 507250 327922 507306 327978
rect 507374 327922 507430 327978
rect 507498 327922 507554 327978
rect 507622 327922 507678 327978
rect 507250 310294 507306 310350
rect 507374 310294 507430 310350
rect 507498 310294 507554 310350
rect 507622 310294 507678 310350
rect 507250 310170 507306 310226
rect 507374 310170 507430 310226
rect 507498 310170 507554 310226
rect 507622 310170 507678 310226
rect 507250 310046 507306 310102
rect 507374 310046 507430 310102
rect 507498 310046 507554 310102
rect 507622 310046 507678 310102
rect 507250 309922 507306 309978
rect 507374 309922 507430 309978
rect 507498 309922 507554 309978
rect 507622 309922 507678 309978
rect 507250 292294 507306 292350
rect 507374 292294 507430 292350
rect 507498 292294 507554 292350
rect 507622 292294 507678 292350
rect 507250 292170 507306 292226
rect 507374 292170 507430 292226
rect 507498 292170 507554 292226
rect 507622 292170 507678 292226
rect 507250 292046 507306 292102
rect 507374 292046 507430 292102
rect 507498 292046 507554 292102
rect 507622 292046 507678 292102
rect 507250 291922 507306 291978
rect 507374 291922 507430 291978
rect 507498 291922 507554 291978
rect 507622 291922 507678 291978
rect 507250 274294 507306 274350
rect 507374 274294 507430 274350
rect 507498 274294 507554 274350
rect 507622 274294 507678 274350
rect 507250 274170 507306 274226
rect 507374 274170 507430 274226
rect 507498 274170 507554 274226
rect 507622 274170 507678 274226
rect 507250 274046 507306 274102
rect 507374 274046 507430 274102
rect 507498 274046 507554 274102
rect 507622 274046 507678 274102
rect 507250 273922 507306 273978
rect 507374 273922 507430 273978
rect 507498 273922 507554 273978
rect 507622 273922 507678 273978
rect 507250 256294 507306 256350
rect 507374 256294 507430 256350
rect 507498 256294 507554 256350
rect 507622 256294 507678 256350
rect 507250 256170 507306 256226
rect 507374 256170 507430 256226
rect 507498 256170 507554 256226
rect 507622 256170 507678 256226
rect 507250 256046 507306 256102
rect 507374 256046 507430 256102
rect 507498 256046 507554 256102
rect 507622 256046 507678 256102
rect 507250 255922 507306 255978
rect 507374 255922 507430 255978
rect 507498 255922 507554 255978
rect 507622 255922 507678 255978
rect 507250 238294 507306 238350
rect 507374 238294 507430 238350
rect 507498 238294 507554 238350
rect 507622 238294 507678 238350
rect 507250 238170 507306 238226
rect 507374 238170 507430 238226
rect 507498 238170 507554 238226
rect 507622 238170 507678 238226
rect 507250 238046 507306 238102
rect 507374 238046 507430 238102
rect 507498 238046 507554 238102
rect 507622 238046 507678 238102
rect 507250 237922 507306 237978
rect 507374 237922 507430 237978
rect 507498 237922 507554 237978
rect 507622 237922 507678 237978
rect 507250 220294 507306 220350
rect 507374 220294 507430 220350
rect 507498 220294 507554 220350
rect 507622 220294 507678 220350
rect 507250 220170 507306 220226
rect 507374 220170 507430 220226
rect 507498 220170 507554 220226
rect 507622 220170 507678 220226
rect 507250 220046 507306 220102
rect 507374 220046 507430 220102
rect 507498 220046 507554 220102
rect 507622 220046 507678 220102
rect 507250 219922 507306 219978
rect 507374 219922 507430 219978
rect 507498 219922 507554 219978
rect 507622 219922 507678 219978
rect 510970 598116 511026 598172
rect 511094 598116 511150 598172
rect 511218 598116 511274 598172
rect 511342 598116 511398 598172
rect 510970 597992 511026 598048
rect 511094 597992 511150 598048
rect 511218 597992 511274 598048
rect 511342 597992 511398 598048
rect 510970 597868 511026 597924
rect 511094 597868 511150 597924
rect 511218 597868 511274 597924
rect 511342 597868 511398 597924
rect 510970 597744 511026 597800
rect 511094 597744 511150 597800
rect 511218 597744 511274 597800
rect 511342 597744 511398 597800
rect 510970 586294 511026 586350
rect 511094 586294 511150 586350
rect 511218 586294 511274 586350
rect 511342 586294 511398 586350
rect 510970 586170 511026 586226
rect 511094 586170 511150 586226
rect 511218 586170 511274 586226
rect 511342 586170 511398 586226
rect 510970 586046 511026 586102
rect 511094 586046 511150 586102
rect 511218 586046 511274 586102
rect 511342 586046 511398 586102
rect 510970 585922 511026 585978
rect 511094 585922 511150 585978
rect 511218 585922 511274 585978
rect 511342 585922 511398 585978
rect 510970 568294 511026 568350
rect 511094 568294 511150 568350
rect 511218 568294 511274 568350
rect 511342 568294 511398 568350
rect 510970 568170 511026 568226
rect 511094 568170 511150 568226
rect 511218 568170 511274 568226
rect 511342 568170 511398 568226
rect 510970 568046 511026 568102
rect 511094 568046 511150 568102
rect 511218 568046 511274 568102
rect 511342 568046 511398 568102
rect 510970 567922 511026 567978
rect 511094 567922 511150 567978
rect 511218 567922 511274 567978
rect 511342 567922 511398 567978
rect 510970 550294 511026 550350
rect 511094 550294 511150 550350
rect 511218 550294 511274 550350
rect 511342 550294 511398 550350
rect 510970 550170 511026 550226
rect 511094 550170 511150 550226
rect 511218 550170 511274 550226
rect 511342 550170 511398 550226
rect 510970 550046 511026 550102
rect 511094 550046 511150 550102
rect 511218 550046 511274 550102
rect 511342 550046 511398 550102
rect 510970 549922 511026 549978
rect 511094 549922 511150 549978
rect 511218 549922 511274 549978
rect 511342 549922 511398 549978
rect 510970 532294 511026 532350
rect 511094 532294 511150 532350
rect 511218 532294 511274 532350
rect 511342 532294 511398 532350
rect 510970 532170 511026 532226
rect 511094 532170 511150 532226
rect 511218 532170 511274 532226
rect 511342 532170 511398 532226
rect 510970 532046 511026 532102
rect 511094 532046 511150 532102
rect 511218 532046 511274 532102
rect 511342 532046 511398 532102
rect 510970 531922 511026 531978
rect 511094 531922 511150 531978
rect 511218 531922 511274 531978
rect 511342 531922 511398 531978
rect 510970 514294 511026 514350
rect 511094 514294 511150 514350
rect 511218 514294 511274 514350
rect 511342 514294 511398 514350
rect 510970 514170 511026 514226
rect 511094 514170 511150 514226
rect 511218 514170 511274 514226
rect 511342 514170 511398 514226
rect 510970 514046 511026 514102
rect 511094 514046 511150 514102
rect 511218 514046 511274 514102
rect 511342 514046 511398 514102
rect 510970 513922 511026 513978
rect 511094 513922 511150 513978
rect 511218 513922 511274 513978
rect 511342 513922 511398 513978
rect 510970 496294 511026 496350
rect 511094 496294 511150 496350
rect 511218 496294 511274 496350
rect 511342 496294 511398 496350
rect 510970 496170 511026 496226
rect 511094 496170 511150 496226
rect 511218 496170 511274 496226
rect 511342 496170 511398 496226
rect 510970 496046 511026 496102
rect 511094 496046 511150 496102
rect 511218 496046 511274 496102
rect 511342 496046 511398 496102
rect 510970 495922 511026 495978
rect 511094 495922 511150 495978
rect 511218 495922 511274 495978
rect 511342 495922 511398 495978
rect 510970 478294 511026 478350
rect 511094 478294 511150 478350
rect 511218 478294 511274 478350
rect 511342 478294 511398 478350
rect 510970 478170 511026 478226
rect 511094 478170 511150 478226
rect 511218 478170 511274 478226
rect 511342 478170 511398 478226
rect 510970 478046 511026 478102
rect 511094 478046 511150 478102
rect 511218 478046 511274 478102
rect 511342 478046 511398 478102
rect 510970 477922 511026 477978
rect 511094 477922 511150 477978
rect 511218 477922 511274 477978
rect 511342 477922 511398 477978
rect 510970 460294 511026 460350
rect 511094 460294 511150 460350
rect 511218 460294 511274 460350
rect 511342 460294 511398 460350
rect 510970 460170 511026 460226
rect 511094 460170 511150 460226
rect 511218 460170 511274 460226
rect 511342 460170 511398 460226
rect 510970 460046 511026 460102
rect 511094 460046 511150 460102
rect 511218 460046 511274 460102
rect 511342 460046 511398 460102
rect 510970 459922 511026 459978
rect 511094 459922 511150 459978
rect 511218 459922 511274 459978
rect 511342 459922 511398 459978
rect 510970 442294 511026 442350
rect 511094 442294 511150 442350
rect 511218 442294 511274 442350
rect 511342 442294 511398 442350
rect 510970 442170 511026 442226
rect 511094 442170 511150 442226
rect 511218 442170 511274 442226
rect 511342 442170 511398 442226
rect 510970 442046 511026 442102
rect 511094 442046 511150 442102
rect 511218 442046 511274 442102
rect 511342 442046 511398 442102
rect 510970 441922 511026 441978
rect 511094 441922 511150 441978
rect 511218 441922 511274 441978
rect 511342 441922 511398 441978
rect 510970 424294 511026 424350
rect 511094 424294 511150 424350
rect 511218 424294 511274 424350
rect 511342 424294 511398 424350
rect 510970 424170 511026 424226
rect 511094 424170 511150 424226
rect 511218 424170 511274 424226
rect 511342 424170 511398 424226
rect 510970 424046 511026 424102
rect 511094 424046 511150 424102
rect 511218 424046 511274 424102
rect 511342 424046 511398 424102
rect 510970 423922 511026 423978
rect 511094 423922 511150 423978
rect 511218 423922 511274 423978
rect 511342 423922 511398 423978
rect 510970 406294 511026 406350
rect 511094 406294 511150 406350
rect 511218 406294 511274 406350
rect 511342 406294 511398 406350
rect 510970 406170 511026 406226
rect 511094 406170 511150 406226
rect 511218 406170 511274 406226
rect 511342 406170 511398 406226
rect 510970 406046 511026 406102
rect 511094 406046 511150 406102
rect 511218 406046 511274 406102
rect 511342 406046 511398 406102
rect 510970 405922 511026 405978
rect 511094 405922 511150 405978
rect 511218 405922 511274 405978
rect 511342 405922 511398 405978
rect 510970 388294 511026 388350
rect 511094 388294 511150 388350
rect 511218 388294 511274 388350
rect 511342 388294 511398 388350
rect 510970 388170 511026 388226
rect 511094 388170 511150 388226
rect 511218 388170 511274 388226
rect 511342 388170 511398 388226
rect 510970 388046 511026 388102
rect 511094 388046 511150 388102
rect 511218 388046 511274 388102
rect 511342 388046 511398 388102
rect 510970 387922 511026 387978
rect 511094 387922 511150 387978
rect 511218 387922 511274 387978
rect 511342 387922 511398 387978
rect 510970 370294 511026 370350
rect 511094 370294 511150 370350
rect 511218 370294 511274 370350
rect 511342 370294 511398 370350
rect 510970 370170 511026 370226
rect 511094 370170 511150 370226
rect 511218 370170 511274 370226
rect 511342 370170 511398 370226
rect 510970 370046 511026 370102
rect 511094 370046 511150 370102
rect 511218 370046 511274 370102
rect 511342 370046 511398 370102
rect 510970 369922 511026 369978
rect 511094 369922 511150 369978
rect 511218 369922 511274 369978
rect 511342 369922 511398 369978
rect 510970 352294 511026 352350
rect 511094 352294 511150 352350
rect 511218 352294 511274 352350
rect 511342 352294 511398 352350
rect 510970 352170 511026 352226
rect 511094 352170 511150 352226
rect 511218 352170 511274 352226
rect 511342 352170 511398 352226
rect 510970 352046 511026 352102
rect 511094 352046 511150 352102
rect 511218 352046 511274 352102
rect 511342 352046 511398 352102
rect 510970 351922 511026 351978
rect 511094 351922 511150 351978
rect 511218 351922 511274 351978
rect 511342 351922 511398 351978
rect 510970 334294 511026 334350
rect 511094 334294 511150 334350
rect 511218 334294 511274 334350
rect 511342 334294 511398 334350
rect 510970 334170 511026 334226
rect 511094 334170 511150 334226
rect 511218 334170 511274 334226
rect 511342 334170 511398 334226
rect 510970 334046 511026 334102
rect 511094 334046 511150 334102
rect 511218 334046 511274 334102
rect 511342 334046 511398 334102
rect 510970 333922 511026 333978
rect 511094 333922 511150 333978
rect 511218 333922 511274 333978
rect 511342 333922 511398 333978
rect 510970 316294 511026 316350
rect 511094 316294 511150 316350
rect 511218 316294 511274 316350
rect 511342 316294 511398 316350
rect 510970 316170 511026 316226
rect 511094 316170 511150 316226
rect 511218 316170 511274 316226
rect 511342 316170 511398 316226
rect 510970 316046 511026 316102
rect 511094 316046 511150 316102
rect 511218 316046 511274 316102
rect 511342 316046 511398 316102
rect 510970 315922 511026 315978
rect 511094 315922 511150 315978
rect 511218 315922 511274 315978
rect 511342 315922 511398 315978
rect 510970 298294 511026 298350
rect 511094 298294 511150 298350
rect 511218 298294 511274 298350
rect 511342 298294 511398 298350
rect 510970 298170 511026 298226
rect 511094 298170 511150 298226
rect 511218 298170 511274 298226
rect 511342 298170 511398 298226
rect 510970 298046 511026 298102
rect 511094 298046 511150 298102
rect 511218 298046 511274 298102
rect 511342 298046 511398 298102
rect 510970 297922 511026 297978
rect 511094 297922 511150 297978
rect 511218 297922 511274 297978
rect 511342 297922 511398 297978
rect 510970 280294 511026 280350
rect 511094 280294 511150 280350
rect 511218 280294 511274 280350
rect 511342 280294 511398 280350
rect 510970 280170 511026 280226
rect 511094 280170 511150 280226
rect 511218 280170 511274 280226
rect 511342 280170 511398 280226
rect 510970 280046 511026 280102
rect 511094 280046 511150 280102
rect 511218 280046 511274 280102
rect 511342 280046 511398 280102
rect 510970 279922 511026 279978
rect 511094 279922 511150 279978
rect 511218 279922 511274 279978
rect 511342 279922 511398 279978
rect 510970 262294 511026 262350
rect 511094 262294 511150 262350
rect 511218 262294 511274 262350
rect 511342 262294 511398 262350
rect 510970 262170 511026 262226
rect 511094 262170 511150 262226
rect 511218 262170 511274 262226
rect 511342 262170 511398 262226
rect 510970 262046 511026 262102
rect 511094 262046 511150 262102
rect 511218 262046 511274 262102
rect 511342 262046 511398 262102
rect 510970 261922 511026 261978
rect 511094 261922 511150 261978
rect 511218 261922 511274 261978
rect 511342 261922 511398 261978
rect 510970 244294 511026 244350
rect 511094 244294 511150 244350
rect 511218 244294 511274 244350
rect 511342 244294 511398 244350
rect 510970 244170 511026 244226
rect 511094 244170 511150 244226
rect 511218 244170 511274 244226
rect 511342 244170 511398 244226
rect 510970 244046 511026 244102
rect 511094 244046 511150 244102
rect 511218 244046 511274 244102
rect 511342 244046 511398 244102
rect 510970 243922 511026 243978
rect 511094 243922 511150 243978
rect 511218 243922 511274 243978
rect 511342 243922 511398 243978
rect 528970 598116 529026 598172
rect 529094 598116 529150 598172
rect 529218 598116 529274 598172
rect 529342 598116 529398 598172
rect 528970 597992 529026 598048
rect 529094 597992 529150 598048
rect 529218 597992 529274 598048
rect 529342 597992 529398 598048
rect 528970 597868 529026 597924
rect 529094 597868 529150 597924
rect 529218 597868 529274 597924
rect 529342 597868 529398 597924
rect 528970 597744 529026 597800
rect 529094 597744 529150 597800
rect 529218 597744 529274 597800
rect 529342 597744 529398 597800
rect 543250 597156 543306 597212
rect 543374 597156 543430 597212
rect 543498 597156 543554 597212
rect 543622 597156 543678 597212
rect 543250 597032 543306 597088
rect 543374 597032 543430 597088
rect 543498 597032 543554 597088
rect 543622 597032 543678 597088
rect 543250 596908 543306 596964
rect 543374 596908 543430 596964
rect 543498 596908 543554 596964
rect 543622 596908 543678 596964
rect 543250 596784 543306 596840
rect 543374 596784 543430 596840
rect 543498 596784 543554 596840
rect 543622 596784 543678 596840
rect 528970 586294 529026 586350
rect 529094 586294 529150 586350
rect 529218 586294 529274 586350
rect 529342 586294 529398 586350
rect 528970 586170 529026 586226
rect 529094 586170 529150 586226
rect 529218 586170 529274 586226
rect 529342 586170 529398 586226
rect 528970 586046 529026 586102
rect 529094 586046 529150 586102
rect 529218 586046 529274 586102
rect 529342 586046 529398 586102
rect 528970 585922 529026 585978
rect 529094 585922 529150 585978
rect 529218 585922 529274 585978
rect 529342 585922 529398 585978
rect 528970 568294 529026 568350
rect 529094 568294 529150 568350
rect 529218 568294 529274 568350
rect 529342 568294 529398 568350
rect 528970 568170 529026 568226
rect 529094 568170 529150 568226
rect 529218 568170 529274 568226
rect 529342 568170 529398 568226
rect 528970 568046 529026 568102
rect 529094 568046 529150 568102
rect 529218 568046 529274 568102
rect 529342 568046 529398 568102
rect 528970 567922 529026 567978
rect 529094 567922 529150 567978
rect 529218 567922 529274 567978
rect 529342 567922 529398 567978
rect 528970 550294 529026 550350
rect 529094 550294 529150 550350
rect 529218 550294 529274 550350
rect 529342 550294 529398 550350
rect 528970 550170 529026 550226
rect 529094 550170 529150 550226
rect 529218 550170 529274 550226
rect 529342 550170 529398 550226
rect 528970 550046 529026 550102
rect 529094 550046 529150 550102
rect 529218 550046 529274 550102
rect 529342 550046 529398 550102
rect 528970 549922 529026 549978
rect 529094 549922 529150 549978
rect 529218 549922 529274 549978
rect 529342 549922 529398 549978
rect 528970 532294 529026 532350
rect 529094 532294 529150 532350
rect 529218 532294 529274 532350
rect 529342 532294 529398 532350
rect 528970 532170 529026 532226
rect 529094 532170 529150 532226
rect 529218 532170 529274 532226
rect 529342 532170 529398 532226
rect 528970 532046 529026 532102
rect 529094 532046 529150 532102
rect 529218 532046 529274 532102
rect 529342 532046 529398 532102
rect 528970 531922 529026 531978
rect 529094 531922 529150 531978
rect 529218 531922 529274 531978
rect 529342 531922 529398 531978
rect 528970 514294 529026 514350
rect 529094 514294 529150 514350
rect 529218 514294 529274 514350
rect 529342 514294 529398 514350
rect 528970 514170 529026 514226
rect 529094 514170 529150 514226
rect 529218 514170 529274 514226
rect 529342 514170 529398 514226
rect 528970 514046 529026 514102
rect 529094 514046 529150 514102
rect 529218 514046 529274 514102
rect 529342 514046 529398 514102
rect 528970 513922 529026 513978
rect 529094 513922 529150 513978
rect 529218 513922 529274 513978
rect 529342 513922 529398 513978
rect 528970 496294 529026 496350
rect 529094 496294 529150 496350
rect 529218 496294 529274 496350
rect 529342 496294 529398 496350
rect 528970 496170 529026 496226
rect 529094 496170 529150 496226
rect 529218 496170 529274 496226
rect 529342 496170 529398 496226
rect 528970 496046 529026 496102
rect 529094 496046 529150 496102
rect 529218 496046 529274 496102
rect 529342 496046 529398 496102
rect 528970 495922 529026 495978
rect 529094 495922 529150 495978
rect 529218 495922 529274 495978
rect 529342 495922 529398 495978
rect 528970 478294 529026 478350
rect 529094 478294 529150 478350
rect 529218 478294 529274 478350
rect 529342 478294 529398 478350
rect 528970 478170 529026 478226
rect 529094 478170 529150 478226
rect 529218 478170 529274 478226
rect 529342 478170 529398 478226
rect 528970 478046 529026 478102
rect 529094 478046 529150 478102
rect 529218 478046 529274 478102
rect 529342 478046 529398 478102
rect 528970 477922 529026 477978
rect 529094 477922 529150 477978
rect 529218 477922 529274 477978
rect 529342 477922 529398 477978
rect 528970 460294 529026 460350
rect 529094 460294 529150 460350
rect 529218 460294 529274 460350
rect 529342 460294 529398 460350
rect 528970 460170 529026 460226
rect 529094 460170 529150 460226
rect 529218 460170 529274 460226
rect 529342 460170 529398 460226
rect 528970 460046 529026 460102
rect 529094 460046 529150 460102
rect 529218 460046 529274 460102
rect 529342 460046 529398 460102
rect 528970 459922 529026 459978
rect 529094 459922 529150 459978
rect 529218 459922 529274 459978
rect 529342 459922 529398 459978
rect 528970 442294 529026 442350
rect 529094 442294 529150 442350
rect 529218 442294 529274 442350
rect 529342 442294 529398 442350
rect 528970 442170 529026 442226
rect 529094 442170 529150 442226
rect 529218 442170 529274 442226
rect 529342 442170 529398 442226
rect 528970 442046 529026 442102
rect 529094 442046 529150 442102
rect 529218 442046 529274 442102
rect 529342 442046 529398 442102
rect 528970 441922 529026 441978
rect 529094 441922 529150 441978
rect 529218 441922 529274 441978
rect 529342 441922 529398 441978
rect 528970 424294 529026 424350
rect 529094 424294 529150 424350
rect 529218 424294 529274 424350
rect 529342 424294 529398 424350
rect 528970 424170 529026 424226
rect 529094 424170 529150 424226
rect 529218 424170 529274 424226
rect 529342 424170 529398 424226
rect 528970 424046 529026 424102
rect 529094 424046 529150 424102
rect 529218 424046 529274 424102
rect 529342 424046 529398 424102
rect 528970 423922 529026 423978
rect 529094 423922 529150 423978
rect 529218 423922 529274 423978
rect 529342 423922 529398 423978
rect 528970 406294 529026 406350
rect 529094 406294 529150 406350
rect 529218 406294 529274 406350
rect 529342 406294 529398 406350
rect 528970 406170 529026 406226
rect 529094 406170 529150 406226
rect 529218 406170 529274 406226
rect 529342 406170 529398 406226
rect 528970 406046 529026 406102
rect 529094 406046 529150 406102
rect 529218 406046 529274 406102
rect 529342 406046 529398 406102
rect 528970 405922 529026 405978
rect 529094 405922 529150 405978
rect 529218 405922 529274 405978
rect 529342 405922 529398 405978
rect 528970 388294 529026 388350
rect 529094 388294 529150 388350
rect 529218 388294 529274 388350
rect 529342 388294 529398 388350
rect 528970 388170 529026 388226
rect 529094 388170 529150 388226
rect 529218 388170 529274 388226
rect 529342 388170 529398 388226
rect 528970 388046 529026 388102
rect 529094 388046 529150 388102
rect 529218 388046 529274 388102
rect 529342 388046 529398 388102
rect 528970 387922 529026 387978
rect 529094 387922 529150 387978
rect 529218 387922 529274 387978
rect 529342 387922 529398 387978
rect 528970 370294 529026 370350
rect 529094 370294 529150 370350
rect 529218 370294 529274 370350
rect 529342 370294 529398 370350
rect 528970 370170 529026 370226
rect 529094 370170 529150 370226
rect 529218 370170 529274 370226
rect 529342 370170 529398 370226
rect 528970 370046 529026 370102
rect 529094 370046 529150 370102
rect 529218 370046 529274 370102
rect 529342 370046 529398 370102
rect 528970 369922 529026 369978
rect 529094 369922 529150 369978
rect 529218 369922 529274 369978
rect 529342 369922 529398 369978
rect 528970 352294 529026 352350
rect 529094 352294 529150 352350
rect 529218 352294 529274 352350
rect 529342 352294 529398 352350
rect 528970 352170 529026 352226
rect 529094 352170 529150 352226
rect 529218 352170 529274 352226
rect 529342 352170 529398 352226
rect 528970 352046 529026 352102
rect 529094 352046 529150 352102
rect 529218 352046 529274 352102
rect 529342 352046 529398 352102
rect 528970 351922 529026 351978
rect 529094 351922 529150 351978
rect 529218 351922 529274 351978
rect 529342 351922 529398 351978
rect 528970 334294 529026 334350
rect 529094 334294 529150 334350
rect 529218 334294 529274 334350
rect 529342 334294 529398 334350
rect 528970 334170 529026 334226
rect 529094 334170 529150 334226
rect 529218 334170 529274 334226
rect 529342 334170 529398 334226
rect 528970 334046 529026 334102
rect 529094 334046 529150 334102
rect 529218 334046 529274 334102
rect 529342 334046 529398 334102
rect 528970 333922 529026 333978
rect 529094 333922 529150 333978
rect 529218 333922 529274 333978
rect 529342 333922 529398 333978
rect 528970 316294 529026 316350
rect 529094 316294 529150 316350
rect 529218 316294 529274 316350
rect 529342 316294 529398 316350
rect 528970 316170 529026 316226
rect 529094 316170 529150 316226
rect 529218 316170 529274 316226
rect 529342 316170 529398 316226
rect 528970 316046 529026 316102
rect 529094 316046 529150 316102
rect 529218 316046 529274 316102
rect 529342 316046 529398 316102
rect 528970 315922 529026 315978
rect 529094 315922 529150 315978
rect 529218 315922 529274 315978
rect 529342 315922 529398 315978
rect 528970 298294 529026 298350
rect 529094 298294 529150 298350
rect 529218 298294 529274 298350
rect 529342 298294 529398 298350
rect 528970 298170 529026 298226
rect 529094 298170 529150 298226
rect 529218 298170 529274 298226
rect 529342 298170 529398 298226
rect 528970 298046 529026 298102
rect 529094 298046 529150 298102
rect 529218 298046 529274 298102
rect 529342 298046 529398 298102
rect 528970 297922 529026 297978
rect 529094 297922 529150 297978
rect 529218 297922 529274 297978
rect 529342 297922 529398 297978
rect 528970 280294 529026 280350
rect 529094 280294 529150 280350
rect 529218 280294 529274 280350
rect 529342 280294 529398 280350
rect 528970 280170 529026 280226
rect 529094 280170 529150 280226
rect 529218 280170 529274 280226
rect 529342 280170 529398 280226
rect 528970 280046 529026 280102
rect 529094 280046 529150 280102
rect 529218 280046 529274 280102
rect 529342 280046 529398 280102
rect 528970 279922 529026 279978
rect 529094 279922 529150 279978
rect 529218 279922 529274 279978
rect 529342 279922 529398 279978
rect 528970 262294 529026 262350
rect 529094 262294 529150 262350
rect 529218 262294 529274 262350
rect 529342 262294 529398 262350
rect 528970 262170 529026 262226
rect 529094 262170 529150 262226
rect 529218 262170 529274 262226
rect 529342 262170 529398 262226
rect 528970 262046 529026 262102
rect 529094 262046 529150 262102
rect 529218 262046 529274 262102
rect 529342 262046 529398 262102
rect 528970 261922 529026 261978
rect 529094 261922 529150 261978
rect 529218 261922 529274 261978
rect 529342 261922 529398 261978
rect 528970 244294 529026 244350
rect 529094 244294 529150 244350
rect 529218 244294 529274 244350
rect 529342 244294 529398 244350
rect 528970 244170 529026 244226
rect 529094 244170 529150 244226
rect 529218 244170 529274 244226
rect 529342 244170 529398 244226
rect 528970 244046 529026 244102
rect 529094 244046 529150 244102
rect 529218 244046 529274 244102
rect 529342 244046 529398 244102
rect 528970 243922 529026 243978
rect 529094 243922 529150 243978
rect 529218 243922 529274 243978
rect 529342 243922 529398 243978
rect 510970 226294 511026 226350
rect 511094 226294 511150 226350
rect 511218 226294 511274 226350
rect 511342 226294 511398 226350
rect 510970 226170 511026 226226
rect 511094 226170 511150 226226
rect 511218 226170 511274 226226
rect 511342 226170 511398 226226
rect 510970 226046 511026 226102
rect 511094 226046 511150 226102
rect 511218 226046 511274 226102
rect 511342 226046 511398 226102
rect 510970 225922 511026 225978
rect 511094 225922 511150 225978
rect 511218 225922 511274 225978
rect 511342 225922 511398 225978
rect 525250 238294 525306 238350
rect 525374 238294 525430 238350
rect 525498 238294 525554 238350
rect 525622 238294 525678 238350
rect 525250 238170 525306 238226
rect 525374 238170 525430 238226
rect 525498 238170 525554 238226
rect 525622 238170 525678 238226
rect 525250 238046 525306 238102
rect 525374 238046 525430 238102
rect 525498 238046 525554 238102
rect 525622 238046 525678 238102
rect 525250 237922 525306 237978
rect 525374 237922 525430 237978
rect 525498 237922 525554 237978
rect 525622 237922 525678 237978
rect 525250 220294 525306 220350
rect 525374 220294 525430 220350
rect 525498 220294 525554 220350
rect 525622 220294 525678 220350
rect 525250 220170 525306 220226
rect 525374 220170 525430 220226
rect 525498 220170 525554 220226
rect 525622 220170 525678 220226
rect 525250 220046 525306 220102
rect 525374 220046 525430 220102
rect 525498 220046 525554 220102
rect 525622 220046 525678 220102
rect 525250 219922 525306 219978
rect 525374 219922 525430 219978
rect 525498 219922 525554 219978
rect 525622 219922 525678 219978
rect 528970 226294 529026 226350
rect 529094 226294 529150 226350
rect 529218 226294 529274 226350
rect 529342 226294 529398 226350
rect 528970 226170 529026 226226
rect 529094 226170 529150 226226
rect 529218 226170 529274 226226
rect 529342 226170 529398 226226
rect 528970 226046 529026 226102
rect 529094 226046 529150 226102
rect 529218 226046 529274 226102
rect 529342 226046 529398 226102
rect 528970 225922 529026 225978
rect 529094 225922 529150 225978
rect 529218 225922 529274 225978
rect 529342 225922 529398 225978
rect 543250 580294 543306 580350
rect 543374 580294 543430 580350
rect 543498 580294 543554 580350
rect 543622 580294 543678 580350
rect 543250 580170 543306 580226
rect 543374 580170 543430 580226
rect 543498 580170 543554 580226
rect 543622 580170 543678 580226
rect 543250 580046 543306 580102
rect 543374 580046 543430 580102
rect 543498 580046 543554 580102
rect 543622 580046 543678 580102
rect 543250 579922 543306 579978
rect 543374 579922 543430 579978
rect 543498 579922 543554 579978
rect 543622 579922 543678 579978
rect 543250 562294 543306 562350
rect 543374 562294 543430 562350
rect 543498 562294 543554 562350
rect 543622 562294 543678 562350
rect 543250 562170 543306 562226
rect 543374 562170 543430 562226
rect 543498 562170 543554 562226
rect 543622 562170 543678 562226
rect 543250 562046 543306 562102
rect 543374 562046 543430 562102
rect 543498 562046 543554 562102
rect 543622 562046 543678 562102
rect 543250 561922 543306 561978
rect 543374 561922 543430 561978
rect 543498 561922 543554 561978
rect 543622 561922 543678 561978
rect 543250 544294 543306 544350
rect 543374 544294 543430 544350
rect 543498 544294 543554 544350
rect 543622 544294 543678 544350
rect 543250 544170 543306 544226
rect 543374 544170 543430 544226
rect 543498 544170 543554 544226
rect 543622 544170 543678 544226
rect 543250 544046 543306 544102
rect 543374 544046 543430 544102
rect 543498 544046 543554 544102
rect 543622 544046 543678 544102
rect 543250 543922 543306 543978
rect 543374 543922 543430 543978
rect 543498 543922 543554 543978
rect 543622 543922 543678 543978
rect 543250 526294 543306 526350
rect 543374 526294 543430 526350
rect 543498 526294 543554 526350
rect 543622 526294 543678 526350
rect 543250 526170 543306 526226
rect 543374 526170 543430 526226
rect 543498 526170 543554 526226
rect 543622 526170 543678 526226
rect 543250 526046 543306 526102
rect 543374 526046 543430 526102
rect 543498 526046 543554 526102
rect 543622 526046 543678 526102
rect 543250 525922 543306 525978
rect 543374 525922 543430 525978
rect 543498 525922 543554 525978
rect 543622 525922 543678 525978
rect 543250 508294 543306 508350
rect 543374 508294 543430 508350
rect 543498 508294 543554 508350
rect 543622 508294 543678 508350
rect 543250 508170 543306 508226
rect 543374 508170 543430 508226
rect 543498 508170 543554 508226
rect 543622 508170 543678 508226
rect 543250 508046 543306 508102
rect 543374 508046 543430 508102
rect 543498 508046 543554 508102
rect 543622 508046 543678 508102
rect 543250 507922 543306 507978
rect 543374 507922 543430 507978
rect 543498 507922 543554 507978
rect 543622 507922 543678 507978
rect 543250 490294 543306 490350
rect 543374 490294 543430 490350
rect 543498 490294 543554 490350
rect 543622 490294 543678 490350
rect 543250 490170 543306 490226
rect 543374 490170 543430 490226
rect 543498 490170 543554 490226
rect 543622 490170 543678 490226
rect 543250 490046 543306 490102
rect 543374 490046 543430 490102
rect 543498 490046 543554 490102
rect 543622 490046 543678 490102
rect 543250 489922 543306 489978
rect 543374 489922 543430 489978
rect 543498 489922 543554 489978
rect 543622 489922 543678 489978
rect 543250 472294 543306 472350
rect 543374 472294 543430 472350
rect 543498 472294 543554 472350
rect 543622 472294 543678 472350
rect 543250 472170 543306 472226
rect 543374 472170 543430 472226
rect 543498 472170 543554 472226
rect 543622 472170 543678 472226
rect 543250 472046 543306 472102
rect 543374 472046 543430 472102
rect 543498 472046 543554 472102
rect 543622 472046 543678 472102
rect 543250 471922 543306 471978
rect 543374 471922 543430 471978
rect 543498 471922 543554 471978
rect 543622 471922 543678 471978
rect 543250 454294 543306 454350
rect 543374 454294 543430 454350
rect 543498 454294 543554 454350
rect 543622 454294 543678 454350
rect 543250 454170 543306 454226
rect 543374 454170 543430 454226
rect 543498 454170 543554 454226
rect 543622 454170 543678 454226
rect 543250 454046 543306 454102
rect 543374 454046 543430 454102
rect 543498 454046 543554 454102
rect 543622 454046 543678 454102
rect 543250 453922 543306 453978
rect 543374 453922 543430 453978
rect 543498 453922 543554 453978
rect 543622 453922 543678 453978
rect 543250 436294 543306 436350
rect 543374 436294 543430 436350
rect 543498 436294 543554 436350
rect 543622 436294 543678 436350
rect 543250 436170 543306 436226
rect 543374 436170 543430 436226
rect 543498 436170 543554 436226
rect 543622 436170 543678 436226
rect 543250 436046 543306 436102
rect 543374 436046 543430 436102
rect 543498 436046 543554 436102
rect 543622 436046 543678 436102
rect 543250 435922 543306 435978
rect 543374 435922 543430 435978
rect 543498 435922 543554 435978
rect 543622 435922 543678 435978
rect 543250 418294 543306 418350
rect 543374 418294 543430 418350
rect 543498 418294 543554 418350
rect 543622 418294 543678 418350
rect 543250 418170 543306 418226
rect 543374 418170 543430 418226
rect 543498 418170 543554 418226
rect 543622 418170 543678 418226
rect 543250 418046 543306 418102
rect 543374 418046 543430 418102
rect 543498 418046 543554 418102
rect 543622 418046 543678 418102
rect 543250 417922 543306 417978
rect 543374 417922 543430 417978
rect 543498 417922 543554 417978
rect 543622 417922 543678 417978
rect 543250 400294 543306 400350
rect 543374 400294 543430 400350
rect 543498 400294 543554 400350
rect 543622 400294 543678 400350
rect 543250 400170 543306 400226
rect 543374 400170 543430 400226
rect 543498 400170 543554 400226
rect 543622 400170 543678 400226
rect 543250 400046 543306 400102
rect 543374 400046 543430 400102
rect 543498 400046 543554 400102
rect 543622 400046 543678 400102
rect 543250 399922 543306 399978
rect 543374 399922 543430 399978
rect 543498 399922 543554 399978
rect 543622 399922 543678 399978
rect 543250 382294 543306 382350
rect 543374 382294 543430 382350
rect 543498 382294 543554 382350
rect 543622 382294 543678 382350
rect 543250 382170 543306 382226
rect 543374 382170 543430 382226
rect 543498 382170 543554 382226
rect 543622 382170 543678 382226
rect 543250 382046 543306 382102
rect 543374 382046 543430 382102
rect 543498 382046 543554 382102
rect 543622 382046 543678 382102
rect 543250 381922 543306 381978
rect 543374 381922 543430 381978
rect 543498 381922 543554 381978
rect 543622 381922 543678 381978
rect 543250 364294 543306 364350
rect 543374 364294 543430 364350
rect 543498 364294 543554 364350
rect 543622 364294 543678 364350
rect 543250 364170 543306 364226
rect 543374 364170 543430 364226
rect 543498 364170 543554 364226
rect 543622 364170 543678 364226
rect 543250 364046 543306 364102
rect 543374 364046 543430 364102
rect 543498 364046 543554 364102
rect 543622 364046 543678 364102
rect 543250 363922 543306 363978
rect 543374 363922 543430 363978
rect 543498 363922 543554 363978
rect 543622 363922 543678 363978
rect 543250 346294 543306 346350
rect 543374 346294 543430 346350
rect 543498 346294 543554 346350
rect 543622 346294 543678 346350
rect 543250 346170 543306 346226
rect 543374 346170 543430 346226
rect 543498 346170 543554 346226
rect 543622 346170 543678 346226
rect 543250 346046 543306 346102
rect 543374 346046 543430 346102
rect 543498 346046 543554 346102
rect 543622 346046 543678 346102
rect 543250 345922 543306 345978
rect 543374 345922 543430 345978
rect 543498 345922 543554 345978
rect 543622 345922 543678 345978
rect 543250 328294 543306 328350
rect 543374 328294 543430 328350
rect 543498 328294 543554 328350
rect 543622 328294 543678 328350
rect 543250 328170 543306 328226
rect 543374 328170 543430 328226
rect 543498 328170 543554 328226
rect 543622 328170 543678 328226
rect 543250 328046 543306 328102
rect 543374 328046 543430 328102
rect 543498 328046 543554 328102
rect 543622 328046 543678 328102
rect 543250 327922 543306 327978
rect 543374 327922 543430 327978
rect 543498 327922 543554 327978
rect 543622 327922 543678 327978
rect 543250 310294 543306 310350
rect 543374 310294 543430 310350
rect 543498 310294 543554 310350
rect 543622 310294 543678 310350
rect 543250 310170 543306 310226
rect 543374 310170 543430 310226
rect 543498 310170 543554 310226
rect 543622 310170 543678 310226
rect 543250 310046 543306 310102
rect 543374 310046 543430 310102
rect 543498 310046 543554 310102
rect 543622 310046 543678 310102
rect 543250 309922 543306 309978
rect 543374 309922 543430 309978
rect 543498 309922 543554 309978
rect 543622 309922 543678 309978
rect 543250 292294 543306 292350
rect 543374 292294 543430 292350
rect 543498 292294 543554 292350
rect 543622 292294 543678 292350
rect 543250 292170 543306 292226
rect 543374 292170 543430 292226
rect 543498 292170 543554 292226
rect 543622 292170 543678 292226
rect 543250 292046 543306 292102
rect 543374 292046 543430 292102
rect 543498 292046 543554 292102
rect 543622 292046 543678 292102
rect 543250 291922 543306 291978
rect 543374 291922 543430 291978
rect 543498 291922 543554 291978
rect 543622 291922 543678 291978
rect 543250 274294 543306 274350
rect 543374 274294 543430 274350
rect 543498 274294 543554 274350
rect 543622 274294 543678 274350
rect 543250 274170 543306 274226
rect 543374 274170 543430 274226
rect 543498 274170 543554 274226
rect 543622 274170 543678 274226
rect 543250 274046 543306 274102
rect 543374 274046 543430 274102
rect 543498 274046 543554 274102
rect 543622 274046 543678 274102
rect 543250 273922 543306 273978
rect 543374 273922 543430 273978
rect 543498 273922 543554 273978
rect 543622 273922 543678 273978
rect 543250 256294 543306 256350
rect 543374 256294 543430 256350
rect 543498 256294 543554 256350
rect 543622 256294 543678 256350
rect 543250 256170 543306 256226
rect 543374 256170 543430 256226
rect 543498 256170 543554 256226
rect 543622 256170 543678 256226
rect 543250 256046 543306 256102
rect 543374 256046 543430 256102
rect 543498 256046 543554 256102
rect 543622 256046 543678 256102
rect 543250 255922 543306 255978
rect 543374 255922 543430 255978
rect 543498 255922 543554 255978
rect 543622 255922 543678 255978
rect 543250 238294 543306 238350
rect 543374 238294 543430 238350
rect 543498 238294 543554 238350
rect 543622 238294 543678 238350
rect 543250 238170 543306 238226
rect 543374 238170 543430 238226
rect 543498 238170 543554 238226
rect 543622 238170 543678 238226
rect 543250 238046 543306 238102
rect 543374 238046 543430 238102
rect 543498 238046 543554 238102
rect 543622 238046 543678 238102
rect 543250 237922 543306 237978
rect 543374 237922 543430 237978
rect 543498 237922 543554 237978
rect 543622 237922 543678 237978
rect 543250 220294 543306 220350
rect 543374 220294 543430 220350
rect 543498 220294 543554 220350
rect 543622 220294 543678 220350
rect 543250 220170 543306 220226
rect 543374 220170 543430 220226
rect 543498 220170 543554 220226
rect 543622 220170 543678 220226
rect 543250 220046 543306 220102
rect 543374 220046 543430 220102
rect 543498 220046 543554 220102
rect 543622 220046 543678 220102
rect 543250 219922 543306 219978
rect 543374 219922 543430 219978
rect 543498 219922 543554 219978
rect 543622 219922 543678 219978
rect 546970 598116 547026 598172
rect 547094 598116 547150 598172
rect 547218 598116 547274 598172
rect 547342 598116 547398 598172
rect 546970 597992 547026 598048
rect 547094 597992 547150 598048
rect 547218 597992 547274 598048
rect 547342 597992 547398 598048
rect 546970 597868 547026 597924
rect 547094 597868 547150 597924
rect 547218 597868 547274 597924
rect 547342 597868 547398 597924
rect 546970 597744 547026 597800
rect 547094 597744 547150 597800
rect 547218 597744 547274 597800
rect 547342 597744 547398 597800
rect 546970 586294 547026 586350
rect 547094 586294 547150 586350
rect 547218 586294 547274 586350
rect 547342 586294 547398 586350
rect 546970 586170 547026 586226
rect 547094 586170 547150 586226
rect 547218 586170 547274 586226
rect 547342 586170 547398 586226
rect 546970 586046 547026 586102
rect 547094 586046 547150 586102
rect 547218 586046 547274 586102
rect 547342 586046 547398 586102
rect 546970 585922 547026 585978
rect 547094 585922 547150 585978
rect 547218 585922 547274 585978
rect 547342 585922 547398 585978
rect 546970 568294 547026 568350
rect 547094 568294 547150 568350
rect 547218 568294 547274 568350
rect 547342 568294 547398 568350
rect 546970 568170 547026 568226
rect 547094 568170 547150 568226
rect 547218 568170 547274 568226
rect 547342 568170 547398 568226
rect 546970 568046 547026 568102
rect 547094 568046 547150 568102
rect 547218 568046 547274 568102
rect 547342 568046 547398 568102
rect 546970 567922 547026 567978
rect 547094 567922 547150 567978
rect 547218 567922 547274 567978
rect 547342 567922 547398 567978
rect 546970 550294 547026 550350
rect 547094 550294 547150 550350
rect 547218 550294 547274 550350
rect 547342 550294 547398 550350
rect 546970 550170 547026 550226
rect 547094 550170 547150 550226
rect 547218 550170 547274 550226
rect 547342 550170 547398 550226
rect 546970 550046 547026 550102
rect 547094 550046 547150 550102
rect 547218 550046 547274 550102
rect 547342 550046 547398 550102
rect 546970 549922 547026 549978
rect 547094 549922 547150 549978
rect 547218 549922 547274 549978
rect 547342 549922 547398 549978
rect 546970 532294 547026 532350
rect 547094 532294 547150 532350
rect 547218 532294 547274 532350
rect 547342 532294 547398 532350
rect 546970 532170 547026 532226
rect 547094 532170 547150 532226
rect 547218 532170 547274 532226
rect 547342 532170 547398 532226
rect 546970 532046 547026 532102
rect 547094 532046 547150 532102
rect 547218 532046 547274 532102
rect 547342 532046 547398 532102
rect 546970 531922 547026 531978
rect 547094 531922 547150 531978
rect 547218 531922 547274 531978
rect 547342 531922 547398 531978
rect 546970 514294 547026 514350
rect 547094 514294 547150 514350
rect 547218 514294 547274 514350
rect 547342 514294 547398 514350
rect 546970 514170 547026 514226
rect 547094 514170 547150 514226
rect 547218 514170 547274 514226
rect 547342 514170 547398 514226
rect 546970 514046 547026 514102
rect 547094 514046 547150 514102
rect 547218 514046 547274 514102
rect 547342 514046 547398 514102
rect 546970 513922 547026 513978
rect 547094 513922 547150 513978
rect 547218 513922 547274 513978
rect 547342 513922 547398 513978
rect 546970 496294 547026 496350
rect 547094 496294 547150 496350
rect 547218 496294 547274 496350
rect 547342 496294 547398 496350
rect 546970 496170 547026 496226
rect 547094 496170 547150 496226
rect 547218 496170 547274 496226
rect 547342 496170 547398 496226
rect 546970 496046 547026 496102
rect 547094 496046 547150 496102
rect 547218 496046 547274 496102
rect 547342 496046 547398 496102
rect 546970 495922 547026 495978
rect 547094 495922 547150 495978
rect 547218 495922 547274 495978
rect 547342 495922 547398 495978
rect 561250 597156 561306 597212
rect 561374 597156 561430 597212
rect 561498 597156 561554 597212
rect 561622 597156 561678 597212
rect 561250 597032 561306 597088
rect 561374 597032 561430 597088
rect 561498 597032 561554 597088
rect 561622 597032 561678 597088
rect 561250 596908 561306 596964
rect 561374 596908 561430 596964
rect 561498 596908 561554 596964
rect 561622 596908 561678 596964
rect 561250 596784 561306 596840
rect 561374 596784 561430 596840
rect 561498 596784 561554 596840
rect 561622 596784 561678 596840
rect 561250 580294 561306 580350
rect 561374 580294 561430 580350
rect 561498 580294 561554 580350
rect 561622 580294 561678 580350
rect 561250 580170 561306 580226
rect 561374 580170 561430 580226
rect 561498 580170 561554 580226
rect 561622 580170 561678 580226
rect 561250 580046 561306 580102
rect 561374 580046 561430 580102
rect 561498 580046 561554 580102
rect 561622 580046 561678 580102
rect 561250 579922 561306 579978
rect 561374 579922 561430 579978
rect 561498 579922 561554 579978
rect 561622 579922 561678 579978
rect 561250 562294 561306 562350
rect 561374 562294 561430 562350
rect 561498 562294 561554 562350
rect 561622 562294 561678 562350
rect 561250 562170 561306 562226
rect 561374 562170 561430 562226
rect 561498 562170 561554 562226
rect 561622 562170 561678 562226
rect 561250 562046 561306 562102
rect 561374 562046 561430 562102
rect 561498 562046 561554 562102
rect 561622 562046 561678 562102
rect 561250 561922 561306 561978
rect 561374 561922 561430 561978
rect 561498 561922 561554 561978
rect 561622 561922 561678 561978
rect 561250 544294 561306 544350
rect 561374 544294 561430 544350
rect 561498 544294 561554 544350
rect 561622 544294 561678 544350
rect 561250 544170 561306 544226
rect 561374 544170 561430 544226
rect 561498 544170 561554 544226
rect 561622 544170 561678 544226
rect 561250 544046 561306 544102
rect 561374 544046 561430 544102
rect 561498 544046 561554 544102
rect 561622 544046 561678 544102
rect 561250 543922 561306 543978
rect 561374 543922 561430 543978
rect 561498 543922 561554 543978
rect 561622 543922 561678 543978
rect 561250 526294 561306 526350
rect 561374 526294 561430 526350
rect 561498 526294 561554 526350
rect 561622 526294 561678 526350
rect 561250 526170 561306 526226
rect 561374 526170 561430 526226
rect 561498 526170 561554 526226
rect 561622 526170 561678 526226
rect 561250 526046 561306 526102
rect 561374 526046 561430 526102
rect 561498 526046 561554 526102
rect 561622 526046 561678 526102
rect 561250 525922 561306 525978
rect 561374 525922 561430 525978
rect 561498 525922 561554 525978
rect 561622 525922 561678 525978
rect 561250 508294 561306 508350
rect 561374 508294 561430 508350
rect 561498 508294 561554 508350
rect 561622 508294 561678 508350
rect 561250 508170 561306 508226
rect 561374 508170 561430 508226
rect 561498 508170 561554 508226
rect 561622 508170 561678 508226
rect 561250 508046 561306 508102
rect 561374 508046 561430 508102
rect 561498 508046 561554 508102
rect 561622 508046 561678 508102
rect 561250 507922 561306 507978
rect 561374 507922 561430 507978
rect 561498 507922 561554 507978
rect 561622 507922 561678 507978
rect 564970 598116 565026 598172
rect 565094 598116 565150 598172
rect 565218 598116 565274 598172
rect 565342 598116 565398 598172
rect 564970 597992 565026 598048
rect 565094 597992 565150 598048
rect 565218 597992 565274 598048
rect 565342 597992 565398 598048
rect 564970 597868 565026 597924
rect 565094 597868 565150 597924
rect 565218 597868 565274 597924
rect 565342 597868 565398 597924
rect 564970 597744 565026 597800
rect 565094 597744 565150 597800
rect 565218 597744 565274 597800
rect 565342 597744 565398 597800
rect 564970 586294 565026 586350
rect 565094 586294 565150 586350
rect 565218 586294 565274 586350
rect 565342 586294 565398 586350
rect 564970 586170 565026 586226
rect 565094 586170 565150 586226
rect 565218 586170 565274 586226
rect 565342 586170 565398 586226
rect 564970 586046 565026 586102
rect 565094 586046 565150 586102
rect 565218 586046 565274 586102
rect 565342 586046 565398 586102
rect 564970 585922 565026 585978
rect 565094 585922 565150 585978
rect 565218 585922 565274 585978
rect 565342 585922 565398 585978
rect 564970 568294 565026 568350
rect 565094 568294 565150 568350
rect 565218 568294 565274 568350
rect 565342 568294 565398 568350
rect 564970 568170 565026 568226
rect 565094 568170 565150 568226
rect 565218 568170 565274 568226
rect 565342 568170 565398 568226
rect 564970 568046 565026 568102
rect 565094 568046 565150 568102
rect 565218 568046 565274 568102
rect 565342 568046 565398 568102
rect 564970 567922 565026 567978
rect 565094 567922 565150 567978
rect 565218 567922 565274 567978
rect 565342 567922 565398 567978
rect 564970 550294 565026 550350
rect 565094 550294 565150 550350
rect 565218 550294 565274 550350
rect 565342 550294 565398 550350
rect 564970 550170 565026 550226
rect 565094 550170 565150 550226
rect 565218 550170 565274 550226
rect 565342 550170 565398 550226
rect 564970 550046 565026 550102
rect 565094 550046 565150 550102
rect 565218 550046 565274 550102
rect 565342 550046 565398 550102
rect 564970 549922 565026 549978
rect 565094 549922 565150 549978
rect 565218 549922 565274 549978
rect 565342 549922 565398 549978
rect 564970 532294 565026 532350
rect 565094 532294 565150 532350
rect 565218 532294 565274 532350
rect 565342 532294 565398 532350
rect 564970 532170 565026 532226
rect 565094 532170 565150 532226
rect 565218 532170 565274 532226
rect 565342 532170 565398 532226
rect 564970 532046 565026 532102
rect 565094 532046 565150 532102
rect 565218 532046 565274 532102
rect 565342 532046 565398 532102
rect 564970 531922 565026 531978
rect 565094 531922 565150 531978
rect 565218 531922 565274 531978
rect 565342 531922 565398 531978
rect 564970 514294 565026 514350
rect 565094 514294 565150 514350
rect 565218 514294 565274 514350
rect 565342 514294 565398 514350
rect 564970 514170 565026 514226
rect 565094 514170 565150 514226
rect 565218 514170 565274 514226
rect 565342 514170 565398 514226
rect 564970 514046 565026 514102
rect 565094 514046 565150 514102
rect 565218 514046 565274 514102
rect 565342 514046 565398 514102
rect 564970 513922 565026 513978
rect 565094 513922 565150 513978
rect 565218 513922 565274 513978
rect 565342 513922 565398 513978
rect 579250 597156 579306 597212
rect 579374 597156 579430 597212
rect 579498 597156 579554 597212
rect 579622 597156 579678 597212
rect 579250 597032 579306 597088
rect 579374 597032 579430 597088
rect 579498 597032 579554 597088
rect 579622 597032 579678 597088
rect 579250 596908 579306 596964
rect 579374 596908 579430 596964
rect 579498 596908 579554 596964
rect 579622 596908 579678 596964
rect 579250 596784 579306 596840
rect 579374 596784 579430 596840
rect 579498 596784 579554 596840
rect 579622 596784 579678 596840
rect 579250 580294 579306 580350
rect 579374 580294 579430 580350
rect 579498 580294 579554 580350
rect 579622 580294 579678 580350
rect 579250 580170 579306 580226
rect 579374 580170 579430 580226
rect 579498 580170 579554 580226
rect 579622 580170 579678 580226
rect 579250 580046 579306 580102
rect 579374 580046 579430 580102
rect 579498 580046 579554 580102
rect 579622 580046 579678 580102
rect 579250 579922 579306 579978
rect 579374 579922 579430 579978
rect 579498 579922 579554 579978
rect 579622 579922 579678 579978
rect 579250 562294 579306 562350
rect 579374 562294 579430 562350
rect 579498 562294 579554 562350
rect 579622 562294 579678 562350
rect 579250 562170 579306 562226
rect 579374 562170 579430 562226
rect 579498 562170 579554 562226
rect 579622 562170 579678 562226
rect 579250 562046 579306 562102
rect 579374 562046 579430 562102
rect 579498 562046 579554 562102
rect 579622 562046 579678 562102
rect 579250 561922 579306 561978
rect 579374 561922 579430 561978
rect 579498 561922 579554 561978
rect 579622 561922 579678 561978
rect 579250 544294 579306 544350
rect 579374 544294 579430 544350
rect 579498 544294 579554 544350
rect 579622 544294 579678 544350
rect 579250 544170 579306 544226
rect 579374 544170 579430 544226
rect 579498 544170 579554 544226
rect 579622 544170 579678 544226
rect 579250 544046 579306 544102
rect 579374 544046 579430 544102
rect 579498 544046 579554 544102
rect 579622 544046 579678 544102
rect 579250 543922 579306 543978
rect 579374 543922 579430 543978
rect 579498 543922 579554 543978
rect 579622 543922 579678 543978
rect 579250 526294 579306 526350
rect 579374 526294 579430 526350
rect 579498 526294 579554 526350
rect 579622 526294 579678 526350
rect 579250 526170 579306 526226
rect 579374 526170 579430 526226
rect 579498 526170 579554 526226
rect 579622 526170 579678 526226
rect 579250 526046 579306 526102
rect 579374 526046 579430 526102
rect 579498 526046 579554 526102
rect 579622 526046 579678 526102
rect 579250 525922 579306 525978
rect 579374 525922 579430 525978
rect 579498 525922 579554 525978
rect 579622 525922 579678 525978
rect 579250 508294 579306 508350
rect 579374 508294 579430 508350
rect 579498 508294 579554 508350
rect 579622 508294 579678 508350
rect 579250 508170 579306 508226
rect 579374 508170 579430 508226
rect 579498 508170 579554 508226
rect 579622 508170 579678 508226
rect 579250 508046 579306 508102
rect 579374 508046 579430 508102
rect 579498 508046 579554 508102
rect 579622 508046 579678 508102
rect 579250 507922 579306 507978
rect 579374 507922 579430 507978
rect 579498 507922 579554 507978
rect 579622 507922 579678 507978
rect 568058 496294 568114 496350
rect 568182 496294 568238 496350
rect 568058 496170 568114 496226
rect 568182 496170 568238 496226
rect 568058 496046 568114 496102
rect 568182 496046 568238 496102
rect 568058 495922 568114 495978
rect 568182 495922 568238 495978
rect 574862 496294 574918 496350
rect 574986 496294 575042 496350
rect 574862 496170 574918 496226
rect 574986 496170 575042 496226
rect 574862 496046 574918 496102
rect 574986 496046 575042 496102
rect 574862 495922 574918 495978
rect 574986 495922 575042 495978
rect 561250 490294 561306 490350
rect 561374 490294 561430 490350
rect 561498 490294 561554 490350
rect 561622 490294 561678 490350
rect 561250 490170 561306 490226
rect 561374 490170 561430 490226
rect 561498 490170 561554 490226
rect 561622 490170 561678 490226
rect 561250 490046 561306 490102
rect 561374 490046 561430 490102
rect 561498 490046 561554 490102
rect 561622 490046 561678 490102
rect 561250 489922 561306 489978
rect 561374 489922 561430 489978
rect 561498 489922 561554 489978
rect 561622 489922 561678 489978
rect 564656 490294 564712 490350
rect 564780 490294 564836 490350
rect 564656 490170 564712 490226
rect 564780 490170 564836 490226
rect 564656 490046 564712 490102
rect 564780 490046 564836 490102
rect 564656 489922 564712 489978
rect 564780 489922 564836 489978
rect 571460 490294 571516 490350
rect 571584 490294 571640 490350
rect 571460 490170 571516 490226
rect 571584 490170 571640 490226
rect 571460 490046 571516 490102
rect 571584 490046 571640 490102
rect 571460 489922 571516 489978
rect 571584 489922 571640 489978
rect 578264 490294 578320 490350
rect 578388 490294 578444 490350
rect 578264 490170 578320 490226
rect 578388 490170 578444 490226
rect 578264 490046 578320 490102
rect 578388 490046 578444 490102
rect 578264 489922 578320 489978
rect 578388 489922 578444 489978
rect 582970 598116 583026 598172
rect 583094 598116 583150 598172
rect 583218 598116 583274 598172
rect 583342 598116 583398 598172
rect 582970 597992 583026 598048
rect 583094 597992 583150 598048
rect 583218 597992 583274 598048
rect 583342 597992 583398 598048
rect 582970 597868 583026 597924
rect 583094 597868 583150 597924
rect 583218 597868 583274 597924
rect 583342 597868 583398 597924
rect 582970 597744 583026 597800
rect 583094 597744 583150 597800
rect 583218 597744 583274 597800
rect 583342 597744 583398 597800
rect 597456 598116 597512 598172
rect 597580 598116 597636 598172
rect 597704 598116 597760 598172
rect 597828 598116 597884 598172
rect 597456 597992 597512 598048
rect 597580 597992 597636 598048
rect 597704 597992 597760 598048
rect 597828 597992 597884 598048
rect 597456 597868 597512 597924
rect 597580 597868 597636 597924
rect 597704 597868 597760 597924
rect 597828 597868 597884 597924
rect 597456 597744 597512 597800
rect 597580 597744 597636 597800
rect 597704 597744 597760 597800
rect 597828 597744 597884 597800
rect 582970 586294 583026 586350
rect 583094 586294 583150 586350
rect 583218 586294 583274 586350
rect 583342 586294 583398 586350
rect 582970 586170 583026 586226
rect 583094 586170 583150 586226
rect 583218 586170 583274 586226
rect 583342 586170 583398 586226
rect 582970 586046 583026 586102
rect 583094 586046 583150 586102
rect 583218 586046 583274 586102
rect 583342 586046 583398 586102
rect 582970 585922 583026 585978
rect 583094 585922 583150 585978
rect 583218 585922 583274 585978
rect 583342 585922 583398 585978
rect 582970 568294 583026 568350
rect 583094 568294 583150 568350
rect 583218 568294 583274 568350
rect 583342 568294 583398 568350
rect 582970 568170 583026 568226
rect 583094 568170 583150 568226
rect 583218 568170 583274 568226
rect 583342 568170 583398 568226
rect 582970 568046 583026 568102
rect 583094 568046 583150 568102
rect 583218 568046 583274 568102
rect 583342 568046 583398 568102
rect 582970 567922 583026 567978
rect 583094 567922 583150 567978
rect 583218 567922 583274 567978
rect 583342 567922 583398 567978
rect 582970 550294 583026 550350
rect 583094 550294 583150 550350
rect 583218 550294 583274 550350
rect 583342 550294 583398 550350
rect 582970 550170 583026 550226
rect 583094 550170 583150 550226
rect 583218 550170 583274 550226
rect 583342 550170 583398 550226
rect 582970 550046 583026 550102
rect 583094 550046 583150 550102
rect 583218 550046 583274 550102
rect 583342 550046 583398 550102
rect 582970 549922 583026 549978
rect 583094 549922 583150 549978
rect 583218 549922 583274 549978
rect 583342 549922 583398 549978
rect 582970 532294 583026 532350
rect 583094 532294 583150 532350
rect 583218 532294 583274 532350
rect 583342 532294 583398 532350
rect 582970 532170 583026 532226
rect 583094 532170 583150 532226
rect 583218 532170 583274 532226
rect 583342 532170 583398 532226
rect 582970 532046 583026 532102
rect 583094 532046 583150 532102
rect 583218 532046 583274 532102
rect 583342 532046 583398 532102
rect 582970 531922 583026 531978
rect 583094 531922 583150 531978
rect 583218 531922 583274 531978
rect 583342 531922 583398 531978
rect 582970 514294 583026 514350
rect 583094 514294 583150 514350
rect 583218 514294 583274 514350
rect 583342 514294 583398 514350
rect 582970 514170 583026 514226
rect 583094 514170 583150 514226
rect 583218 514170 583274 514226
rect 583342 514170 583398 514226
rect 582970 514046 583026 514102
rect 583094 514046 583150 514102
rect 583218 514046 583274 514102
rect 583342 514046 583398 514102
rect 582970 513922 583026 513978
rect 583094 513922 583150 513978
rect 583218 513922 583274 513978
rect 583342 513922 583398 513978
rect 581666 496294 581722 496350
rect 581790 496294 581846 496350
rect 581666 496170 581722 496226
rect 581790 496170 581846 496226
rect 581666 496046 581722 496102
rect 581790 496046 581846 496102
rect 581666 495922 581722 495978
rect 581790 495922 581846 495978
rect 596496 597156 596552 597212
rect 596620 597156 596676 597212
rect 596744 597156 596800 597212
rect 596868 597156 596924 597212
rect 596496 597032 596552 597088
rect 596620 597032 596676 597088
rect 596744 597032 596800 597088
rect 596868 597032 596924 597088
rect 596496 596908 596552 596964
rect 596620 596908 596676 596964
rect 596744 596908 596800 596964
rect 596868 596908 596924 596964
rect 596496 596784 596552 596840
rect 596620 596784 596676 596840
rect 596744 596784 596800 596840
rect 596868 596784 596924 596840
rect 596496 580294 596552 580350
rect 596620 580294 596676 580350
rect 596744 580294 596800 580350
rect 596868 580294 596924 580350
rect 596496 580170 596552 580226
rect 596620 580170 596676 580226
rect 596744 580170 596800 580226
rect 596868 580170 596924 580226
rect 596496 580046 596552 580102
rect 596620 580046 596676 580102
rect 596744 580046 596800 580102
rect 596868 580046 596924 580102
rect 596496 579922 596552 579978
rect 596620 579922 596676 579978
rect 596744 579922 596800 579978
rect 596868 579922 596924 579978
rect 596496 562294 596552 562350
rect 596620 562294 596676 562350
rect 596744 562294 596800 562350
rect 596868 562294 596924 562350
rect 596496 562170 596552 562226
rect 596620 562170 596676 562226
rect 596744 562170 596800 562226
rect 596868 562170 596924 562226
rect 596496 562046 596552 562102
rect 596620 562046 596676 562102
rect 596744 562046 596800 562102
rect 596868 562046 596924 562102
rect 596496 561922 596552 561978
rect 596620 561922 596676 561978
rect 596744 561922 596800 561978
rect 596868 561922 596924 561978
rect 596496 544294 596552 544350
rect 596620 544294 596676 544350
rect 596744 544294 596800 544350
rect 596868 544294 596924 544350
rect 596496 544170 596552 544226
rect 596620 544170 596676 544226
rect 596744 544170 596800 544226
rect 596868 544170 596924 544226
rect 596496 544046 596552 544102
rect 596620 544046 596676 544102
rect 596744 544046 596800 544102
rect 596868 544046 596924 544102
rect 596496 543922 596552 543978
rect 596620 543922 596676 543978
rect 596744 543922 596800 543978
rect 596868 543922 596924 543978
rect 596496 526294 596552 526350
rect 596620 526294 596676 526350
rect 596744 526294 596800 526350
rect 596868 526294 596924 526350
rect 596496 526170 596552 526226
rect 596620 526170 596676 526226
rect 596744 526170 596800 526226
rect 596868 526170 596924 526226
rect 596496 526046 596552 526102
rect 596620 526046 596676 526102
rect 596744 526046 596800 526102
rect 596868 526046 596924 526102
rect 596496 525922 596552 525978
rect 596620 525922 596676 525978
rect 596744 525922 596800 525978
rect 596868 525922 596924 525978
rect 596496 508294 596552 508350
rect 596620 508294 596676 508350
rect 596744 508294 596800 508350
rect 596868 508294 596924 508350
rect 596496 508170 596552 508226
rect 596620 508170 596676 508226
rect 596744 508170 596800 508226
rect 596868 508170 596924 508226
rect 596496 508046 596552 508102
rect 596620 508046 596676 508102
rect 596744 508046 596800 508102
rect 596868 508046 596924 508102
rect 596496 507922 596552 507978
rect 596620 507922 596676 507978
rect 596744 507922 596800 507978
rect 596868 507922 596924 507978
rect 582970 496294 583026 496350
rect 583094 496294 583150 496350
rect 583218 496294 583274 496350
rect 583342 496294 583398 496350
rect 582970 496170 583026 496226
rect 583094 496170 583150 496226
rect 583218 496170 583274 496226
rect 583342 496170 583398 496226
rect 582970 496046 583026 496102
rect 583094 496046 583150 496102
rect 583218 496046 583274 496102
rect 583342 496046 583398 496102
rect 582970 495922 583026 495978
rect 583094 495922 583150 495978
rect 583218 495922 583274 495978
rect 583342 495922 583398 495978
rect 579250 490294 579306 490350
rect 579374 490294 579430 490350
rect 579498 490294 579554 490350
rect 579622 490294 579678 490350
rect 579250 490170 579306 490226
rect 579374 490170 579430 490226
rect 579498 490170 579554 490226
rect 579622 490170 579678 490226
rect 579250 490046 579306 490102
rect 579374 490046 579430 490102
rect 579498 490046 579554 490102
rect 579622 490046 579678 490102
rect 579250 489922 579306 489978
rect 579374 489922 579430 489978
rect 579498 489922 579554 489978
rect 579622 489922 579678 489978
rect 588470 496294 588526 496350
rect 588594 496294 588650 496350
rect 588470 496170 588526 496226
rect 588594 496170 588650 496226
rect 588470 496046 588526 496102
rect 588594 496046 588650 496102
rect 588470 495922 588526 495978
rect 588594 495922 588650 495978
rect 585068 490294 585124 490350
rect 585192 490294 585248 490350
rect 585068 490170 585124 490226
rect 585192 490170 585248 490226
rect 585068 490046 585124 490102
rect 585192 490046 585248 490102
rect 585068 489922 585124 489978
rect 585192 489922 585248 489978
rect 596496 490294 596552 490350
rect 596620 490294 596676 490350
rect 596744 490294 596800 490350
rect 596868 490294 596924 490350
rect 596496 490170 596552 490226
rect 596620 490170 596676 490226
rect 596744 490170 596800 490226
rect 596868 490170 596924 490226
rect 596496 490046 596552 490102
rect 596620 490046 596676 490102
rect 596744 490046 596800 490102
rect 596868 490046 596924 490102
rect 596496 489922 596552 489978
rect 596620 489922 596676 489978
rect 596744 489922 596800 489978
rect 596868 489922 596924 489978
rect 546970 478294 547026 478350
rect 547094 478294 547150 478350
rect 547218 478294 547274 478350
rect 547342 478294 547398 478350
rect 546970 478170 547026 478226
rect 547094 478170 547150 478226
rect 547218 478170 547274 478226
rect 547342 478170 547398 478226
rect 546970 478046 547026 478102
rect 547094 478046 547150 478102
rect 547218 478046 547274 478102
rect 547342 478046 547398 478102
rect 546970 477922 547026 477978
rect 547094 477922 547150 477978
rect 547218 477922 547274 477978
rect 547342 477922 547398 477978
rect 568058 478294 568114 478350
rect 568182 478294 568238 478350
rect 568058 478170 568114 478226
rect 568182 478170 568238 478226
rect 568058 478046 568114 478102
rect 568182 478046 568238 478102
rect 568058 477922 568114 477978
rect 568182 477922 568238 477978
rect 574862 478294 574918 478350
rect 574986 478294 575042 478350
rect 574862 478170 574918 478226
rect 574986 478170 575042 478226
rect 574862 478046 574918 478102
rect 574986 478046 575042 478102
rect 574862 477922 574918 477978
rect 574986 477922 575042 477978
rect 581666 478294 581722 478350
rect 581790 478294 581846 478350
rect 581666 478170 581722 478226
rect 581790 478170 581846 478226
rect 581666 478046 581722 478102
rect 581790 478046 581846 478102
rect 581666 477922 581722 477978
rect 581790 477922 581846 477978
rect 588470 478294 588526 478350
rect 588594 478294 588650 478350
rect 588470 478170 588526 478226
rect 588594 478170 588650 478226
rect 588470 478046 588526 478102
rect 588594 478046 588650 478102
rect 588470 477922 588526 477978
rect 588594 477922 588650 477978
rect 564656 472294 564712 472350
rect 564780 472294 564836 472350
rect 564656 472170 564712 472226
rect 564780 472170 564836 472226
rect 564656 472046 564712 472102
rect 564780 472046 564836 472102
rect 564656 471922 564712 471978
rect 564780 471922 564836 471978
rect 571460 472294 571516 472350
rect 571584 472294 571640 472350
rect 571460 472170 571516 472226
rect 571584 472170 571640 472226
rect 571460 472046 571516 472102
rect 571584 472046 571640 472102
rect 571460 471922 571516 471978
rect 571584 471922 571640 471978
rect 578264 472294 578320 472350
rect 578388 472294 578444 472350
rect 578264 472170 578320 472226
rect 578388 472170 578444 472226
rect 578264 472046 578320 472102
rect 578388 472046 578444 472102
rect 578264 471922 578320 471978
rect 578388 471922 578444 471978
rect 585068 472294 585124 472350
rect 585192 472294 585248 472350
rect 585068 472170 585124 472226
rect 585192 472170 585248 472226
rect 585068 472046 585124 472102
rect 585192 472046 585248 472102
rect 585068 471922 585124 471978
rect 585192 471922 585248 471978
rect 596496 472294 596552 472350
rect 596620 472294 596676 472350
rect 596744 472294 596800 472350
rect 596868 472294 596924 472350
rect 596496 472170 596552 472226
rect 596620 472170 596676 472226
rect 596744 472170 596800 472226
rect 596868 472170 596924 472226
rect 596496 472046 596552 472102
rect 596620 472046 596676 472102
rect 596744 472046 596800 472102
rect 596868 472046 596924 472102
rect 596496 471922 596552 471978
rect 596620 471922 596676 471978
rect 596744 471922 596800 471978
rect 596868 471922 596924 471978
rect 546970 460294 547026 460350
rect 547094 460294 547150 460350
rect 547218 460294 547274 460350
rect 547342 460294 547398 460350
rect 546970 460170 547026 460226
rect 547094 460170 547150 460226
rect 547218 460170 547274 460226
rect 547342 460170 547398 460226
rect 546970 460046 547026 460102
rect 547094 460046 547150 460102
rect 547218 460046 547274 460102
rect 547342 460046 547398 460102
rect 546970 459922 547026 459978
rect 547094 459922 547150 459978
rect 547218 459922 547274 459978
rect 547342 459922 547398 459978
rect 546970 442294 547026 442350
rect 547094 442294 547150 442350
rect 547218 442294 547274 442350
rect 547342 442294 547398 442350
rect 546970 442170 547026 442226
rect 547094 442170 547150 442226
rect 547218 442170 547274 442226
rect 547342 442170 547398 442226
rect 546970 442046 547026 442102
rect 547094 442046 547150 442102
rect 547218 442046 547274 442102
rect 547342 442046 547398 442102
rect 546970 441922 547026 441978
rect 547094 441922 547150 441978
rect 547218 441922 547274 441978
rect 547342 441922 547398 441978
rect 546970 424294 547026 424350
rect 547094 424294 547150 424350
rect 547218 424294 547274 424350
rect 547342 424294 547398 424350
rect 546970 424170 547026 424226
rect 547094 424170 547150 424226
rect 547218 424170 547274 424226
rect 547342 424170 547398 424226
rect 546970 424046 547026 424102
rect 547094 424046 547150 424102
rect 547218 424046 547274 424102
rect 547342 424046 547398 424102
rect 546970 423922 547026 423978
rect 547094 423922 547150 423978
rect 547218 423922 547274 423978
rect 547342 423922 547398 423978
rect 546970 406294 547026 406350
rect 547094 406294 547150 406350
rect 547218 406294 547274 406350
rect 547342 406294 547398 406350
rect 546970 406170 547026 406226
rect 547094 406170 547150 406226
rect 547218 406170 547274 406226
rect 547342 406170 547398 406226
rect 546970 406046 547026 406102
rect 547094 406046 547150 406102
rect 547218 406046 547274 406102
rect 547342 406046 547398 406102
rect 546970 405922 547026 405978
rect 547094 405922 547150 405978
rect 547218 405922 547274 405978
rect 547342 405922 547398 405978
rect 546970 388294 547026 388350
rect 547094 388294 547150 388350
rect 547218 388294 547274 388350
rect 547342 388294 547398 388350
rect 546970 388170 547026 388226
rect 547094 388170 547150 388226
rect 547218 388170 547274 388226
rect 547342 388170 547398 388226
rect 546970 388046 547026 388102
rect 547094 388046 547150 388102
rect 547218 388046 547274 388102
rect 547342 388046 547398 388102
rect 546970 387922 547026 387978
rect 547094 387922 547150 387978
rect 547218 387922 547274 387978
rect 547342 387922 547398 387978
rect 546970 370294 547026 370350
rect 547094 370294 547150 370350
rect 547218 370294 547274 370350
rect 547342 370294 547398 370350
rect 546970 370170 547026 370226
rect 547094 370170 547150 370226
rect 547218 370170 547274 370226
rect 547342 370170 547398 370226
rect 546970 370046 547026 370102
rect 547094 370046 547150 370102
rect 547218 370046 547274 370102
rect 547342 370046 547398 370102
rect 546970 369922 547026 369978
rect 547094 369922 547150 369978
rect 547218 369922 547274 369978
rect 547342 369922 547398 369978
rect 546970 352294 547026 352350
rect 547094 352294 547150 352350
rect 547218 352294 547274 352350
rect 547342 352294 547398 352350
rect 546970 352170 547026 352226
rect 547094 352170 547150 352226
rect 547218 352170 547274 352226
rect 547342 352170 547398 352226
rect 546970 352046 547026 352102
rect 547094 352046 547150 352102
rect 547218 352046 547274 352102
rect 547342 352046 547398 352102
rect 546970 351922 547026 351978
rect 547094 351922 547150 351978
rect 547218 351922 547274 351978
rect 547342 351922 547398 351978
rect 546970 334294 547026 334350
rect 547094 334294 547150 334350
rect 547218 334294 547274 334350
rect 547342 334294 547398 334350
rect 546970 334170 547026 334226
rect 547094 334170 547150 334226
rect 547218 334170 547274 334226
rect 547342 334170 547398 334226
rect 546970 334046 547026 334102
rect 547094 334046 547150 334102
rect 547218 334046 547274 334102
rect 547342 334046 547398 334102
rect 546970 333922 547026 333978
rect 547094 333922 547150 333978
rect 547218 333922 547274 333978
rect 547342 333922 547398 333978
rect 546970 316294 547026 316350
rect 547094 316294 547150 316350
rect 547218 316294 547274 316350
rect 547342 316294 547398 316350
rect 546970 316170 547026 316226
rect 547094 316170 547150 316226
rect 547218 316170 547274 316226
rect 547342 316170 547398 316226
rect 546970 316046 547026 316102
rect 547094 316046 547150 316102
rect 547218 316046 547274 316102
rect 547342 316046 547398 316102
rect 546970 315922 547026 315978
rect 547094 315922 547150 315978
rect 547218 315922 547274 315978
rect 547342 315922 547398 315978
rect 546970 298294 547026 298350
rect 547094 298294 547150 298350
rect 547218 298294 547274 298350
rect 547342 298294 547398 298350
rect 546970 298170 547026 298226
rect 547094 298170 547150 298226
rect 547218 298170 547274 298226
rect 547342 298170 547398 298226
rect 546970 298046 547026 298102
rect 547094 298046 547150 298102
rect 547218 298046 547274 298102
rect 547342 298046 547398 298102
rect 546970 297922 547026 297978
rect 547094 297922 547150 297978
rect 547218 297922 547274 297978
rect 547342 297922 547398 297978
rect 546970 280294 547026 280350
rect 547094 280294 547150 280350
rect 547218 280294 547274 280350
rect 547342 280294 547398 280350
rect 546970 280170 547026 280226
rect 547094 280170 547150 280226
rect 547218 280170 547274 280226
rect 547342 280170 547398 280226
rect 546970 280046 547026 280102
rect 547094 280046 547150 280102
rect 547218 280046 547274 280102
rect 547342 280046 547398 280102
rect 546970 279922 547026 279978
rect 547094 279922 547150 279978
rect 547218 279922 547274 279978
rect 547342 279922 547398 279978
rect 546970 262294 547026 262350
rect 547094 262294 547150 262350
rect 547218 262294 547274 262350
rect 547342 262294 547398 262350
rect 546970 262170 547026 262226
rect 547094 262170 547150 262226
rect 547218 262170 547274 262226
rect 547342 262170 547398 262226
rect 546970 262046 547026 262102
rect 547094 262046 547150 262102
rect 547218 262046 547274 262102
rect 547342 262046 547398 262102
rect 546970 261922 547026 261978
rect 547094 261922 547150 261978
rect 547218 261922 547274 261978
rect 547342 261922 547398 261978
rect 546970 244294 547026 244350
rect 547094 244294 547150 244350
rect 547218 244294 547274 244350
rect 547342 244294 547398 244350
rect 546970 244170 547026 244226
rect 547094 244170 547150 244226
rect 547218 244170 547274 244226
rect 547342 244170 547398 244226
rect 546970 244046 547026 244102
rect 547094 244046 547150 244102
rect 547218 244046 547274 244102
rect 547342 244046 547398 244102
rect 546970 243922 547026 243978
rect 547094 243922 547150 243978
rect 547218 243922 547274 243978
rect 547342 243922 547398 243978
rect 546970 226294 547026 226350
rect 547094 226294 547150 226350
rect 547218 226294 547274 226350
rect 547342 226294 547398 226350
rect 546970 226170 547026 226226
rect 547094 226170 547150 226226
rect 547218 226170 547274 226226
rect 547342 226170 547398 226226
rect 546970 226046 547026 226102
rect 547094 226046 547150 226102
rect 547218 226046 547274 226102
rect 547342 226046 547398 226102
rect 546970 225922 547026 225978
rect 547094 225922 547150 225978
rect 547218 225922 547274 225978
rect 547342 225922 547398 225978
rect 348970 208294 349026 208350
rect 349094 208294 349150 208350
rect 349218 208294 349274 208350
rect 349342 208294 349398 208350
rect 348970 208170 349026 208226
rect 349094 208170 349150 208226
rect 349218 208170 349274 208226
rect 349342 208170 349398 208226
rect 348970 208046 349026 208102
rect 349094 208046 349150 208102
rect 349218 208046 349274 208102
rect 349342 208046 349398 208102
rect 348970 207922 349026 207978
rect 349094 207922 349150 207978
rect 349218 207922 349274 207978
rect 349342 207922 349398 207978
rect 364022 208356 364078 208412
rect 364146 208356 364202 208412
rect 364270 208356 364326 208412
rect 364394 208356 364450 208412
rect 364518 208356 364574 208412
rect 364642 208356 364698 208412
rect 364766 208356 364822 208412
rect 364890 208356 364946 208412
rect 365014 208356 365070 208412
rect 365138 208356 365194 208412
rect 364022 208232 364078 208288
rect 364146 208232 364202 208288
rect 364270 208232 364326 208288
rect 364394 208232 364450 208288
rect 364518 208232 364574 208288
rect 364642 208232 364698 208288
rect 364766 208232 364822 208288
rect 364890 208232 364946 208288
rect 365014 208232 365070 208288
rect 365138 208232 365194 208288
rect 364022 208108 364078 208164
rect 364146 208108 364202 208164
rect 364270 208108 364326 208164
rect 364394 208108 364450 208164
rect 364518 208108 364574 208164
rect 364642 208108 364698 208164
rect 364766 208108 364822 208164
rect 364890 208108 364946 208164
rect 365014 208108 365070 208164
rect 365138 208108 365194 208164
rect 364022 207984 364078 208040
rect 364146 207984 364202 208040
rect 364270 207984 364326 208040
rect 364394 207984 364450 208040
rect 364518 207984 364574 208040
rect 364642 207984 364698 208040
rect 364766 207984 364822 208040
rect 364890 207984 364946 208040
rect 365014 207984 365070 208040
rect 365138 207984 365194 208040
rect 364022 207860 364078 207916
rect 364146 207860 364202 207916
rect 364270 207860 364326 207916
rect 364394 207860 364450 207916
rect 364518 207860 364574 207916
rect 364642 207860 364698 207916
rect 364766 207860 364822 207916
rect 364890 207860 364946 207916
rect 365014 207860 365070 207916
rect 365138 207860 365194 207916
rect 384022 208356 384078 208412
rect 384146 208356 384202 208412
rect 384270 208356 384326 208412
rect 384394 208356 384450 208412
rect 384518 208356 384574 208412
rect 384642 208356 384698 208412
rect 384766 208356 384822 208412
rect 384890 208356 384946 208412
rect 385014 208356 385070 208412
rect 385138 208356 385194 208412
rect 384022 208232 384078 208288
rect 384146 208232 384202 208288
rect 384270 208232 384326 208288
rect 384394 208232 384450 208288
rect 384518 208232 384574 208288
rect 384642 208232 384698 208288
rect 384766 208232 384822 208288
rect 384890 208232 384946 208288
rect 385014 208232 385070 208288
rect 385138 208232 385194 208288
rect 384022 208108 384078 208164
rect 384146 208108 384202 208164
rect 384270 208108 384326 208164
rect 384394 208108 384450 208164
rect 384518 208108 384574 208164
rect 384642 208108 384698 208164
rect 384766 208108 384822 208164
rect 384890 208108 384946 208164
rect 385014 208108 385070 208164
rect 385138 208108 385194 208164
rect 384022 207984 384078 208040
rect 384146 207984 384202 208040
rect 384270 207984 384326 208040
rect 384394 207984 384450 208040
rect 384518 207984 384574 208040
rect 384642 207984 384698 208040
rect 384766 207984 384822 208040
rect 384890 207984 384946 208040
rect 385014 207984 385070 208040
rect 385138 207984 385194 208040
rect 384022 207860 384078 207916
rect 384146 207860 384202 207916
rect 384270 207860 384326 207916
rect 384394 207860 384450 207916
rect 384518 207860 384574 207916
rect 384642 207860 384698 207916
rect 384766 207860 384822 207916
rect 384890 207860 384946 207916
rect 385014 207860 385070 207916
rect 385138 207860 385194 207916
rect 404022 208356 404078 208412
rect 404146 208356 404202 208412
rect 404270 208356 404326 208412
rect 404394 208356 404450 208412
rect 404518 208356 404574 208412
rect 404642 208356 404698 208412
rect 404766 208356 404822 208412
rect 404890 208356 404946 208412
rect 405014 208356 405070 208412
rect 405138 208356 405194 208412
rect 404022 208232 404078 208288
rect 404146 208232 404202 208288
rect 404270 208232 404326 208288
rect 404394 208232 404450 208288
rect 404518 208232 404574 208288
rect 404642 208232 404698 208288
rect 404766 208232 404822 208288
rect 404890 208232 404946 208288
rect 405014 208232 405070 208288
rect 405138 208232 405194 208288
rect 404022 208108 404078 208164
rect 404146 208108 404202 208164
rect 404270 208108 404326 208164
rect 404394 208108 404450 208164
rect 404518 208108 404574 208164
rect 404642 208108 404698 208164
rect 404766 208108 404822 208164
rect 404890 208108 404946 208164
rect 405014 208108 405070 208164
rect 405138 208108 405194 208164
rect 404022 207984 404078 208040
rect 404146 207984 404202 208040
rect 404270 207984 404326 208040
rect 404394 207984 404450 208040
rect 404518 207984 404574 208040
rect 404642 207984 404698 208040
rect 404766 207984 404822 208040
rect 404890 207984 404946 208040
rect 405014 207984 405070 208040
rect 405138 207984 405194 208040
rect 404022 207860 404078 207916
rect 404146 207860 404202 207916
rect 404270 207860 404326 207916
rect 404394 207860 404450 207916
rect 404518 207860 404574 207916
rect 404642 207860 404698 207916
rect 404766 207860 404822 207916
rect 404890 207860 404946 207916
rect 405014 207860 405070 207916
rect 405138 207860 405194 207916
rect 424022 208356 424078 208412
rect 424146 208356 424202 208412
rect 424270 208356 424326 208412
rect 424394 208356 424450 208412
rect 424518 208356 424574 208412
rect 424642 208356 424698 208412
rect 424766 208356 424822 208412
rect 424890 208356 424946 208412
rect 425014 208356 425070 208412
rect 425138 208356 425194 208412
rect 424022 208232 424078 208288
rect 424146 208232 424202 208288
rect 424270 208232 424326 208288
rect 424394 208232 424450 208288
rect 424518 208232 424574 208288
rect 424642 208232 424698 208288
rect 424766 208232 424822 208288
rect 424890 208232 424946 208288
rect 425014 208232 425070 208288
rect 425138 208232 425194 208288
rect 424022 208108 424078 208164
rect 424146 208108 424202 208164
rect 424270 208108 424326 208164
rect 424394 208108 424450 208164
rect 424518 208108 424574 208164
rect 424642 208108 424698 208164
rect 424766 208108 424822 208164
rect 424890 208108 424946 208164
rect 425014 208108 425070 208164
rect 425138 208108 425194 208164
rect 424022 207984 424078 208040
rect 424146 207984 424202 208040
rect 424270 207984 424326 208040
rect 424394 207984 424450 208040
rect 424518 207984 424574 208040
rect 424642 207984 424698 208040
rect 424766 207984 424822 208040
rect 424890 207984 424946 208040
rect 425014 207984 425070 208040
rect 425138 207984 425194 208040
rect 424022 207860 424078 207916
rect 424146 207860 424202 207916
rect 424270 207860 424326 207916
rect 424394 207860 424450 207916
rect 424518 207860 424574 207916
rect 424642 207860 424698 207916
rect 424766 207860 424822 207916
rect 424890 207860 424946 207916
rect 425014 207860 425070 207916
rect 425138 207860 425194 207916
rect 444022 208356 444078 208412
rect 444146 208356 444202 208412
rect 444270 208356 444326 208412
rect 444394 208356 444450 208412
rect 444518 208356 444574 208412
rect 444642 208356 444698 208412
rect 444766 208356 444822 208412
rect 444890 208356 444946 208412
rect 445014 208356 445070 208412
rect 445138 208356 445194 208412
rect 444022 208232 444078 208288
rect 444146 208232 444202 208288
rect 444270 208232 444326 208288
rect 444394 208232 444450 208288
rect 444518 208232 444574 208288
rect 444642 208232 444698 208288
rect 444766 208232 444822 208288
rect 444890 208232 444946 208288
rect 445014 208232 445070 208288
rect 445138 208232 445194 208288
rect 444022 208108 444078 208164
rect 444146 208108 444202 208164
rect 444270 208108 444326 208164
rect 444394 208108 444450 208164
rect 444518 208108 444574 208164
rect 444642 208108 444698 208164
rect 444766 208108 444822 208164
rect 444890 208108 444946 208164
rect 445014 208108 445070 208164
rect 445138 208108 445194 208164
rect 444022 207984 444078 208040
rect 444146 207984 444202 208040
rect 444270 207984 444326 208040
rect 444394 207984 444450 208040
rect 444518 207984 444574 208040
rect 444642 207984 444698 208040
rect 444766 207984 444822 208040
rect 444890 207984 444946 208040
rect 445014 207984 445070 208040
rect 445138 207984 445194 208040
rect 444022 207860 444078 207916
rect 444146 207860 444202 207916
rect 444270 207860 444326 207916
rect 444394 207860 444450 207916
rect 444518 207860 444574 207916
rect 444642 207860 444698 207916
rect 444766 207860 444822 207916
rect 444890 207860 444946 207916
rect 445014 207860 445070 207916
rect 445138 207860 445194 207916
rect 464022 208356 464078 208412
rect 464146 208356 464202 208412
rect 464270 208356 464326 208412
rect 464394 208356 464450 208412
rect 464518 208356 464574 208412
rect 464642 208356 464698 208412
rect 464766 208356 464822 208412
rect 464890 208356 464946 208412
rect 465014 208356 465070 208412
rect 465138 208356 465194 208412
rect 464022 208232 464078 208288
rect 464146 208232 464202 208288
rect 464270 208232 464326 208288
rect 464394 208232 464450 208288
rect 464518 208232 464574 208288
rect 464642 208232 464698 208288
rect 464766 208232 464822 208288
rect 464890 208232 464946 208288
rect 465014 208232 465070 208288
rect 465138 208232 465194 208288
rect 464022 208108 464078 208164
rect 464146 208108 464202 208164
rect 464270 208108 464326 208164
rect 464394 208108 464450 208164
rect 464518 208108 464574 208164
rect 464642 208108 464698 208164
rect 464766 208108 464822 208164
rect 464890 208108 464946 208164
rect 465014 208108 465070 208164
rect 465138 208108 465194 208164
rect 464022 207984 464078 208040
rect 464146 207984 464202 208040
rect 464270 207984 464326 208040
rect 464394 207984 464450 208040
rect 464518 207984 464574 208040
rect 464642 207984 464698 208040
rect 464766 207984 464822 208040
rect 464890 207984 464946 208040
rect 465014 207984 465070 208040
rect 465138 207984 465194 208040
rect 464022 207860 464078 207916
rect 464146 207860 464202 207916
rect 464270 207860 464326 207916
rect 464394 207860 464450 207916
rect 464518 207860 464574 207916
rect 464642 207860 464698 207916
rect 464766 207860 464822 207916
rect 464890 207860 464946 207916
rect 465014 207860 465070 207916
rect 465138 207860 465194 207916
rect 484022 208356 484078 208412
rect 484146 208356 484202 208412
rect 484270 208356 484326 208412
rect 484394 208356 484450 208412
rect 484518 208356 484574 208412
rect 484642 208356 484698 208412
rect 484766 208356 484822 208412
rect 484890 208356 484946 208412
rect 485014 208356 485070 208412
rect 485138 208356 485194 208412
rect 484022 208232 484078 208288
rect 484146 208232 484202 208288
rect 484270 208232 484326 208288
rect 484394 208232 484450 208288
rect 484518 208232 484574 208288
rect 484642 208232 484698 208288
rect 484766 208232 484822 208288
rect 484890 208232 484946 208288
rect 485014 208232 485070 208288
rect 485138 208232 485194 208288
rect 484022 208108 484078 208164
rect 484146 208108 484202 208164
rect 484270 208108 484326 208164
rect 484394 208108 484450 208164
rect 484518 208108 484574 208164
rect 484642 208108 484698 208164
rect 484766 208108 484822 208164
rect 484890 208108 484946 208164
rect 485014 208108 485070 208164
rect 485138 208108 485194 208164
rect 484022 207984 484078 208040
rect 484146 207984 484202 208040
rect 484270 207984 484326 208040
rect 484394 207984 484450 208040
rect 484518 207984 484574 208040
rect 484642 207984 484698 208040
rect 484766 207984 484822 208040
rect 484890 207984 484946 208040
rect 485014 207984 485070 208040
rect 485138 207984 485194 208040
rect 484022 207860 484078 207916
rect 484146 207860 484202 207916
rect 484270 207860 484326 207916
rect 484394 207860 484450 207916
rect 484518 207860 484574 207916
rect 484642 207860 484698 207916
rect 484766 207860 484822 207916
rect 484890 207860 484946 207916
rect 485014 207860 485070 207916
rect 485138 207860 485194 207916
rect 504022 208356 504078 208412
rect 504146 208356 504202 208412
rect 504270 208356 504326 208412
rect 504394 208356 504450 208412
rect 504518 208356 504574 208412
rect 504642 208356 504698 208412
rect 504766 208356 504822 208412
rect 504890 208356 504946 208412
rect 505014 208356 505070 208412
rect 505138 208356 505194 208412
rect 504022 208232 504078 208288
rect 504146 208232 504202 208288
rect 504270 208232 504326 208288
rect 504394 208232 504450 208288
rect 504518 208232 504574 208288
rect 504642 208232 504698 208288
rect 504766 208232 504822 208288
rect 504890 208232 504946 208288
rect 505014 208232 505070 208288
rect 505138 208232 505194 208288
rect 504022 208108 504078 208164
rect 504146 208108 504202 208164
rect 504270 208108 504326 208164
rect 504394 208108 504450 208164
rect 504518 208108 504574 208164
rect 504642 208108 504698 208164
rect 504766 208108 504822 208164
rect 504890 208108 504946 208164
rect 505014 208108 505070 208164
rect 505138 208108 505194 208164
rect 504022 207984 504078 208040
rect 504146 207984 504202 208040
rect 504270 207984 504326 208040
rect 504394 207984 504450 208040
rect 504518 207984 504574 208040
rect 504642 207984 504698 208040
rect 504766 207984 504822 208040
rect 504890 207984 504946 208040
rect 505014 207984 505070 208040
rect 505138 207984 505194 208040
rect 504022 207860 504078 207916
rect 504146 207860 504202 207916
rect 504270 207860 504326 207916
rect 504394 207860 504450 207916
rect 504518 207860 504574 207916
rect 504642 207860 504698 207916
rect 504766 207860 504822 207916
rect 504890 207860 504946 207916
rect 505014 207860 505070 207916
rect 505138 207860 505194 207916
rect 524022 208356 524078 208412
rect 524146 208356 524202 208412
rect 524270 208356 524326 208412
rect 524394 208356 524450 208412
rect 524518 208356 524574 208412
rect 524642 208356 524698 208412
rect 524766 208356 524822 208412
rect 524890 208356 524946 208412
rect 525014 208356 525070 208412
rect 525138 208356 525194 208412
rect 524022 208232 524078 208288
rect 524146 208232 524202 208288
rect 524270 208232 524326 208288
rect 524394 208232 524450 208288
rect 524518 208232 524574 208288
rect 524642 208232 524698 208288
rect 524766 208232 524822 208288
rect 524890 208232 524946 208288
rect 525014 208232 525070 208288
rect 525138 208232 525194 208288
rect 524022 208108 524078 208164
rect 524146 208108 524202 208164
rect 524270 208108 524326 208164
rect 524394 208108 524450 208164
rect 524518 208108 524574 208164
rect 524642 208108 524698 208164
rect 524766 208108 524822 208164
rect 524890 208108 524946 208164
rect 525014 208108 525070 208164
rect 525138 208108 525194 208164
rect 524022 207984 524078 208040
rect 524146 207984 524202 208040
rect 524270 207984 524326 208040
rect 524394 207984 524450 208040
rect 524518 207984 524574 208040
rect 524642 207984 524698 208040
rect 524766 207984 524822 208040
rect 524890 207984 524946 208040
rect 525014 207984 525070 208040
rect 525138 207984 525194 208040
rect 524022 207860 524078 207916
rect 524146 207860 524202 207916
rect 524270 207860 524326 207916
rect 524394 207860 524450 207916
rect 524518 207860 524574 207916
rect 524642 207860 524698 207916
rect 524766 207860 524822 207916
rect 524890 207860 524946 207916
rect 525014 207860 525070 207916
rect 525138 207860 525194 207916
rect 544022 208356 544078 208412
rect 544146 208356 544202 208412
rect 544270 208356 544326 208412
rect 544394 208356 544450 208412
rect 544518 208356 544574 208412
rect 544642 208356 544698 208412
rect 544766 208356 544822 208412
rect 544890 208356 544946 208412
rect 545014 208356 545070 208412
rect 545138 208356 545194 208412
rect 544022 208232 544078 208288
rect 544146 208232 544202 208288
rect 544270 208232 544326 208288
rect 544394 208232 544450 208288
rect 544518 208232 544574 208288
rect 544642 208232 544698 208288
rect 544766 208232 544822 208288
rect 544890 208232 544946 208288
rect 545014 208232 545070 208288
rect 545138 208232 545194 208288
rect 544022 208108 544078 208164
rect 544146 208108 544202 208164
rect 544270 208108 544326 208164
rect 544394 208108 544450 208164
rect 544518 208108 544574 208164
rect 544642 208108 544698 208164
rect 544766 208108 544822 208164
rect 544890 208108 544946 208164
rect 545014 208108 545070 208164
rect 545138 208108 545194 208164
rect 544022 207984 544078 208040
rect 544146 207984 544202 208040
rect 544270 207984 544326 208040
rect 544394 207984 544450 208040
rect 544518 207984 544574 208040
rect 544642 207984 544698 208040
rect 544766 207984 544822 208040
rect 544890 207984 544946 208040
rect 545014 207984 545070 208040
rect 545138 207984 545194 208040
rect 544022 207860 544078 207916
rect 544146 207860 544202 207916
rect 544270 207860 544326 207916
rect 544394 207860 544450 207916
rect 544518 207860 544574 207916
rect 544642 207860 544698 207916
rect 544766 207860 544822 207916
rect 544890 207860 544946 207916
rect 545014 207860 545070 207916
rect 545138 207860 545194 207916
rect 354022 202356 354078 202412
rect 354146 202356 354202 202412
rect 354270 202356 354326 202412
rect 354394 202356 354450 202412
rect 354518 202356 354574 202412
rect 354642 202356 354698 202412
rect 354766 202356 354822 202412
rect 354890 202356 354946 202412
rect 355014 202356 355070 202412
rect 355138 202356 355194 202412
rect 354022 202232 354078 202288
rect 354146 202232 354202 202288
rect 354270 202232 354326 202288
rect 354394 202232 354450 202288
rect 354518 202232 354574 202288
rect 354642 202232 354698 202288
rect 354766 202232 354822 202288
rect 354890 202232 354946 202288
rect 355014 202232 355070 202288
rect 355138 202232 355194 202288
rect 354022 202108 354078 202164
rect 354146 202108 354202 202164
rect 354270 202108 354326 202164
rect 354394 202108 354450 202164
rect 354518 202108 354574 202164
rect 354642 202108 354698 202164
rect 354766 202108 354822 202164
rect 354890 202108 354946 202164
rect 355014 202108 355070 202164
rect 355138 202108 355194 202164
rect 354022 201984 354078 202040
rect 354146 201984 354202 202040
rect 354270 201984 354326 202040
rect 354394 201984 354450 202040
rect 354518 201984 354574 202040
rect 354642 201984 354698 202040
rect 354766 201984 354822 202040
rect 354890 201984 354946 202040
rect 355014 201984 355070 202040
rect 355138 201984 355194 202040
rect 354022 201860 354078 201916
rect 354146 201860 354202 201916
rect 354270 201860 354326 201916
rect 354394 201860 354450 201916
rect 354518 201860 354574 201916
rect 354642 201860 354698 201916
rect 354766 201860 354822 201916
rect 354890 201860 354946 201916
rect 355014 201860 355070 201916
rect 355138 201860 355194 201916
rect 374022 202356 374078 202412
rect 374146 202356 374202 202412
rect 374270 202356 374326 202412
rect 374394 202356 374450 202412
rect 374518 202356 374574 202412
rect 374642 202356 374698 202412
rect 374766 202356 374822 202412
rect 374890 202356 374946 202412
rect 375014 202356 375070 202412
rect 375138 202356 375194 202412
rect 374022 202232 374078 202288
rect 374146 202232 374202 202288
rect 374270 202232 374326 202288
rect 374394 202232 374450 202288
rect 374518 202232 374574 202288
rect 374642 202232 374698 202288
rect 374766 202232 374822 202288
rect 374890 202232 374946 202288
rect 375014 202232 375070 202288
rect 375138 202232 375194 202288
rect 374022 202108 374078 202164
rect 374146 202108 374202 202164
rect 374270 202108 374326 202164
rect 374394 202108 374450 202164
rect 374518 202108 374574 202164
rect 374642 202108 374698 202164
rect 374766 202108 374822 202164
rect 374890 202108 374946 202164
rect 375014 202108 375070 202164
rect 375138 202108 375194 202164
rect 374022 201984 374078 202040
rect 374146 201984 374202 202040
rect 374270 201984 374326 202040
rect 374394 201984 374450 202040
rect 374518 201984 374574 202040
rect 374642 201984 374698 202040
rect 374766 201984 374822 202040
rect 374890 201984 374946 202040
rect 375014 201984 375070 202040
rect 375138 201984 375194 202040
rect 374022 201860 374078 201916
rect 374146 201860 374202 201916
rect 374270 201860 374326 201916
rect 374394 201860 374450 201916
rect 374518 201860 374574 201916
rect 374642 201860 374698 201916
rect 374766 201860 374822 201916
rect 374890 201860 374946 201916
rect 375014 201860 375070 201916
rect 375138 201860 375194 201916
rect 394022 202356 394078 202412
rect 394146 202356 394202 202412
rect 394270 202356 394326 202412
rect 394394 202356 394450 202412
rect 394518 202356 394574 202412
rect 394642 202356 394698 202412
rect 394766 202356 394822 202412
rect 394890 202356 394946 202412
rect 395014 202356 395070 202412
rect 395138 202356 395194 202412
rect 394022 202232 394078 202288
rect 394146 202232 394202 202288
rect 394270 202232 394326 202288
rect 394394 202232 394450 202288
rect 394518 202232 394574 202288
rect 394642 202232 394698 202288
rect 394766 202232 394822 202288
rect 394890 202232 394946 202288
rect 395014 202232 395070 202288
rect 395138 202232 395194 202288
rect 394022 202108 394078 202164
rect 394146 202108 394202 202164
rect 394270 202108 394326 202164
rect 394394 202108 394450 202164
rect 394518 202108 394574 202164
rect 394642 202108 394698 202164
rect 394766 202108 394822 202164
rect 394890 202108 394946 202164
rect 395014 202108 395070 202164
rect 395138 202108 395194 202164
rect 394022 201984 394078 202040
rect 394146 201984 394202 202040
rect 394270 201984 394326 202040
rect 394394 201984 394450 202040
rect 394518 201984 394574 202040
rect 394642 201984 394698 202040
rect 394766 201984 394822 202040
rect 394890 201984 394946 202040
rect 395014 201984 395070 202040
rect 395138 201984 395194 202040
rect 394022 201860 394078 201916
rect 394146 201860 394202 201916
rect 394270 201860 394326 201916
rect 394394 201860 394450 201916
rect 394518 201860 394574 201916
rect 394642 201860 394698 201916
rect 394766 201860 394822 201916
rect 394890 201860 394946 201916
rect 395014 201860 395070 201916
rect 395138 201860 395194 201916
rect 414022 202356 414078 202412
rect 414146 202356 414202 202412
rect 414270 202356 414326 202412
rect 414394 202356 414450 202412
rect 414518 202356 414574 202412
rect 414642 202356 414698 202412
rect 414766 202356 414822 202412
rect 414890 202356 414946 202412
rect 415014 202356 415070 202412
rect 415138 202356 415194 202412
rect 414022 202232 414078 202288
rect 414146 202232 414202 202288
rect 414270 202232 414326 202288
rect 414394 202232 414450 202288
rect 414518 202232 414574 202288
rect 414642 202232 414698 202288
rect 414766 202232 414822 202288
rect 414890 202232 414946 202288
rect 415014 202232 415070 202288
rect 415138 202232 415194 202288
rect 414022 202108 414078 202164
rect 414146 202108 414202 202164
rect 414270 202108 414326 202164
rect 414394 202108 414450 202164
rect 414518 202108 414574 202164
rect 414642 202108 414698 202164
rect 414766 202108 414822 202164
rect 414890 202108 414946 202164
rect 415014 202108 415070 202164
rect 415138 202108 415194 202164
rect 414022 201984 414078 202040
rect 414146 201984 414202 202040
rect 414270 201984 414326 202040
rect 414394 201984 414450 202040
rect 414518 201984 414574 202040
rect 414642 201984 414698 202040
rect 414766 201984 414822 202040
rect 414890 201984 414946 202040
rect 415014 201984 415070 202040
rect 415138 201984 415194 202040
rect 414022 201860 414078 201916
rect 414146 201860 414202 201916
rect 414270 201860 414326 201916
rect 414394 201860 414450 201916
rect 414518 201860 414574 201916
rect 414642 201860 414698 201916
rect 414766 201860 414822 201916
rect 414890 201860 414946 201916
rect 415014 201860 415070 201916
rect 415138 201860 415194 201916
rect 434022 202356 434078 202412
rect 434146 202356 434202 202412
rect 434270 202356 434326 202412
rect 434394 202356 434450 202412
rect 434518 202356 434574 202412
rect 434642 202356 434698 202412
rect 434766 202356 434822 202412
rect 434890 202356 434946 202412
rect 435014 202356 435070 202412
rect 435138 202356 435194 202412
rect 434022 202232 434078 202288
rect 434146 202232 434202 202288
rect 434270 202232 434326 202288
rect 434394 202232 434450 202288
rect 434518 202232 434574 202288
rect 434642 202232 434698 202288
rect 434766 202232 434822 202288
rect 434890 202232 434946 202288
rect 435014 202232 435070 202288
rect 435138 202232 435194 202288
rect 434022 202108 434078 202164
rect 434146 202108 434202 202164
rect 434270 202108 434326 202164
rect 434394 202108 434450 202164
rect 434518 202108 434574 202164
rect 434642 202108 434698 202164
rect 434766 202108 434822 202164
rect 434890 202108 434946 202164
rect 435014 202108 435070 202164
rect 435138 202108 435194 202164
rect 434022 201984 434078 202040
rect 434146 201984 434202 202040
rect 434270 201984 434326 202040
rect 434394 201984 434450 202040
rect 434518 201984 434574 202040
rect 434642 201984 434698 202040
rect 434766 201984 434822 202040
rect 434890 201984 434946 202040
rect 435014 201984 435070 202040
rect 435138 201984 435194 202040
rect 434022 201860 434078 201916
rect 434146 201860 434202 201916
rect 434270 201860 434326 201916
rect 434394 201860 434450 201916
rect 434518 201860 434574 201916
rect 434642 201860 434698 201916
rect 434766 201860 434822 201916
rect 434890 201860 434946 201916
rect 435014 201860 435070 201916
rect 435138 201860 435194 201916
rect 454022 202356 454078 202412
rect 454146 202356 454202 202412
rect 454270 202356 454326 202412
rect 454394 202356 454450 202412
rect 454518 202356 454574 202412
rect 454642 202356 454698 202412
rect 454766 202356 454822 202412
rect 454890 202356 454946 202412
rect 455014 202356 455070 202412
rect 455138 202356 455194 202412
rect 454022 202232 454078 202288
rect 454146 202232 454202 202288
rect 454270 202232 454326 202288
rect 454394 202232 454450 202288
rect 454518 202232 454574 202288
rect 454642 202232 454698 202288
rect 454766 202232 454822 202288
rect 454890 202232 454946 202288
rect 455014 202232 455070 202288
rect 455138 202232 455194 202288
rect 454022 202108 454078 202164
rect 454146 202108 454202 202164
rect 454270 202108 454326 202164
rect 454394 202108 454450 202164
rect 454518 202108 454574 202164
rect 454642 202108 454698 202164
rect 454766 202108 454822 202164
rect 454890 202108 454946 202164
rect 455014 202108 455070 202164
rect 455138 202108 455194 202164
rect 454022 201984 454078 202040
rect 454146 201984 454202 202040
rect 454270 201984 454326 202040
rect 454394 201984 454450 202040
rect 454518 201984 454574 202040
rect 454642 201984 454698 202040
rect 454766 201984 454822 202040
rect 454890 201984 454946 202040
rect 455014 201984 455070 202040
rect 455138 201984 455194 202040
rect 454022 201860 454078 201916
rect 454146 201860 454202 201916
rect 454270 201860 454326 201916
rect 454394 201860 454450 201916
rect 454518 201860 454574 201916
rect 454642 201860 454698 201916
rect 454766 201860 454822 201916
rect 454890 201860 454946 201916
rect 455014 201860 455070 201916
rect 455138 201860 455194 201916
rect 474022 202356 474078 202412
rect 474146 202356 474202 202412
rect 474270 202356 474326 202412
rect 474394 202356 474450 202412
rect 474518 202356 474574 202412
rect 474642 202356 474698 202412
rect 474766 202356 474822 202412
rect 474890 202356 474946 202412
rect 475014 202356 475070 202412
rect 475138 202356 475194 202412
rect 474022 202232 474078 202288
rect 474146 202232 474202 202288
rect 474270 202232 474326 202288
rect 474394 202232 474450 202288
rect 474518 202232 474574 202288
rect 474642 202232 474698 202288
rect 474766 202232 474822 202288
rect 474890 202232 474946 202288
rect 475014 202232 475070 202288
rect 475138 202232 475194 202288
rect 474022 202108 474078 202164
rect 474146 202108 474202 202164
rect 474270 202108 474326 202164
rect 474394 202108 474450 202164
rect 474518 202108 474574 202164
rect 474642 202108 474698 202164
rect 474766 202108 474822 202164
rect 474890 202108 474946 202164
rect 475014 202108 475070 202164
rect 475138 202108 475194 202164
rect 474022 201984 474078 202040
rect 474146 201984 474202 202040
rect 474270 201984 474326 202040
rect 474394 201984 474450 202040
rect 474518 201984 474574 202040
rect 474642 201984 474698 202040
rect 474766 201984 474822 202040
rect 474890 201984 474946 202040
rect 475014 201984 475070 202040
rect 475138 201984 475194 202040
rect 474022 201860 474078 201916
rect 474146 201860 474202 201916
rect 474270 201860 474326 201916
rect 474394 201860 474450 201916
rect 474518 201860 474574 201916
rect 474642 201860 474698 201916
rect 474766 201860 474822 201916
rect 474890 201860 474946 201916
rect 475014 201860 475070 201916
rect 475138 201860 475194 201916
rect 494022 202356 494078 202412
rect 494146 202356 494202 202412
rect 494270 202356 494326 202412
rect 494394 202356 494450 202412
rect 494518 202356 494574 202412
rect 494642 202356 494698 202412
rect 494766 202356 494822 202412
rect 494890 202356 494946 202412
rect 495014 202356 495070 202412
rect 495138 202356 495194 202412
rect 494022 202232 494078 202288
rect 494146 202232 494202 202288
rect 494270 202232 494326 202288
rect 494394 202232 494450 202288
rect 494518 202232 494574 202288
rect 494642 202232 494698 202288
rect 494766 202232 494822 202288
rect 494890 202232 494946 202288
rect 495014 202232 495070 202288
rect 495138 202232 495194 202288
rect 494022 202108 494078 202164
rect 494146 202108 494202 202164
rect 494270 202108 494326 202164
rect 494394 202108 494450 202164
rect 494518 202108 494574 202164
rect 494642 202108 494698 202164
rect 494766 202108 494822 202164
rect 494890 202108 494946 202164
rect 495014 202108 495070 202164
rect 495138 202108 495194 202164
rect 494022 201984 494078 202040
rect 494146 201984 494202 202040
rect 494270 201984 494326 202040
rect 494394 201984 494450 202040
rect 494518 201984 494574 202040
rect 494642 201984 494698 202040
rect 494766 201984 494822 202040
rect 494890 201984 494946 202040
rect 495014 201984 495070 202040
rect 495138 201984 495194 202040
rect 494022 201860 494078 201916
rect 494146 201860 494202 201916
rect 494270 201860 494326 201916
rect 494394 201860 494450 201916
rect 494518 201860 494574 201916
rect 494642 201860 494698 201916
rect 494766 201860 494822 201916
rect 494890 201860 494946 201916
rect 495014 201860 495070 201916
rect 495138 201860 495194 201916
rect 514022 202356 514078 202412
rect 514146 202356 514202 202412
rect 514270 202356 514326 202412
rect 514394 202356 514450 202412
rect 514518 202356 514574 202412
rect 514642 202356 514698 202412
rect 514766 202356 514822 202412
rect 514890 202356 514946 202412
rect 515014 202356 515070 202412
rect 515138 202356 515194 202412
rect 514022 202232 514078 202288
rect 514146 202232 514202 202288
rect 514270 202232 514326 202288
rect 514394 202232 514450 202288
rect 514518 202232 514574 202288
rect 514642 202232 514698 202288
rect 514766 202232 514822 202288
rect 514890 202232 514946 202288
rect 515014 202232 515070 202288
rect 515138 202232 515194 202288
rect 514022 202108 514078 202164
rect 514146 202108 514202 202164
rect 514270 202108 514326 202164
rect 514394 202108 514450 202164
rect 514518 202108 514574 202164
rect 514642 202108 514698 202164
rect 514766 202108 514822 202164
rect 514890 202108 514946 202164
rect 515014 202108 515070 202164
rect 515138 202108 515194 202164
rect 514022 201984 514078 202040
rect 514146 201984 514202 202040
rect 514270 201984 514326 202040
rect 514394 201984 514450 202040
rect 514518 201984 514574 202040
rect 514642 201984 514698 202040
rect 514766 201984 514822 202040
rect 514890 201984 514946 202040
rect 515014 201984 515070 202040
rect 515138 201984 515194 202040
rect 514022 201860 514078 201916
rect 514146 201860 514202 201916
rect 514270 201860 514326 201916
rect 514394 201860 514450 201916
rect 514518 201860 514574 201916
rect 514642 201860 514698 201916
rect 514766 201860 514822 201916
rect 514890 201860 514946 201916
rect 515014 201860 515070 201916
rect 515138 201860 515194 201916
rect 534022 202356 534078 202412
rect 534146 202356 534202 202412
rect 534270 202356 534326 202412
rect 534394 202356 534450 202412
rect 534518 202356 534574 202412
rect 534642 202356 534698 202412
rect 534766 202356 534822 202412
rect 534890 202356 534946 202412
rect 535014 202356 535070 202412
rect 535138 202356 535194 202412
rect 534022 202232 534078 202288
rect 534146 202232 534202 202288
rect 534270 202232 534326 202288
rect 534394 202232 534450 202288
rect 534518 202232 534574 202288
rect 534642 202232 534698 202288
rect 534766 202232 534822 202288
rect 534890 202232 534946 202288
rect 535014 202232 535070 202288
rect 535138 202232 535194 202288
rect 534022 202108 534078 202164
rect 534146 202108 534202 202164
rect 534270 202108 534326 202164
rect 534394 202108 534450 202164
rect 534518 202108 534574 202164
rect 534642 202108 534698 202164
rect 534766 202108 534822 202164
rect 534890 202108 534946 202164
rect 535014 202108 535070 202164
rect 535138 202108 535194 202164
rect 534022 201984 534078 202040
rect 534146 201984 534202 202040
rect 534270 201984 534326 202040
rect 534394 201984 534450 202040
rect 534518 201984 534574 202040
rect 534642 201984 534698 202040
rect 534766 201984 534822 202040
rect 534890 201984 534946 202040
rect 535014 201984 535070 202040
rect 535138 201984 535194 202040
rect 534022 201860 534078 201916
rect 534146 201860 534202 201916
rect 534270 201860 534326 201916
rect 534394 201860 534450 201916
rect 534518 201860 534574 201916
rect 534642 201860 534698 201916
rect 534766 201860 534822 201916
rect 534890 201860 534946 201916
rect 535014 201860 535070 201916
rect 535138 201860 535194 201916
rect 348970 190294 349026 190350
rect 349094 190294 349150 190350
rect 349218 190294 349274 190350
rect 349342 190294 349398 190350
rect 348970 190170 349026 190226
rect 349094 190170 349150 190226
rect 349218 190170 349274 190226
rect 349342 190170 349398 190226
rect 348970 190046 349026 190102
rect 349094 190046 349150 190102
rect 349218 190046 349274 190102
rect 349342 190046 349398 190102
rect 348970 189922 349026 189978
rect 349094 189922 349150 189978
rect 349218 189922 349274 189978
rect 349342 189922 349398 189978
rect 345250 166294 345306 166350
rect 345374 166294 345430 166350
rect 345498 166294 345554 166350
rect 345622 166294 345678 166350
rect 345250 166170 345306 166226
rect 345374 166170 345430 166226
rect 345498 166170 345554 166226
rect 345622 166170 345678 166226
rect 345250 166046 345306 166102
rect 345374 166046 345430 166102
rect 345498 166046 345554 166102
rect 345622 166046 345678 166102
rect 345250 165922 345306 165978
rect 345374 165922 345430 165978
rect 345498 165922 345554 165978
rect 345622 165922 345678 165978
rect 345250 148294 345306 148350
rect 345374 148294 345430 148350
rect 345498 148294 345554 148350
rect 345622 148294 345678 148350
rect 345250 148170 345306 148226
rect 345374 148170 345430 148226
rect 345498 148170 345554 148226
rect 345622 148170 345678 148226
rect 345250 148046 345306 148102
rect 345374 148046 345430 148102
rect 345498 148046 345554 148102
rect 345622 148046 345678 148102
rect 345250 147922 345306 147978
rect 345374 147922 345430 147978
rect 345498 147922 345554 147978
rect 345622 147922 345678 147978
rect 345250 130294 345306 130350
rect 345374 130294 345430 130350
rect 345498 130294 345554 130350
rect 345622 130294 345678 130350
rect 345250 130170 345306 130226
rect 345374 130170 345430 130226
rect 345498 130170 345554 130226
rect 345622 130170 345678 130226
rect 345250 130046 345306 130102
rect 345374 130046 345430 130102
rect 345498 130046 345554 130102
rect 345622 130046 345678 130102
rect 345250 129922 345306 129978
rect 345374 129922 345430 129978
rect 345498 129922 345554 129978
rect 345622 129922 345678 129978
rect 345250 112294 345306 112350
rect 345374 112294 345430 112350
rect 345498 112294 345554 112350
rect 345622 112294 345678 112350
rect 345250 112170 345306 112226
rect 345374 112170 345430 112226
rect 345498 112170 345554 112226
rect 345622 112170 345678 112226
rect 345250 112046 345306 112102
rect 345374 112046 345430 112102
rect 345498 112046 345554 112102
rect 345622 112046 345678 112102
rect 345250 111922 345306 111978
rect 345374 111922 345430 111978
rect 345498 111922 345554 111978
rect 345622 111922 345678 111978
rect 345250 94294 345306 94350
rect 345374 94294 345430 94350
rect 345498 94294 345554 94350
rect 345622 94294 345678 94350
rect 345250 94170 345306 94226
rect 345374 94170 345430 94226
rect 345498 94170 345554 94226
rect 345622 94170 345678 94226
rect 345250 94046 345306 94102
rect 345374 94046 345430 94102
rect 345498 94046 345554 94102
rect 345622 94046 345678 94102
rect 345250 93922 345306 93978
rect 345374 93922 345430 93978
rect 345498 93922 345554 93978
rect 345622 93922 345678 93978
rect 345250 76294 345306 76350
rect 345374 76294 345430 76350
rect 345498 76294 345554 76350
rect 345622 76294 345678 76350
rect 345250 76170 345306 76226
rect 345374 76170 345430 76226
rect 345498 76170 345554 76226
rect 345622 76170 345678 76226
rect 345250 76046 345306 76102
rect 345374 76046 345430 76102
rect 345498 76046 345554 76102
rect 345622 76046 345678 76102
rect 345250 75922 345306 75978
rect 345374 75922 345430 75978
rect 345498 75922 345554 75978
rect 345622 75922 345678 75978
rect 345250 58294 345306 58350
rect 345374 58294 345430 58350
rect 345498 58294 345554 58350
rect 345622 58294 345678 58350
rect 345250 58170 345306 58226
rect 345374 58170 345430 58226
rect 345498 58170 345554 58226
rect 345622 58170 345678 58226
rect 345250 58046 345306 58102
rect 345374 58046 345430 58102
rect 345498 58046 345554 58102
rect 345622 58046 345678 58102
rect 345250 57922 345306 57978
rect 345374 57922 345430 57978
rect 345498 57922 345554 57978
rect 345622 57922 345678 57978
rect 330970 46294 331026 46350
rect 331094 46294 331150 46350
rect 331218 46294 331274 46350
rect 331342 46294 331398 46350
rect 330970 46170 331026 46226
rect 331094 46170 331150 46226
rect 331218 46170 331274 46226
rect 331342 46170 331398 46226
rect 330970 46046 331026 46102
rect 331094 46046 331150 46102
rect 331218 46046 331274 46102
rect 331342 46046 331398 46102
rect 330970 45922 331026 45978
rect 331094 45922 331150 45978
rect 331218 45922 331274 45978
rect 331342 45922 331398 45978
rect 345250 40294 345306 40350
rect 345374 40294 345430 40350
rect 345498 40294 345554 40350
rect 345622 40294 345678 40350
rect 345250 40170 345306 40226
rect 345374 40170 345430 40226
rect 345498 40170 345554 40226
rect 345622 40170 345678 40226
rect 345250 40046 345306 40102
rect 345374 40046 345430 40102
rect 345498 40046 345554 40102
rect 345622 40046 345678 40102
rect 345250 39922 345306 39978
rect 345374 39922 345430 39978
rect 345498 39922 345554 39978
rect 345622 39922 345678 39978
rect 330970 28294 331026 28350
rect 331094 28294 331150 28350
rect 331218 28294 331274 28350
rect 331342 28294 331398 28350
rect 330970 28170 331026 28226
rect 331094 28170 331150 28226
rect 331218 28170 331274 28226
rect 331342 28170 331398 28226
rect 330970 28046 331026 28102
rect 331094 28046 331150 28102
rect 331218 28046 331274 28102
rect 331342 28046 331398 28102
rect 330970 27922 331026 27978
rect 331094 27922 331150 27978
rect 331218 27922 331274 27978
rect 331342 27922 331398 27978
rect 330970 10294 331026 10350
rect 331094 10294 331150 10350
rect 331218 10294 331274 10350
rect 331342 10294 331398 10350
rect 330970 10170 331026 10226
rect 331094 10170 331150 10226
rect 331218 10170 331274 10226
rect 331342 10170 331398 10226
rect 330970 10046 331026 10102
rect 331094 10046 331150 10102
rect 331218 10046 331274 10102
rect 331342 10046 331398 10102
rect 330970 9922 331026 9978
rect 331094 9922 331150 9978
rect 331218 9922 331274 9978
rect 331342 9922 331398 9978
rect 330970 -1176 331026 -1120
rect 331094 -1176 331150 -1120
rect 331218 -1176 331274 -1120
rect 331342 -1176 331398 -1120
rect 330970 -1300 331026 -1244
rect 331094 -1300 331150 -1244
rect 331218 -1300 331274 -1244
rect 331342 -1300 331398 -1244
rect 330970 -1424 331026 -1368
rect 331094 -1424 331150 -1368
rect 331218 -1424 331274 -1368
rect 331342 -1424 331398 -1368
rect 330970 -1548 331026 -1492
rect 331094 -1548 331150 -1492
rect 331218 -1548 331274 -1492
rect 331342 -1548 331398 -1492
rect 346780 42722 346836 42778
rect 348970 172294 349026 172350
rect 349094 172294 349150 172350
rect 349218 172294 349274 172350
rect 349342 172294 349398 172350
rect 348970 172170 349026 172226
rect 349094 172170 349150 172226
rect 349218 172170 349274 172226
rect 349342 172170 349398 172226
rect 348970 172046 349026 172102
rect 349094 172046 349150 172102
rect 349218 172046 349274 172102
rect 349342 172046 349398 172102
rect 348970 171922 349026 171978
rect 349094 171922 349150 171978
rect 349218 171922 349274 171978
rect 349342 171922 349398 171978
rect 348970 154294 349026 154350
rect 349094 154294 349150 154350
rect 349218 154294 349274 154350
rect 349342 154294 349398 154350
rect 348970 154170 349026 154226
rect 349094 154170 349150 154226
rect 349218 154170 349274 154226
rect 349342 154170 349398 154226
rect 348970 154046 349026 154102
rect 349094 154046 349150 154102
rect 349218 154046 349274 154102
rect 349342 154046 349398 154102
rect 348970 153922 349026 153978
rect 349094 153922 349150 153978
rect 349218 153922 349274 153978
rect 349342 153922 349398 153978
rect 348970 136294 349026 136350
rect 349094 136294 349150 136350
rect 349218 136294 349274 136350
rect 349342 136294 349398 136350
rect 348970 136170 349026 136226
rect 349094 136170 349150 136226
rect 349218 136170 349274 136226
rect 349342 136170 349398 136226
rect 348970 136046 349026 136102
rect 349094 136046 349150 136102
rect 349218 136046 349274 136102
rect 349342 136046 349398 136102
rect 348970 135922 349026 135978
rect 349094 135922 349150 135978
rect 349218 135922 349274 135978
rect 349342 135922 349398 135978
rect 348970 118294 349026 118350
rect 349094 118294 349150 118350
rect 349218 118294 349274 118350
rect 349342 118294 349398 118350
rect 348970 118170 349026 118226
rect 349094 118170 349150 118226
rect 349218 118170 349274 118226
rect 349342 118170 349398 118226
rect 348970 118046 349026 118102
rect 349094 118046 349150 118102
rect 349218 118046 349274 118102
rect 349342 118046 349398 118102
rect 348970 117922 349026 117978
rect 349094 117922 349150 117978
rect 349218 117922 349274 117978
rect 349342 117922 349398 117978
rect 348970 100294 349026 100350
rect 349094 100294 349150 100350
rect 349218 100294 349274 100350
rect 349342 100294 349398 100350
rect 348970 100170 349026 100226
rect 349094 100170 349150 100226
rect 349218 100170 349274 100226
rect 349342 100170 349398 100226
rect 348970 100046 349026 100102
rect 349094 100046 349150 100102
rect 349218 100046 349274 100102
rect 349342 100046 349398 100102
rect 348970 99922 349026 99978
rect 349094 99922 349150 99978
rect 349218 99922 349274 99978
rect 349342 99922 349398 99978
rect 348970 82294 349026 82350
rect 349094 82294 349150 82350
rect 349218 82294 349274 82350
rect 349342 82294 349398 82350
rect 348970 82170 349026 82226
rect 349094 82170 349150 82226
rect 349218 82170 349274 82226
rect 349342 82170 349398 82226
rect 348970 82046 349026 82102
rect 349094 82046 349150 82102
rect 349218 82046 349274 82102
rect 349342 82046 349398 82102
rect 348970 81922 349026 81978
rect 349094 81922 349150 81978
rect 349218 81922 349274 81978
rect 349342 81922 349398 81978
rect 348970 64294 349026 64350
rect 349094 64294 349150 64350
rect 349218 64294 349274 64350
rect 349342 64294 349398 64350
rect 348970 64170 349026 64226
rect 349094 64170 349150 64226
rect 349218 64170 349274 64226
rect 349342 64170 349398 64226
rect 348970 64046 349026 64102
rect 349094 64046 349150 64102
rect 349218 64046 349274 64102
rect 349342 64046 349398 64102
rect 348970 63922 349026 63978
rect 349094 63922 349150 63978
rect 349218 63922 349274 63978
rect 349342 63922 349398 63978
rect 548940 59822 548996 59878
rect 348970 46294 349026 46350
rect 349094 46294 349150 46350
rect 349218 46294 349274 46350
rect 349342 46294 349398 46350
rect 348970 46170 349026 46226
rect 349094 46170 349150 46226
rect 349218 46170 349274 46226
rect 349342 46170 349398 46226
rect 348970 46046 349026 46102
rect 349094 46046 349150 46102
rect 349218 46046 349274 46102
rect 349342 46046 349398 46102
rect 348970 45922 349026 45978
rect 349094 45922 349150 45978
rect 349218 45922 349274 45978
rect 349342 45922 349398 45978
rect 348970 28294 349026 28350
rect 349094 28294 349150 28350
rect 349218 28294 349274 28350
rect 349342 28294 349398 28350
rect 348970 28170 349026 28226
rect 349094 28170 349150 28226
rect 349218 28170 349274 28226
rect 349342 28170 349398 28226
rect 348970 28046 349026 28102
rect 349094 28046 349150 28102
rect 349218 28046 349274 28102
rect 349342 28046 349398 28102
rect 348970 27922 349026 27978
rect 349094 27922 349150 27978
rect 349218 27922 349274 27978
rect 349342 27922 349398 27978
rect 345250 22294 345306 22350
rect 345374 22294 345430 22350
rect 345498 22294 345554 22350
rect 345622 22294 345678 22350
rect 345250 22170 345306 22226
rect 345374 22170 345430 22226
rect 345498 22170 345554 22226
rect 345622 22170 345678 22226
rect 345250 22046 345306 22102
rect 345374 22046 345430 22102
rect 345498 22046 345554 22102
rect 345622 22046 345678 22102
rect 345250 21922 345306 21978
rect 345374 21922 345430 21978
rect 345498 21922 345554 21978
rect 345622 21922 345678 21978
rect 345250 4294 345306 4350
rect 345374 4294 345430 4350
rect 345498 4294 345554 4350
rect 345622 4294 345678 4350
rect 345250 4170 345306 4226
rect 345374 4170 345430 4226
rect 345498 4170 345554 4226
rect 345622 4170 345678 4226
rect 345250 4046 345306 4102
rect 345374 4046 345430 4102
rect 345498 4046 345554 4102
rect 345622 4046 345678 4102
rect 345250 3922 345306 3978
rect 345374 3922 345430 3978
rect 345498 3922 345554 3978
rect 345622 3922 345678 3978
rect 345250 -216 345306 -160
rect 345374 -216 345430 -160
rect 345498 -216 345554 -160
rect 345622 -216 345678 -160
rect 345250 -340 345306 -284
rect 345374 -340 345430 -284
rect 345498 -340 345554 -284
rect 345622 -340 345678 -284
rect 345250 -464 345306 -408
rect 345374 -464 345430 -408
rect 345498 -464 345554 -408
rect 345622 -464 345678 -408
rect 345250 -588 345306 -532
rect 345374 -588 345430 -532
rect 345498 -588 345554 -532
rect 345622 -588 345678 -532
rect 548716 54602 548772 54658
rect 350252 25082 350308 25138
rect 525308 43082 525364 43138
rect 516460 42902 516516 42958
rect 436268 41282 436324 41338
rect 363250 40294 363306 40350
rect 363374 40294 363430 40350
rect 363498 40294 363554 40350
rect 363622 40294 363678 40350
rect 363250 40170 363306 40226
rect 363374 40170 363430 40226
rect 363498 40170 363554 40226
rect 363622 40170 363678 40226
rect 363250 40046 363306 40102
rect 363374 40046 363430 40102
rect 363498 40046 363554 40102
rect 363622 40046 363678 40102
rect 363250 39922 363306 39978
rect 363374 39922 363430 39978
rect 363498 39922 363554 39978
rect 363622 39922 363678 39978
rect 354508 37716 354564 37738
rect 354508 37682 354564 37716
rect 362908 36988 362964 37018
rect 362908 36962 362964 36988
rect 363250 22294 363306 22350
rect 363374 22294 363430 22350
rect 363498 22294 363554 22350
rect 363622 22294 363678 22350
rect 363250 22170 363306 22226
rect 363374 22170 363430 22226
rect 363498 22170 363554 22226
rect 363622 22170 363678 22226
rect 363250 22046 363306 22102
rect 363374 22046 363430 22102
rect 363498 22046 363554 22102
rect 363622 22046 363678 22102
rect 363250 21922 363306 21978
rect 363374 21922 363430 21978
rect 363498 21922 363554 21978
rect 363622 21922 363678 21978
rect 348970 10294 349026 10350
rect 349094 10294 349150 10350
rect 349218 10294 349274 10350
rect 349342 10294 349398 10350
rect 348970 10170 349026 10226
rect 349094 10170 349150 10226
rect 349218 10170 349274 10226
rect 349342 10170 349398 10226
rect 348970 10046 349026 10102
rect 349094 10046 349150 10102
rect 349218 10046 349274 10102
rect 349342 10046 349398 10102
rect 348970 9922 349026 9978
rect 349094 9922 349150 9978
rect 349218 9922 349274 9978
rect 349342 9922 349398 9978
rect 348970 -1176 349026 -1120
rect 349094 -1176 349150 -1120
rect 349218 -1176 349274 -1120
rect 349342 -1176 349398 -1120
rect 348970 -1300 349026 -1244
rect 349094 -1300 349150 -1244
rect 349218 -1300 349274 -1244
rect 349342 -1300 349398 -1244
rect 348970 -1424 349026 -1368
rect 349094 -1424 349150 -1368
rect 349218 -1424 349274 -1368
rect 349342 -1424 349398 -1368
rect 348970 -1548 349026 -1492
rect 349094 -1548 349150 -1492
rect 349218 -1548 349274 -1492
rect 349342 -1548 349398 -1492
rect 363250 4294 363306 4350
rect 363374 4294 363430 4350
rect 363498 4294 363554 4350
rect 363622 4294 363678 4350
rect 363250 4170 363306 4226
rect 363374 4170 363430 4226
rect 363498 4170 363554 4226
rect 363622 4170 363678 4226
rect 363250 4046 363306 4102
rect 363374 4046 363430 4102
rect 363498 4046 363554 4102
rect 363622 4046 363678 4102
rect 363250 3922 363306 3978
rect 363374 3922 363430 3978
rect 363498 3922 363554 3978
rect 363622 3922 363678 3978
rect 363250 -216 363306 -160
rect 363374 -216 363430 -160
rect 363498 -216 363554 -160
rect 363622 -216 363678 -160
rect 363250 -340 363306 -284
rect 363374 -340 363430 -284
rect 363498 -340 363554 -284
rect 363622 -340 363678 -284
rect 363250 -464 363306 -408
rect 363374 -464 363430 -408
rect 363498 -464 363554 -408
rect 363622 -464 363678 -408
rect 363250 -588 363306 -532
rect 363374 -588 363430 -532
rect 363498 -588 363554 -532
rect 363622 -588 363678 -532
rect 381250 40294 381306 40350
rect 381374 40294 381430 40350
rect 381498 40294 381554 40350
rect 381622 40294 381678 40350
rect 381250 40170 381306 40226
rect 381374 40170 381430 40226
rect 381498 40170 381554 40226
rect 381622 40170 381678 40226
rect 381250 40046 381306 40102
rect 381374 40046 381430 40102
rect 381498 40046 381554 40102
rect 381622 40046 381678 40102
rect 381250 39922 381306 39978
rect 381374 39922 381430 39978
rect 381498 39922 381554 39978
rect 381622 39922 381678 39978
rect 366970 28294 367026 28350
rect 367094 28294 367150 28350
rect 367218 28294 367274 28350
rect 367342 28294 367398 28350
rect 366970 28170 367026 28226
rect 367094 28170 367150 28226
rect 367218 28170 367274 28226
rect 367342 28170 367398 28226
rect 366970 28046 367026 28102
rect 367094 28046 367150 28102
rect 367218 28046 367274 28102
rect 367342 28046 367398 28102
rect 366970 27922 367026 27978
rect 367094 27922 367150 27978
rect 367218 27922 367274 27978
rect 367342 27922 367398 27978
rect 371308 24902 371364 24958
rect 366970 10294 367026 10350
rect 367094 10294 367150 10350
rect 367218 10294 367274 10350
rect 367342 10294 367398 10350
rect 366970 10170 367026 10226
rect 367094 10170 367150 10226
rect 367218 10170 367274 10226
rect 367342 10170 367398 10226
rect 366970 10046 367026 10102
rect 367094 10046 367150 10102
rect 367218 10046 367274 10102
rect 367342 10046 367398 10102
rect 366970 9922 367026 9978
rect 367094 9922 367150 9978
rect 367218 9922 367274 9978
rect 367342 9922 367398 9978
rect 366970 -1176 367026 -1120
rect 367094 -1176 367150 -1120
rect 367218 -1176 367274 -1120
rect 367342 -1176 367398 -1120
rect 366970 -1300 367026 -1244
rect 367094 -1300 367150 -1244
rect 367218 -1300 367274 -1244
rect 367342 -1300 367398 -1244
rect 366970 -1424 367026 -1368
rect 367094 -1424 367150 -1368
rect 367218 -1424 367274 -1368
rect 367342 -1424 367398 -1368
rect 366970 -1548 367026 -1492
rect 367094 -1548 367150 -1492
rect 367218 -1548 367274 -1492
rect 367342 -1548 367398 -1492
rect 383852 24362 383908 24418
rect 399250 40294 399306 40350
rect 399374 40294 399430 40350
rect 399498 40294 399554 40350
rect 399622 40294 399678 40350
rect 399250 40170 399306 40226
rect 399374 40170 399430 40226
rect 399498 40170 399554 40226
rect 399622 40170 399678 40226
rect 399250 40046 399306 40102
rect 399374 40046 399430 40102
rect 399498 40046 399554 40102
rect 399622 40046 399678 40102
rect 399250 39922 399306 39978
rect 399374 39922 399430 39978
rect 399498 39922 399554 39978
rect 399622 39922 399678 39978
rect 394828 29596 394884 29638
rect 394828 29582 394884 29596
rect 384970 28294 385026 28350
rect 385094 28294 385150 28350
rect 385218 28294 385274 28350
rect 385342 28294 385398 28350
rect 384970 28170 385026 28226
rect 385094 28170 385150 28226
rect 385218 28170 385274 28226
rect 385342 28170 385398 28226
rect 384970 28046 385026 28102
rect 385094 28046 385150 28102
rect 385218 28046 385274 28102
rect 385342 28046 385398 28102
rect 384970 27922 385026 27978
rect 385094 27922 385150 27978
rect 385218 27922 385274 27978
rect 385342 27922 385398 27978
rect 381250 22294 381306 22350
rect 381374 22294 381430 22350
rect 381498 22294 381554 22350
rect 381622 22294 381678 22350
rect 381250 22170 381306 22226
rect 381374 22170 381430 22226
rect 381498 22170 381554 22226
rect 381622 22170 381678 22226
rect 381250 22046 381306 22102
rect 381374 22046 381430 22102
rect 381498 22046 381554 22102
rect 381622 22046 381678 22102
rect 381250 21922 381306 21978
rect 381374 21922 381430 21978
rect 381498 21922 381554 21978
rect 381622 21922 381678 21978
rect 381250 4294 381306 4350
rect 381374 4294 381430 4350
rect 381498 4294 381554 4350
rect 381622 4294 381678 4350
rect 381250 4170 381306 4226
rect 381374 4170 381430 4226
rect 381498 4170 381554 4226
rect 381622 4170 381678 4226
rect 381250 4046 381306 4102
rect 381374 4046 381430 4102
rect 381498 4046 381554 4102
rect 381622 4046 381678 4102
rect 381250 3922 381306 3978
rect 381374 3922 381430 3978
rect 381498 3922 381554 3978
rect 381622 3922 381678 3978
rect 381250 -216 381306 -160
rect 381374 -216 381430 -160
rect 381498 -216 381554 -160
rect 381622 -216 381678 -160
rect 381250 -340 381306 -284
rect 381374 -340 381430 -284
rect 381498 -340 381554 -284
rect 381622 -340 381678 -284
rect 381250 -464 381306 -408
rect 381374 -464 381430 -408
rect 381498 -464 381554 -408
rect 381622 -464 381678 -408
rect 381250 -588 381306 -532
rect 381374 -588 381430 -532
rect 381498 -588 381554 -532
rect 381622 -588 381678 -532
rect 384970 10294 385026 10350
rect 385094 10294 385150 10350
rect 385218 10294 385274 10350
rect 385342 10294 385398 10350
rect 384970 10170 385026 10226
rect 385094 10170 385150 10226
rect 385218 10170 385274 10226
rect 385342 10170 385398 10226
rect 384970 10046 385026 10102
rect 385094 10046 385150 10102
rect 385218 10046 385274 10102
rect 385342 10046 385398 10102
rect 384970 9922 385026 9978
rect 385094 9922 385150 9978
rect 385218 9922 385274 9978
rect 385342 9922 385398 9978
rect 384970 -1176 385026 -1120
rect 385094 -1176 385150 -1120
rect 385218 -1176 385274 -1120
rect 385342 -1176 385398 -1120
rect 384970 -1300 385026 -1244
rect 385094 -1300 385150 -1244
rect 385218 -1300 385274 -1244
rect 385342 -1300 385398 -1244
rect 384970 -1424 385026 -1368
rect 385094 -1424 385150 -1368
rect 385218 -1424 385274 -1368
rect 385342 -1424 385398 -1368
rect 384970 -1548 385026 -1492
rect 385094 -1548 385150 -1492
rect 385218 -1548 385274 -1492
rect 385342 -1548 385398 -1492
rect 399250 22294 399306 22350
rect 399374 22294 399430 22350
rect 399498 22294 399554 22350
rect 399622 22294 399678 22350
rect 399250 22170 399306 22226
rect 399374 22170 399430 22226
rect 399498 22170 399554 22226
rect 399622 22170 399678 22226
rect 399250 22046 399306 22102
rect 399374 22046 399430 22102
rect 399498 22046 399554 22102
rect 399622 22046 399678 22102
rect 399250 21922 399306 21978
rect 399374 21922 399430 21978
rect 399498 21922 399554 21978
rect 399622 21922 399678 21978
rect 399250 4294 399306 4350
rect 399374 4294 399430 4350
rect 399498 4294 399554 4350
rect 399622 4294 399678 4350
rect 399250 4170 399306 4226
rect 399374 4170 399430 4226
rect 399498 4170 399554 4226
rect 399622 4170 399678 4226
rect 399250 4046 399306 4102
rect 399374 4046 399430 4102
rect 399498 4046 399554 4102
rect 399622 4046 399678 4102
rect 399250 3922 399306 3978
rect 399374 3922 399430 3978
rect 399498 3922 399554 3978
rect 399622 3922 399678 3978
rect 399250 -216 399306 -160
rect 399374 -216 399430 -160
rect 399498 -216 399554 -160
rect 399622 -216 399678 -160
rect 399250 -340 399306 -284
rect 399374 -340 399430 -284
rect 399498 -340 399554 -284
rect 399622 -340 399678 -284
rect 399250 -464 399306 -408
rect 399374 -464 399430 -408
rect 399498 -464 399554 -408
rect 399622 -464 399678 -408
rect 399250 -588 399306 -532
rect 399374 -588 399430 -532
rect 399498 -588 399554 -532
rect 399622 -588 399678 -532
rect 402970 28294 403026 28350
rect 403094 28294 403150 28350
rect 403218 28294 403274 28350
rect 403342 28294 403398 28350
rect 402970 28170 403026 28226
rect 403094 28170 403150 28226
rect 403218 28170 403274 28226
rect 403342 28170 403398 28226
rect 402970 28046 403026 28102
rect 403094 28046 403150 28102
rect 403218 28046 403274 28102
rect 403342 28046 403398 28102
rect 402970 27922 403026 27978
rect 403094 27922 403150 27978
rect 403218 27922 403274 27978
rect 403342 27922 403398 27978
rect 402970 10294 403026 10350
rect 403094 10294 403150 10350
rect 403218 10294 403274 10350
rect 403342 10294 403398 10350
rect 402970 10170 403026 10226
rect 403094 10170 403150 10226
rect 403218 10170 403274 10226
rect 403342 10170 403398 10226
rect 402970 10046 403026 10102
rect 403094 10046 403150 10102
rect 403218 10046 403274 10102
rect 403342 10046 403398 10102
rect 402970 9922 403026 9978
rect 403094 9922 403150 9978
rect 403218 9922 403274 9978
rect 403342 9922 403398 9978
rect 402970 -1176 403026 -1120
rect 403094 -1176 403150 -1120
rect 403218 -1176 403274 -1120
rect 403342 -1176 403398 -1120
rect 402970 -1300 403026 -1244
rect 403094 -1300 403150 -1244
rect 403218 -1300 403274 -1244
rect 403342 -1300 403398 -1244
rect 402970 -1424 403026 -1368
rect 403094 -1424 403150 -1368
rect 403218 -1424 403274 -1368
rect 403342 -1424 403398 -1368
rect 402970 -1548 403026 -1492
rect 403094 -1548 403150 -1492
rect 403218 -1548 403274 -1492
rect 403342 -1548 403398 -1492
rect 417250 40294 417306 40350
rect 417374 40294 417430 40350
rect 417498 40294 417554 40350
rect 417622 40294 417678 40350
rect 417250 40170 417306 40226
rect 417374 40170 417430 40226
rect 417498 40170 417554 40226
rect 417622 40170 417678 40226
rect 417250 40046 417306 40102
rect 417374 40046 417430 40102
rect 417498 40046 417554 40102
rect 417622 40046 417678 40102
rect 417250 39922 417306 39978
rect 417374 39922 417430 39978
rect 417498 39922 417554 39978
rect 417622 39922 417678 39978
rect 418348 39662 418404 39718
rect 419692 39676 419748 39718
rect 419692 39662 419748 39676
rect 418348 34442 418404 34498
rect 417250 22294 417306 22350
rect 417374 22294 417430 22350
rect 417498 22294 417554 22350
rect 417622 22294 417678 22350
rect 417250 22170 417306 22226
rect 417374 22170 417430 22226
rect 417498 22170 417554 22226
rect 417622 22170 417678 22226
rect 417250 22046 417306 22102
rect 417374 22046 417430 22102
rect 417498 22046 417554 22102
rect 417622 22046 417678 22102
rect 417250 21922 417306 21978
rect 417374 21922 417430 21978
rect 417498 21922 417554 21978
rect 417622 21922 417678 21978
rect 417250 4294 417306 4350
rect 417374 4294 417430 4350
rect 417498 4294 417554 4350
rect 417622 4294 417678 4350
rect 417250 4170 417306 4226
rect 417374 4170 417430 4226
rect 417498 4170 417554 4226
rect 417622 4170 417678 4226
rect 417250 4046 417306 4102
rect 417374 4046 417430 4102
rect 417498 4046 417554 4102
rect 417622 4046 417678 4102
rect 417250 3922 417306 3978
rect 417374 3922 417430 3978
rect 417498 3922 417554 3978
rect 417622 3922 417678 3978
rect 417250 -216 417306 -160
rect 417374 -216 417430 -160
rect 417498 -216 417554 -160
rect 417622 -216 417678 -160
rect 417250 -340 417306 -284
rect 417374 -340 417430 -284
rect 417498 -340 417554 -284
rect 417622 -340 417678 -284
rect 417250 -464 417306 -408
rect 417374 -464 417430 -408
rect 417498 -464 417554 -408
rect 417622 -464 417678 -408
rect 417250 -588 417306 -532
rect 417374 -588 417430 -532
rect 417498 -588 417554 -532
rect 417622 -588 417678 -532
rect 431788 41102 431844 41158
rect 423388 35162 423444 35218
rect 431788 29402 431844 29458
rect 435250 40294 435306 40350
rect 435374 40294 435430 40350
rect 435498 40294 435554 40350
rect 435622 40294 435678 40350
rect 435250 40170 435306 40226
rect 435374 40170 435430 40226
rect 435498 40170 435554 40226
rect 435622 40170 435678 40226
rect 435250 40046 435306 40102
rect 435374 40046 435430 40102
rect 435498 40046 435554 40102
rect 435622 40046 435678 40102
rect 435250 39922 435306 39978
rect 435374 39922 435430 39978
rect 435498 39922 435554 39978
rect 435622 39922 435678 39978
rect 420970 28294 421026 28350
rect 421094 28294 421150 28350
rect 421218 28294 421274 28350
rect 421342 28294 421398 28350
rect 420970 28170 421026 28226
rect 421094 28170 421150 28226
rect 421218 28170 421274 28226
rect 421342 28170 421398 28226
rect 420970 28046 421026 28102
rect 421094 28046 421150 28102
rect 421218 28046 421274 28102
rect 421342 28046 421398 28102
rect 420970 27922 421026 27978
rect 421094 27922 421150 27978
rect 421218 27922 421274 27978
rect 421342 27922 421398 27978
rect 420970 10294 421026 10350
rect 421094 10294 421150 10350
rect 421218 10294 421274 10350
rect 421342 10294 421398 10350
rect 420970 10170 421026 10226
rect 421094 10170 421150 10226
rect 421218 10170 421274 10226
rect 421342 10170 421398 10226
rect 420970 10046 421026 10102
rect 421094 10046 421150 10102
rect 421218 10046 421274 10102
rect 421342 10046 421398 10102
rect 420970 9922 421026 9978
rect 421094 9922 421150 9978
rect 421218 9922 421274 9978
rect 421342 9922 421398 9978
rect 420970 -1176 421026 -1120
rect 421094 -1176 421150 -1120
rect 421218 -1176 421274 -1120
rect 421342 -1176 421398 -1120
rect 420970 -1300 421026 -1244
rect 421094 -1300 421150 -1244
rect 421218 -1300 421274 -1244
rect 421342 -1300 421398 -1244
rect 420970 -1424 421026 -1368
rect 421094 -1424 421150 -1368
rect 421218 -1424 421274 -1368
rect 421342 -1424 421398 -1368
rect 420970 -1548 421026 -1492
rect 421094 -1548 421150 -1492
rect 421218 -1548 421274 -1492
rect 421342 -1548 421398 -1492
rect 435250 22294 435306 22350
rect 435374 22294 435430 22350
rect 435498 22294 435554 22350
rect 435622 22294 435678 22350
rect 435250 22170 435306 22226
rect 435374 22170 435430 22226
rect 435498 22170 435554 22226
rect 435622 22170 435678 22226
rect 435250 22046 435306 22102
rect 435374 22046 435430 22102
rect 435498 22046 435554 22102
rect 435622 22046 435678 22102
rect 435250 21922 435306 21978
rect 435374 21922 435430 21978
rect 435498 21922 435554 21978
rect 435622 21922 435678 21978
rect 435250 4294 435306 4350
rect 435374 4294 435430 4350
rect 435498 4294 435554 4350
rect 435622 4294 435678 4350
rect 435250 4170 435306 4226
rect 435374 4170 435430 4226
rect 435498 4170 435554 4226
rect 435622 4170 435678 4226
rect 435250 4046 435306 4102
rect 435374 4046 435430 4102
rect 435498 4046 435554 4102
rect 435622 4046 435678 4102
rect 435250 3922 435306 3978
rect 435374 3922 435430 3978
rect 435498 3922 435554 3978
rect 435622 3922 435678 3978
rect 435250 -216 435306 -160
rect 435374 -216 435430 -160
rect 435498 -216 435554 -160
rect 435622 -216 435678 -160
rect 435250 -340 435306 -284
rect 435374 -340 435430 -284
rect 435498 -340 435554 -284
rect 435622 -340 435678 -284
rect 435250 -464 435306 -408
rect 435374 -464 435430 -408
rect 435498 -464 435554 -408
rect 435622 -464 435678 -408
rect 435250 -588 435306 -532
rect 435374 -588 435430 -532
rect 435498 -588 435554 -532
rect 435622 -588 435678 -532
rect 453250 40294 453306 40350
rect 453374 40294 453430 40350
rect 453498 40294 453554 40350
rect 453622 40294 453678 40350
rect 453250 40170 453306 40226
rect 453374 40170 453430 40226
rect 453498 40170 453554 40226
rect 453622 40170 453678 40226
rect 453250 40046 453306 40102
rect 453374 40046 453430 40102
rect 453498 40046 453554 40102
rect 453622 40046 453678 40102
rect 453250 39922 453306 39978
rect 453374 39922 453430 39978
rect 453498 39922 453554 39978
rect 453622 39922 453678 39978
rect 451948 39508 452004 39538
rect 451948 39482 452004 39508
rect 438970 28294 439026 28350
rect 439094 28294 439150 28350
rect 439218 28294 439274 28350
rect 439342 28294 439398 28350
rect 438970 28170 439026 28226
rect 439094 28170 439150 28226
rect 439218 28170 439274 28226
rect 439342 28170 439398 28226
rect 438970 28046 439026 28102
rect 439094 28046 439150 28102
rect 439218 28046 439274 28102
rect 439342 28046 439398 28102
rect 438970 27922 439026 27978
rect 439094 27922 439150 27978
rect 439218 27922 439274 27978
rect 439342 27922 439398 27978
rect 438970 10294 439026 10350
rect 439094 10294 439150 10350
rect 439218 10294 439274 10350
rect 439342 10294 439398 10350
rect 438970 10170 439026 10226
rect 439094 10170 439150 10226
rect 439218 10170 439274 10226
rect 439342 10170 439398 10226
rect 438970 10046 439026 10102
rect 439094 10046 439150 10102
rect 439218 10046 439274 10102
rect 439342 10046 439398 10102
rect 438970 9922 439026 9978
rect 439094 9922 439150 9978
rect 439218 9922 439274 9978
rect 439342 9922 439398 9978
rect 438970 -1176 439026 -1120
rect 439094 -1176 439150 -1120
rect 439218 -1176 439274 -1120
rect 439342 -1176 439398 -1120
rect 438970 -1300 439026 -1244
rect 439094 -1300 439150 -1244
rect 439218 -1300 439274 -1244
rect 439342 -1300 439398 -1244
rect 438970 -1424 439026 -1368
rect 439094 -1424 439150 -1368
rect 439218 -1424 439274 -1368
rect 439342 -1424 439398 -1368
rect 438970 -1548 439026 -1492
rect 439094 -1548 439150 -1492
rect 439218 -1548 439274 -1492
rect 439342 -1548 439398 -1492
rect 453250 22294 453306 22350
rect 453374 22294 453430 22350
rect 453498 22294 453554 22350
rect 453622 22294 453678 22350
rect 453250 22170 453306 22226
rect 453374 22170 453430 22226
rect 453498 22170 453554 22226
rect 453622 22170 453678 22226
rect 453250 22046 453306 22102
rect 453374 22046 453430 22102
rect 453498 22046 453554 22102
rect 453622 22046 453678 22102
rect 453250 21922 453306 21978
rect 453374 21922 453430 21978
rect 453498 21922 453554 21978
rect 453622 21922 453678 21978
rect 453250 4294 453306 4350
rect 453374 4294 453430 4350
rect 453498 4294 453554 4350
rect 453622 4294 453678 4350
rect 453250 4170 453306 4226
rect 453374 4170 453430 4226
rect 453498 4170 453554 4226
rect 453622 4170 453678 4226
rect 453250 4046 453306 4102
rect 453374 4046 453430 4102
rect 453498 4046 453554 4102
rect 453622 4046 453678 4102
rect 453250 3922 453306 3978
rect 453374 3922 453430 3978
rect 453498 3922 453554 3978
rect 453622 3922 453678 3978
rect 453250 -216 453306 -160
rect 453374 -216 453430 -160
rect 453498 -216 453554 -160
rect 453622 -216 453678 -160
rect 453250 -340 453306 -284
rect 453374 -340 453430 -284
rect 453498 -340 453554 -284
rect 453622 -340 453678 -284
rect 453250 -464 453306 -408
rect 453374 -464 453430 -408
rect 453498 -464 453554 -408
rect 453622 -464 453678 -408
rect 453250 -588 453306 -532
rect 453374 -588 453430 -532
rect 453498 -588 453554 -532
rect 453622 -588 453678 -532
rect 460012 39340 460068 39358
rect 460012 39302 460068 39340
rect 471250 40294 471306 40350
rect 471374 40294 471430 40350
rect 471498 40294 471554 40350
rect 471622 40294 471678 40350
rect 471250 40170 471306 40226
rect 471374 40170 471430 40226
rect 471498 40170 471554 40226
rect 471622 40170 471678 40226
rect 471250 40046 471306 40102
rect 471374 40046 471430 40102
rect 471498 40046 471554 40102
rect 471622 40046 471678 40102
rect 471250 39922 471306 39978
rect 471374 39922 471430 39978
rect 471498 39922 471554 39978
rect 471622 39922 471678 39978
rect 463708 31742 463764 31798
rect 456970 28294 457026 28350
rect 457094 28294 457150 28350
rect 457218 28294 457274 28350
rect 457342 28294 457398 28350
rect 456970 28170 457026 28226
rect 457094 28170 457150 28226
rect 457218 28170 457274 28226
rect 457342 28170 457398 28226
rect 456970 28046 457026 28102
rect 457094 28046 457150 28102
rect 457218 28046 457274 28102
rect 457342 28046 457398 28102
rect 456970 27922 457026 27978
rect 457094 27922 457150 27978
rect 457218 27922 457274 27978
rect 457342 27922 457398 27978
rect 456970 10294 457026 10350
rect 457094 10294 457150 10350
rect 457218 10294 457274 10350
rect 457342 10294 457398 10350
rect 456970 10170 457026 10226
rect 457094 10170 457150 10226
rect 457218 10170 457274 10226
rect 457342 10170 457398 10226
rect 456970 10046 457026 10102
rect 457094 10046 457150 10102
rect 457218 10046 457274 10102
rect 457342 10046 457398 10102
rect 456970 9922 457026 9978
rect 457094 9922 457150 9978
rect 457218 9922 457274 9978
rect 457342 9922 457398 9978
rect 456970 -1176 457026 -1120
rect 457094 -1176 457150 -1120
rect 457218 -1176 457274 -1120
rect 457342 -1176 457398 -1120
rect 456970 -1300 457026 -1244
rect 457094 -1300 457150 -1244
rect 457218 -1300 457274 -1244
rect 457342 -1300 457398 -1244
rect 456970 -1424 457026 -1368
rect 457094 -1424 457150 -1368
rect 457218 -1424 457274 -1368
rect 457342 -1424 457398 -1368
rect 456970 -1548 457026 -1492
rect 457094 -1548 457150 -1492
rect 457218 -1548 457274 -1492
rect 457342 -1548 457398 -1492
rect 471250 22294 471306 22350
rect 471374 22294 471430 22350
rect 471498 22294 471554 22350
rect 471622 22294 471678 22350
rect 471250 22170 471306 22226
rect 471374 22170 471430 22226
rect 471498 22170 471554 22226
rect 471622 22170 471678 22226
rect 471250 22046 471306 22102
rect 471374 22046 471430 22102
rect 471498 22046 471554 22102
rect 471622 22046 471678 22102
rect 471250 21922 471306 21978
rect 471374 21922 471430 21978
rect 471498 21922 471554 21978
rect 471622 21922 471678 21978
rect 471250 4294 471306 4350
rect 471374 4294 471430 4350
rect 471498 4294 471554 4350
rect 471622 4294 471678 4350
rect 471250 4170 471306 4226
rect 471374 4170 471430 4226
rect 471498 4170 471554 4226
rect 471622 4170 471678 4226
rect 471250 4046 471306 4102
rect 471374 4046 471430 4102
rect 471498 4046 471554 4102
rect 471622 4046 471678 4102
rect 471250 3922 471306 3978
rect 471374 3922 471430 3978
rect 471498 3922 471554 3978
rect 471622 3922 471678 3978
rect 471250 -216 471306 -160
rect 471374 -216 471430 -160
rect 471498 -216 471554 -160
rect 471622 -216 471678 -160
rect 471250 -340 471306 -284
rect 471374 -340 471430 -284
rect 471498 -340 471554 -284
rect 471622 -340 471678 -284
rect 471250 -464 471306 -408
rect 471374 -464 471430 -408
rect 471498 -464 471554 -408
rect 471622 -464 471678 -408
rect 471250 -588 471306 -532
rect 471374 -588 471430 -532
rect 471498 -588 471554 -532
rect 471622 -588 471678 -532
rect 489250 40294 489306 40350
rect 489374 40294 489430 40350
rect 489498 40294 489554 40350
rect 489622 40294 489678 40350
rect 489250 40170 489306 40226
rect 489374 40170 489430 40226
rect 489498 40170 489554 40226
rect 489622 40170 489678 40226
rect 489250 40046 489306 40102
rect 489374 40046 489430 40102
rect 489498 40046 489554 40102
rect 489622 40046 489678 40102
rect 489250 39922 489306 39978
rect 489374 39922 489430 39978
rect 489498 39922 489554 39978
rect 489622 39922 489678 39978
rect 478828 31562 478884 31618
rect 483868 31382 483924 31438
rect 487228 31202 487284 31258
rect 474970 28294 475026 28350
rect 475094 28294 475150 28350
rect 475218 28294 475274 28350
rect 475342 28294 475398 28350
rect 474970 28170 475026 28226
rect 475094 28170 475150 28226
rect 475218 28170 475274 28226
rect 475342 28170 475398 28226
rect 474970 28046 475026 28102
rect 475094 28046 475150 28102
rect 475218 28046 475274 28102
rect 475342 28046 475398 28102
rect 474970 27922 475026 27978
rect 475094 27922 475150 27978
rect 475218 27922 475274 27978
rect 475342 27922 475398 27978
rect 474970 10294 475026 10350
rect 475094 10294 475150 10350
rect 475218 10294 475274 10350
rect 475342 10294 475398 10350
rect 474970 10170 475026 10226
rect 475094 10170 475150 10226
rect 475218 10170 475274 10226
rect 475342 10170 475398 10226
rect 474970 10046 475026 10102
rect 475094 10046 475150 10102
rect 475218 10046 475274 10102
rect 475342 10046 475398 10102
rect 474970 9922 475026 9978
rect 475094 9922 475150 9978
rect 475218 9922 475274 9978
rect 475342 9922 475398 9978
rect 474970 -1176 475026 -1120
rect 475094 -1176 475150 -1120
rect 475218 -1176 475274 -1120
rect 475342 -1176 475398 -1120
rect 474970 -1300 475026 -1244
rect 475094 -1300 475150 -1244
rect 475218 -1300 475274 -1244
rect 475342 -1300 475398 -1244
rect 474970 -1424 475026 -1368
rect 475094 -1424 475150 -1368
rect 475218 -1424 475274 -1368
rect 475342 -1424 475398 -1368
rect 474970 -1548 475026 -1492
rect 475094 -1548 475150 -1492
rect 475218 -1548 475274 -1492
rect 475342 -1548 475398 -1492
rect 489250 22294 489306 22350
rect 489374 22294 489430 22350
rect 489498 22294 489554 22350
rect 489622 22294 489678 22350
rect 489250 22170 489306 22226
rect 489374 22170 489430 22226
rect 489498 22170 489554 22226
rect 489622 22170 489678 22226
rect 489250 22046 489306 22102
rect 489374 22046 489430 22102
rect 489498 22046 489554 22102
rect 489622 22046 489678 22102
rect 489250 21922 489306 21978
rect 489374 21922 489430 21978
rect 489498 21922 489554 21978
rect 489622 21922 489678 21978
rect 489250 4294 489306 4350
rect 489374 4294 489430 4350
rect 489498 4294 489554 4350
rect 489622 4294 489678 4350
rect 489250 4170 489306 4226
rect 489374 4170 489430 4226
rect 489498 4170 489554 4226
rect 489622 4170 489678 4226
rect 489250 4046 489306 4102
rect 489374 4046 489430 4102
rect 489498 4046 489554 4102
rect 489622 4046 489678 4102
rect 489250 3922 489306 3978
rect 489374 3922 489430 3978
rect 489498 3922 489554 3978
rect 489622 3922 489678 3978
rect 489250 -216 489306 -160
rect 489374 -216 489430 -160
rect 489498 -216 489554 -160
rect 489622 -216 489678 -160
rect 489250 -340 489306 -284
rect 489374 -340 489430 -284
rect 489498 -340 489554 -284
rect 489622 -340 489678 -284
rect 489250 -464 489306 -408
rect 489374 -464 489430 -408
rect 489498 -464 489554 -408
rect 489622 -464 489678 -408
rect 489250 -588 489306 -532
rect 489374 -588 489430 -532
rect 489498 -588 489554 -532
rect 489622 -588 489678 -532
rect 507250 40294 507306 40350
rect 507374 40294 507430 40350
rect 507498 40294 507554 40350
rect 507622 40294 507678 40350
rect 507250 40170 507306 40226
rect 507374 40170 507430 40226
rect 507498 40170 507554 40226
rect 507622 40170 507678 40226
rect 507250 40046 507306 40102
rect 507374 40046 507430 40102
rect 507498 40046 507554 40102
rect 507622 40046 507678 40102
rect 507250 39922 507306 39978
rect 507374 39922 507430 39978
rect 507498 39922 507554 39978
rect 507622 39922 507678 39978
rect 504812 31022 504868 31078
rect 500332 29762 500388 29818
rect 492970 28294 493026 28350
rect 493094 28294 493150 28350
rect 493218 28294 493274 28350
rect 493342 28294 493398 28350
rect 492970 28170 493026 28226
rect 493094 28170 493150 28226
rect 493218 28170 493274 28226
rect 493342 28170 493398 28226
rect 492970 28046 493026 28102
rect 493094 28046 493150 28102
rect 493218 28046 493274 28102
rect 493342 28046 493398 28102
rect 492970 27922 493026 27978
rect 493094 27922 493150 27978
rect 493218 27922 493274 27978
rect 493342 27922 493398 27978
rect 492970 10294 493026 10350
rect 493094 10294 493150 10350
rect 493218 10294 493274 10350
rect 493342 10294 493398 10350
rect 492970 10170 493026 10226
rect 493094 10170 493150 10226
rect 493218 10170 493274 10226
rect 493342 10170 493398 10226
rect 492970 10046 493026 10102
rect 493094 10046 493150 10102
rect 493218 10046 493274 10102
rect 493342 10046 493398 10102
rect 492970 9922 493026 9978
rect 493094 9922 493150 9978
rect 493218 9922 493274 9978
rect 493342 9922 493398 9978
rect 492970 -1176 493026 -1120
rect 493094 -1176 493150 -1120
rect 493218 -1176 493274 -1120
rect 493342 -1176 493398 -1120
rect 492970 -1300 493026 -1244
rect 493094 -1300 493150 -1244
rect 493218 -1300 493274 -1244
rect 493342 -1300 493398 -1244
rect 492970 -1424 493026 -1368
rect 493094 -1424 493150 -1368
rect 493218 -1424 493274 -1368
rect 493342 -1424 493398 -1368
rect 492970 -1548 493026 -1492
rect 493094 -1548 493150 -1492
rect 493218 -1548 493274 -1492
rect 493342 -1548 493398 -1492
rect 507250 22294 507306 22350
rect 507374 22294 507430 22350
rect 507498 22294 507554 22350
rect 507622 22294 507678 22350
rect 507250 22170 507306 22226
rect 507374 22170 507430 22226
rect 507498 22170 507554 22226
rect 507622 22170 507678 22226
rect 507250 22046 507306 22102
rect 507374 22046 507430 22102
rect 507498 22046 507554 22102
rect 507622 22046 507678 22102
rect 507250 21922 507306 21978
rect 507374 21922 507430 21978
rect 507498 21922 507554 21978
rect 507622 21922 507678 21978
rect 507250 4294 507306 4350
rect 507374 4294 507430 4350
rect 507498 4294 507554 4350
rect 507622 4294 507678 4350
rect 507250 4170 507306 4226
rect 507374 4170 507430 4226
rect 507498 4170 507554 4226
rect 507622 4170 507678 4226
rect 507250 4046 507306 4102
rect 507374 4046 507430 4102
rect 507498 4046 507554 4102
rect 507622 4046 507678 4102
rect 507250 3922 507306 3978
rect 507374 3922 507430 3978
rect 507498 3922 507554 3978
rect 507622 3922 507678 3978
rect 507250 -216 507306 -160
rect 507374 -216 507430 -160
rect 507498 -216 507554 -160
rect 507622 -216 507678 -160
rect 507250 -340 507306 -284
rect 507374 -340 507430 -284
rect 507498 -340 507554 -284
rect 507622 -340 507678 -284
rect 507250 -464 507306 -408
rect 507374 -464 507430 -408
rect 507498 -464 507554 -408
rect 507622 -464 507678 -408
rect 507250 -588 507306 -532
rect 507374 -588 507430 -532
rect 507498 -588 507554 -532
rect 507622 -588 507678 -532
rect 512428 33182 512484 33238
rect 532700 41462 532756 41518
rect 525250 40294 525306 40350
rect 525374 40294 525430 40350
rect 525498 40294 525554 40350
rect 525622 40294 525678 40350
rect 525250 40170 525306 40226
rect 525374 40170 525430 40226
rect 525498 40170 525554 40226
rect 525622 40170 525678 40226
rect 525250 40046 525306 40102
rect 525374 40046 525430 40102
rect 525498 40046 525554 40102
rect 525622 40046 525678 40102
rect 525250 39922 525306 39978
rect 525374 39922 525430 39978
rect 525498 39922 525554 39978
rect 525622 39922 525678 39978
rect 524524 33002 524580 33058
rect 519148 30122 519204 30178
rect 516460 29942 516516 29998
rect 510970 28294 511026 28350
rect 511094 28294 511150 28350
rect 511218 28294 511274 28350
rect 511342 28294 511398 28350
rect 510970 28170 511026 28226
rect 511094 28170 511150 28226
rect 511218 28170 511274 28226
rect 511342 28170 511398 28226
rect 510970 28046 511026 28102
rect 511094 28046 511150 28102
rect 511218 28046 511274 28102
rect 511342 28046 511398 28102
rect 510970 27922 511026 27978
rect 511094 27922 511150 27978
rect 511218 27922 511274 27978
rect 511342 27922 511398 27978
rect 510970 10294 511026 10350
rect 511094 10294 511150 10350
rect 511218 10294 511274 10350
rect 511342 10294 511398 10350
rect 510970 10170 511026 10226
rect 511094 10170 511150 10226
rect 511218 10170 511274 10226
rect 511342 10170 511398 10226
rect 510970 10046 511026 10102
rect 511094 10046 511150 10102
rect 511218 10046 511274 10102
rect 511342 10046 511398 10102
rect 510970 9922 511026 9978
rect 511094 9922 511150 9978
rect 511218 9922 511274 9978
rect 511342 9922 511398 9978
rect 510970 -1176 511026 -1120
rect 511094 -1176 511150 -1120
rect 511218 -1176 511274 -1120
rect 511342 -1176 511398 -1120
rect 510970 -1300 511026 -1244
rect 511094 -1300 511150 -1244
rect 511218 -1300 511274 -1244
rect 511342 -1300 511398 -1244
rect 510970 -1424 511026 -1368
rect 511094 -1424 511150 -1368
rect 511218 -1424 511274 -1368
rect 511342 -1424 511398 -1368
rect 510970 -1548 511026 -1492
rect 511094 -1548 511150 -1492
rect 511218 -1548 511274 -1492
rect 511342 -1548 511398 -1492
rect 528556 32822 528612 32878
rect 525250 22294 525306 22350
rect 525374 22294 525430 22350
rect 525498 22294 525554 22350
rect 525622 22294 525678 22350
rect 525250 22170 525306 22226
rect 525374 22170 525430 22226
rect 525498 22170 525554 22226
rect 525622 22170 525678 22226
rect 525250 22046 525306 22102
rect 525374 22046 525430 22102
rect 525498 22046 525554 22102
rect 525622 22046 525678 22102
rect 525250 21922 525306 21978
rect 525374 21922 525430 21978
rect 525498 21922 525554 21978
rect 525622 21922 525678 21978
rect 525250 4294 525306 4350
rect 525374 4294 525430 4350
rect 525498 4294 525554 4350
rect 525622 4294 525678 4350
rect 525250 4170 525306 4226
rect 525374 4170 525430 4226
rect 525498 4170 525554 4226
rect 525622 4170 525678 4226
rect 525250 4046 525306 4102
rect 525374 4046 525430 4102
rect 525498 4046 525554 4102
rect 525622 4046 525678 4102
rect 525250 3922 525306 3978
rect 525374 3922 525430 3978
rect 525498 3922 525554 3978
rect 525622 3922 525678 3978
rect 525250 -216 525306 -160
rect 525374 -216 525430 -160
rect 525498 -216 525554 -160
rect 525622 -216 525678 -160
rect 525250 -340 525306 -284
rect 525374 -340 525430 -284
rect 525498 -340 525554 -284
rect 525622 -340 525678 -284
rect 525250 -464 525306 -408
rect 525374 -464 525430 -408
rect 525498 -464 525554 -408
rect 525622 -464 525678 -408
rect 525250 -588 525306 -532
rect 525374 -588 525430 -532
rect 525498 -588 525554 -532
rect 525622 -588 525678 -532
rect 543250 40294 543306 40350
rect 543374 40294 543430 40350
rect 543498 40294 543554 40350
rect 543622 40294 543678 40350
rect 543250 40170 543306 40226
rect 543374 40170 543430 40226
rect 543498 40170 543554 40226
rect 543622 40170 543678 40226
rect 543250 40046 543306 40102
rect 543374 40046 543430 40102
rect 543498 40046 543554 40102
rect 543622 40046 543678 40102
rect 543250 39922 543306 39978
rect 543374 39922 543430 39978
rect 543498 39922 543554 39978
rect 543622 39922 543678 39978
rect 532588 32642 532644 32698
rect 528970 28294 529026 28350
rect 529094 28294 529150 28350
rect 529218 28294 529274 28350
rect 529342 28294 529398 28350
rect 528970 28170 529026 28226
rect 529094 28170 529150 28226
rect 529218 28170 529274 28226
rect 529342 28170 529398 28226
rect 528970 28046 529026 28102
rect 529094 28046 529150 28102
rect 529218 28046 529274 28102
rect 529342 28046 529398 28102
rect 528970 27922 529026 27978
rect 529094 27922 529150 27978
rect 529218 27922 529274 27978
rect 529342 27922 529398 27978
rect 528970 10294 529026 10350
rect 529094 10294 529150 10350
rect 529218 10294 529274 10350
rect 529342 10294 529398 10350
rect 528970 10170 529026 10226
rect 529094 10170 529150 10226
rect 529218 10170 529274 10226
rect 529342 10170 529398 10226
rect 528970 10046 529026 10102
rect 529094 10046 529150 10102
rect 529218 10046 529274 10102
rect 529342 10046 529398 10102
rect 528970 9922 529026 9978
rect 529094 9922 529150 9978
rect 529218 9922 529274 9978
rect 529342 9922 529398 9978
rect 528970 -1176 529026 -1120
rect 529094 -1176 529150 -1120
rect 529218 -1176 529274 -1120
rect 529342 -1176 529398 -1120
rect 528970 -1300 529026 -1244
rect 529094 -1300 529150 -1244
rect 529218 -1300 529274 -1244
rect 529342 -1300 529398 -1244
rect 528970 -1424 529026 -1368
rect 529094 -1424 529150 -1368
rect 529218 -1424 529274 -1368
rect 529342 -1424 529398 -1368
rect 528970 -1548 529026 -1492
rect 529094 -1548 529150 -1492
rect 529218 -1548 529274 -1492
rect 529342 -1548 529398 -1492
rect 546028 37884 546084 37918
rect 546028 37862 546084 37884
rect 543250 22294 543306 22350
rect 543374 22294 543430 22350
rect 543498 22294 543554 22350
rect 543622 22294 543678 22350
rect 543250 22170 543306 22226
rect 543374 22170 543430 22226
rect 543498 22170 543554 22226
rect 543622 22170 543678 22226
rect 543250 22046 543306 22102
rect 543374 22046 543430 22102
rect 543498 22046 543554 22102
rect 543622 22046 543678 22102
rect 543250 21922 543306 21978
rect 543374 21922 543430 21978
rect 543498 21922 543554 21978
rect 543622 21922 543678 21978
rect 543250 4294 543306 4350
rect 543374 4294 543430 4350
rect 543498 4294 543554 4350
rect 543622 4294 543678 4350
rect 543250 4170 543306 4226
rect 543374 4170 543430 4226
rect 543498 4170 543554 4226
rect 543622 4170 543678 4226
rect 543250 4046 543306 4102
rect 543374 4046 543430 4102
rect 543498 4046 543554 4102
rect 543622 4046 543678 4102
rect 543250 3922 543306 3978
rect 543374 3922 543430 3978
rect 543498 3922 543554 3978
rect 543622 3922 543678 3978
rect 543250 -216 543306 -160
rect 543374 -216 543430 -160
rect 543498 -216 543554 -160
rect 543622 -216 543678 -160
rect 543250 -340 543306 -284
rect 543374 -340 543430 -284
rect 543498 -340 543554 -284
rect 543622 -340 543678 -284
rect 543250 -464 543306 -408
rect 543374 -464 543430 -408
rect 543498 -464 543554 -408
rect 543622 -464 543678 -408
rect 543250 -588 543306 -532
rect 543374 -588 543430 -532
rect 543498 -588 543554 -532
rect 543622 -588 543678 -532
rect 546970 28294 547026 28350
rect 547094 28294 547150 28350
rect 547218 28294 547274 28350
rect 547342 28294 547398 28350
rect 546970 28170 547026 28226
rect 547094 28170 547150 28226
rect 547218 28170 547274 28226
rect 547342 28170 547398 28226
rect 546970 28046 547026 28102
rect 547094 28046 547150 28102
rect 547218 28046 547274 28102
rect 547342 28046 547398 28102
rect 546970 27922 547026 27978
rect 547094 27922 547150 27978
rect 547218 27922 547274 27978
rect 547342 27922 547398 27978
rect 548716 51542 548772 51598
rect 548604 49742 548660 49798
rect 546970 10294 547026 10350
rect 547094 10294 547150 10350
rect 547218 10294 547274 10350
rect 547342 10294 547398 10350
rect 546970 10170 547026 10226
rect 547094 10170 547150 10226
rect 547218 10170 547274 10226
rect 547342 10170 547398 10226
rect 546970 10046 547026 10102
rect 547094 10046 547150 10102
rect 547218 10046 547274 10102
rect 547342 10046 547398 10102
rect 546970 9922 547026 9978
rect 547094 9922 547150 9978
rect 547218 9922 547274 9978
rect 547342 9922 547398 9978
rect 549388 54602 549444 54658
rect 549388 51542 549444 51598
rect 549388 49756 549444 49798
rect 549388 49742 549444 49756
rect 550060 59822 550116 59878
rect 549276 35162 549332 35218
rect 550284 41462 550340 41518
rect 550844 38052 550900 38098
rect 550844 38042 550900 38052
rect 551068 42722 551124 42778
rect 551516 27602 551572 27658
rect 551292 27422 551348 27478
rect 551068 11582 551124 11638
rect 553980 44162 554036 44218
rect 554540 41282 554596 41338
rect 555324 44162 555380 44218
rect 556892 42902 556948 42958
rect 554540 37862 554596 37918
rect 554316 36782 554372 36838
rect 557340 47762 557396 47818
rect 557004 37682 557060 37738
rect 554540 29402 554596 29458
rect 554428 26522 554484 26578
rect 554540 25982 554596 26038
rect 554540 25802 554596 25858
rect 552636 11582 552692 11638
rect 552636 10682 552692 10738
rect 556892 29402 556948 29458
rect 557228 38042 557284 38098
rect 557116 26522 557172 26578
rect 557228 13022 557284 13078
rect 559356 43082 559412 43138
rect 558022 40356 558078 40412
rect 558146 40356 558202 40412
rect 558270 40356 558326 40412
rect 558394 40356 558450 40412
rect 558518 40356 558574 40412
rect 558642 40356 558698 40412
rect 558766 40356 558822 40412
rect 558890 40356 558946 40412
rect 559014 40356 559070 40412
rect 559138 40356 559194 40412
rect 558022 40232 558078 40288
rect 558146 40232 558202 40288
rect 558270 40232 558326 40288
rect 558394 40232 558450 40288
rect 558518 40232 558574 40288
rect 558642 40232 558698 40288
rect 558766 40232 558822 40288
rect 558890 40232 558946 40288
rect 559014 40232 559070 40288
rect 559138 40232 559194 40288
rect 558022 40108 558078 40164
rect 558146 40108 558202 40164
rect 558270 40108 558326 40164
rect 558394 40108 558450 40164
rect 558518 40108 558574 40164
rect 558642 40108 558698 40164
rect 558766 40108 558822 40164
rect 558890 40108 558946 40164
rect 559014 40108 559070 40164
rect 559138 40108 559194 40164
rect 558022 39984 558078 40040
rect 558146 39984 558202 40040
rect 558270 39984 558326 40040
rect 558394 39984 558450 40040
rect 558518 39984 558574 40040
rect 558642 39984 558698 40040
rect 558766 39984 558822 40040
rect 558890 39984 558946 40040
rect 559014 39984 559070 40040
rect 559138 39984 559194 40040
rect 558022 39860 558078 39916
rect 558146 39860 558202 39916
rect 558270 39860 558326 39916
rect 558394 39860 558450 39916
rect 558518 39860 558574 39916
rect 558642 39860 558698 39916
rect 558766 39860 558822 39916
rect 558890 39860 558946 39916
rect 559014 39860 559070 39916
rect 559138 39860 559194 39916
rect 568058 460294 568114 460350
rect 568182 460294 568238 460350
rect 568058 460170 568114 460226
rect 568182 460170 568238 460226
rect 568058 460046 568114 460102
rect 568182 460046 568238 460102
rect 568058 459922 568114 459978
rect 568182 459922 568238 459978
rect 574862 460294 574918 460350
rect 574986 460294 575042 460350
rect 574862 460170 574918 460226
rect 574986 460170 575042 460226
rect 574862 460046 574918 460102
rect 574986 460046 575042 460102
rect 574862 459922 574918 459978
rect 574986 459922 575042 459978
rect 581666 460294 581722 460350
rect 581790 460294 581846 460350
rect 581666 460170 581722 460226
rect 581790 460170 581846 460226
rect 581666 460046 581722 460102
rect 581790 460046 581846 460102
rect 581666 459922 581722 459978
rect 581790 459922 581846 459978
rect 588470 460294 588526 460350
rect 588594 460294 588650 460350
rect 588470 460170 588526 460226
rect 588594 460170 588650 460226
rect 588470 460046 588526 460102
rect 588594 460046 588650 460102
rect 588470 459922 588526 459978
rect 588594 459922 588650 459978
rect 559916 41102 559972 41158
rect 564656 454294 564712 454350
rect 564780 454294 564836 454350
rect 564656 454170 564712 454226
rect 564780 454170 564836 454226
rect 564656 454046 564712 454102
rect 564780 454046 564836 454102
rect 564656 453922 564712 453978
rect 564780 453922 564836 453978
rect 571460 454294 571516 454350
rect 571584 454294 571640 454350
rect 571460 454170 571516 454226
rect 571584 454170 571640 454226
rect 571460 454046 571516 454102
rect 571584 454046 571640 454102
rect 571460 453922 571516 453978
rect 571584 453922 571640 453978
rect 578264 454294 578320 454350
rect 578388 454294 578444 454350
rect 578264 454170 578320 454226
rect 578388 454170 578444 454226
rect 578264 454046 578320 454102
rect 578388 454046 578444 454102
rect 578264 453922 578320 453978
rect 578388 453922 578444 453978
rect 585068 454294 585124 454350
rect 585192 454294 585248 454350
rect 585068 454170 585124 454226
rect 585192 454170 585248 454226
rect 585068 454046 585124 454102
rect 585192 454046 585248 454102
rect 585068 453922 585124 453978
rect 585192 453922 585248 453978
rect 596496 454294 596552 454350
rect 596620 454294 596676 454350
rect 596744 454294 596800 454350
rect 596868 454294 596924 454350
rect 596496 454170 596552 454226
rect 596620 454170 596676 454226
rect 596744 454170 596800 454226
rect 596868 454170 596924 454226
rect 596496 454046 596552 454102
rect 596620 454046 596676 454102
rect 596744 454046 596800 454102
rect 596868 454046 596924 454102
rect 596496 453922 596552 453978
rect 596620 453922 596676 453978
rect 596744 453922 596800 453978
rect 596868 453922 596924 453978
rect 568058 442294 568114 442350
rect 568182 442294 568238 442350
rect 568058 442170 568114 442226
rect 568182 442170 568238 442226
rect 568058 442046 568114 442102
rect 568182 442046 568238 442102
rect 568058 441922 568114 441978
rect 568182 441922 568238 441978
rect 574862 442294 574918 442350
rect 574986 442294 575042 442350
rect 574862 442170 574918 442226
rect 574986 442170 575042 442226
rect 574862 442046 574918 442102
rect 574986 442046 575042 442102
rect 574862 441922 574918 441978
rect 574986 441922 575042 441978
rect 581666 442294 581722 442350
rect 581790 442294 581846 442350
rect 581666 442170 581722 442226
rect 581790 442170 581846 442226
rect 581666 442046 581722 442102
rect 581790 442046 581846 442102
rect 581666 441922 581722 441978
rect 581790 441922 581846 441978
rect 588470 442294 588526 442350
rect 588594 442294 588650 442350
rect 588470 442170 588526 442226
rect 588594 442170 588650 442226
rect 588470 442046 588526 442102
rect 588594 442046 588650 442102
rect 588470 441922 588526 441978
rect 588594 441922 588650 441978
rect 564656 436294 564712 436350
rect 564780 436294 564836 436350
rect 564656 436170 564712 436226
rect 564780 436170 564836 436226
rect 564656 436046 564712 436102
rect 564780 436046 564836 436102
rect 564656 435922 564712 435978
rect 564780 435922 564836 435978
rect 571460 436294 571516 436350
rect 571584 436294 571640 436350
rect 571460 436170 571516 436226
rect 571584 436170 571640 436226
rect 571460 436046 571516 436102
rect 571584 436046 571640 436102
rect 571460 435922 571516 435978
rect 571584 435922 571640 435978
rect 578264 436294 578320 436350
rect 578388 436294 578444 436350
rect 578264 436170 578320 436226
rect 578388 436170 578444 436226
rect 578264 436046 578320 436102
rect 578388 436046 578444 436102
rect 578264 435922 578320 435978
rect 578388 435922 578444 435978
rect 585068 436294 585124 436350
rect 585192 436294 585248 436350
rect 585068 436170 585124 436226
rect 585192 436170 585248 436226
rect 585068 436046 585124 436102
rect 585192 436046 585248 436102
rect 585068 435922 585124 435978
rect 585192 435922 585248 435978
rect 596496 436294 596552 436350
rect 596620 436294 596676 436350
rect 596744 436294 596800 436350
rect 596868 436294 596924 436350
rect 596496 436170 596552 436226
rect 596620 436170 596676 436226
rect 596744 436170 596800 436226
rect 596868 436170 596924 436226
rect 596496 436046 596552 436102
rect 596620 436046 596676 436102
rect 596744 436046 596800 436102
rect 596868 436046 596924 436102
rect 596496 435922 596552 435978
rect 596620 435922 596676 435978
rect 596744 435922 596800 435978
rect 596868 435922 596924 435978
rect 568058 424294 568114 424350
rect 568182 424294 568238 424350
rect 568058 424170 568114 424226
rect 568182 424170 568238 424226
rect 568058 424046 568114 424102
rect 568182 424046 568238 424102
rect 568058 423922 568114 423978
rect 568182 423922 568238 423978
rect 574862 424294 574918 424350
rect 574986 424294 575042 424350
rect 574862 424170 574918 424226
rect 574986 424170 575042 424226
rect 574862 424046 574918 424102
rect 574986 424046 575042 424102
rect 574862 423922 574918 423978
rect 574986 423922 575042 423978
rect 581666 424294 581722 424350
rect 581790 424294 581846 424350
rect 581666 424170 581722 424226
rect 581790 424170 581846 424226
rect 581666 424046 581722 424102
rect 581790 424046 581846 424102
rect 581666 423922 581722 423978
rect 581790 423922 581846 423978
rect 588470 424294 588526 424350
rect 588594 424294 588650 424350
rect 588470 424170 588526 424226
rect 588594 424170 588650 424226
rect 588470 424046 588526 424102
rect 588594 424046 588650 424102
rect 588470 423922 588526 423978
rect 588594 423922 588650 423978
rect 564656 418294 564712 418350
rect 564780 418294 564836 418350
rect 564656 418170 564712 418226
rect 564780 418170 564836 418226
rect 564656 418046 564712 418102
rect 564780 418046 564836 418102
rect 564656 417922 564712 417978
rect 564780 417922 564836 417978
rect 571460 418294 571516 418350
rect 571584 418294 571640 418350
rect 571460 418170 571516 418226
rect 571584 418170 571640 418226
rect 571460 418046 571516 418102
rect 571584 418046 571640 418102
rect 571460 417922 571516 417978
rect 571584 417922 571640 417978
rect 578264 418294 578320 418350
rect 578388 418294 578444 418350
rect 578264 418170 578320 418226
rect 578388 418170 578444 418226
rect 578264 418046 578320 418102
rect 578388 418046 578444 418102
rect 578264 417922 578320 417978
rect 578388 417922 578444 417978
rect 585068 418294 585124 418350
rect 585192 418294 585248 418350
rect 585068 418170 585124 418226
rect 585192 418170 585248 418226
rect 585068 418046 585124 418102
rect 585192 418046 585248 418102
rect 585068 417922 585124 417978
rect 585192 417922 585248 417978
rect 596496 418294 596552 418350
rect 596620 418294 596676 418350
rect 596744 418294 596800 418350
rect 596868 418294 596924 418350
rect 596496 418170 596552 418226
rect 596620 418170 596676 418226
rect 596744 418170 596800 418226
rect 596868 418170 596924 418226
rect 596496 418046 596552 418102
rect 596620 418046 596676 418102
rect 596744 418046 596800 418102
rect 596868 418046 596924 418102
rect 596496 417922 596552 417978
rect 596620 417922 596676 417978
rect 596744 417922 596800 417978
rect 596868 417922 596924 417978
rect 568058 406294 568114 406350
rect 568182 406294 568238 406350
rect 568058 406170 568114 406226
rect 568182 406170 568238 406226
rect 568058 406046 568114 406102
rect 568182 406046 568238 406102
rect 568058 405922 568114 405978
rect 568182 405922 568238 405978
rect 574862 406294 574918 406350
rect 574986 406294 575042 406350
rect 574862 406170 574918 406226
rect 574986 406170 575042 406226
rect 574862 406046 574918 406102
rect 574986 406046 575042 406102
rect 574862 405922 574918 405978
rect 574986 405922 575042 405978
rect 581666 406294 581722 406350
rect 581790 406294 581846 406350
rect 581666 406170 581722 406226
rect 581790 406170 581846 406226
rect 581666 406046 581722 406102
rect 581790 406046 581846 406102
rect 581666 405922 581722 405978
rect 581790 405922 581846 405978
rect 588470 406294 588526 406350
rect 588594 406294 588650 406350
rect 588470 406170 588526 406226
rect 588594 406170 588650 406226
rect 588470 406046 588526 406102
rect 588594 406046 588650 406102
rect 588470 405922 588526 405978
rect 588594 405922 588650 405978
rect 564656 400294 564712 400350
rect 564780 400294 564836 400350
rect 564656 400170 564712 400226
rect 564780 400170 564836 400226
rect 564656 400046 564712 400102
rect 564780 400046 564836 400102
rect 564656 399922 564712 399978
rect 564780 399922 564836 399978
rect 571460 400294 571516 400350
rect 571584 400294 571640 400350
rect 571460 400170 571516 400226
rect 571584 400170 571640 400226
rect 571460 400046 571516 400102
rect 571584 400046 571640 400102
rect 571460 399922 571516 399978
rect 571584 399922 571640 399978
rect 578264 400294 578320 400350
rect 578388 400294 578444 400350
rect 578264 400170 578320 400226
rect 578388 400170 578444 400226
rect 578264 400046 578320 400102
rect 578388 400046 578444 400102
rect 578264 399922 578320 399978
rect 578388 399922 578444 399978
rect 585068 400294 585124 400350
rect 585192 400294 585248 400350
rect 585068 400170 585124 400226
rect 585192 400170 585248 400226
rect 585068 400046 585124 400102
rect 585192 400046 585248 400102
rect 585068 399922 585124 399978
rect 585192 399922 585248 399978
rect 596496 400294 596552 400350
rect 596620 400294 596676 400350
rect 596744 400294 596800 400350
rect 596868 400294 596924 400350
rect 596496 400170 596552 400226
rect 596620 400170 596676 400226
rect 596744 400170 596800 400226
rect 596868 400170 596924 400226
rect 596496 400046 596552 400102
rect 596620 400046 596676 400102
rect 596744 400046 596800 400102
rect 596868 400046 596924 400102
rect 596496 399922 596552 399978
rect 596620 399922 596676 399978
rect 596744 399922 596800 399978
rect 596868 399922 596924 399978
rect 568058 388294 568114 388350
rect 568182 388294 568238 388350
rect 568058 388170 568114 388226
rect 568182 388170 568238 388226
rect 568058 388046 568114 388102
rect 568182 388046 568238 388102
rect 568058 387922 568114 387978
rect 568182 387922 568238 387978
rect 574862 388294 574918 388350
rect 574986 388294 575042 388350
rect 574862 388170 574918 388226
rect 574986 388170 575042 388226
rect 574862 388046 574918 388102
rect 574986 388046 575042 388102
rect 574862 387922 574918 387978
rect 574986 387922 575042 387978
rect 581666 388294 581722 388350
rect 581790 388294 581846 388350
rect 581666 388170 581722 388226
rect 581790 388170 581846 388226
rect 581666 388046 581722 388102
rect 581790 388046 581846 388102
rect 581666 387922 581722 387978
rect 581790 387922 581846 387978
rect 588470 388294 588526 388350
rect 588594 388294 588650 388350
rect 588470 388170 588526 388226
rect 588594 388170 588650 388226
rect 588470 388046 588526 388102
rect 588594 388046 588650 388102
rect 588470 387922 588526 387978
rect 588594 387922 588650 387978
rect 564656 382294 564712 382350
rect 564780 382294 564836 382350
rect 564656 382170 564712 382226
rect 564780 382170 564836 382226
rect 564656 382046 564712 382102
rect 564780 382046 564836 382102
rect 564656 381922 564712 381978
rect 564780 381922 564836 381978
rect 571460 382294 571516 382350
rect 571584 382294 571640 382350
rect 571460 382170 571516 382226
rect 571584 382170 571640 382226
rect 571460 382046 571516 382102
rect 571584 382046 571640 382102
rect 571460 381922 571516 381978
rect 571584 381922 571640 381978
rect 578264 382294 578320 382350
rect 578388 382294 578444 382350
rect 578264 382170 578320 382226
rect 578388 382170 578444 382226
rect 578264 382046 578320 382102
rect 578388 382046 578444 382102
rect 578264 381922 578320 381978
rect 578388 381922 578444 381978
rect 585068 382294 585124 382350
rect 585192 382294 585248 382350
rect 585068 382170 585124 382226
rect 585192 382170 585248 382226
rect 585068 382046 585124 382102
rect 585192 382046 585248 382102
rect 585068 381922 585124 381978
rect 585192 381922 585248 381978
rect 596496 382294 596552 382350
rect 596620 382294 596676 382350
rect 596744 382294 596800 382350
rect 596868 382294 596924 382350
rect 596496 382170 596552 382226
rect 596620 382170 596676 382226
rect 596744 382170 596800 382226
rect 596868 382170 596924 382226
rect 596496 382046 596552 382102
rect 596620 382046 596676 382102
rect 596744 382046 596800 382102
rect 596868 382046 596924 382102
rect 596496 381922 596552 381978
rect 596620 381922 596676 381978
rect 596744 381922 596800 381978
rect 596868 381922 596924 381978
rect 561250 364294 561306 364350
rect 561374 364294 561430 364350
rect 561498 364294 561554 364350
rect 561622 364294 561678 364350
rect 561250 364170 561306 364226
rect 561374 364170 561430 364226
rect 561498 364170 561554 364226
rect 561622 364170 561678 364226
rect 561250 364046 561306 364102
rect 561374 364046 561430 364102
rect 561498 364046 561554 364102
rect 561622 364046 561678 364102
rect 561250 363922 561306 363978
rect 561374 363922 561430 363978
rect 561498 363922 561554 363978
rect 561622 363922 561678 363978
rect 561250 346294 561306 346350
rect 561374 346294 561430 346350
rect 561498 346294 561554 346350
rect 561622 346294 561678 346350
rect 561250 346170 561306 346226
rect 561374 346170 561430 346226
rect 561498 346170 561554 346226
rect 561622 346170 561678 346226
rect 561250 346046 561306 346102
rect 561374 346046 561430 346102
rect 561498 346046 561554 346102
rect 561622 346046 561678 346102
rect 561250 345922 561306 345978
rect 561374 345922 561430 345978
rect 561498 345922 561554 345978
rect 561622 345922 561678 345978
rect 561250 328294 561306 328350
rect 561374 328294 561430 328350
rect 561498 328294 561554 328350
rect 561622 328294 561678 328350
rect 561250 328170 561306 328226
rect 561374 328170 561430 328226
rect 561498 328170 561554 328226
rect 561622 328170 561678 328226
rect 561250 328046 561306 328102
rect 561374 328046 561430 328102
rect 561498 328046 561554 328102
rect 561622 328046 561678 328102
rect 561250 327922 561306 327978
rect 561374 327922 561430 327978
rect 561498 327922 561554 327978
rect 561622 327922 561678 327978
rect 561250 310294 561306 310350
rect 561374 310294 561430 310350
rect 561498 310294 561554 310350
rect 561622 310294 561678 310350
rect 561250 310170 561306 310226
rect 561374 310170 561430 310226
rect 561498 310170 561554 310226
rect 561622 310170 561678 310226
rect 561250 310046 561306 310102
rect 561374 310046 561430 310102
rect 561498 310046 561554 310102
rect 561622 310046 561678 310102
rect 561250 309922 561306 309978
rect 561374 309922 561430 309978
rect 561498 309922 561554 309978
rect 561622 309922 561678 309978
rect 561250 292294 561306 292350
rect 561374 292294 561430 292350
rect 561498 292294 561554 292350
rect 561622 292294 561678 292350
rect 561250 292170 561306 292226
rect 561374 292170 561430 292226
rect 561498 292170 561554 292226
rect 561622 292170 561678 292226
rect 561250 292046 561306 292102
rect 561374 292046 561430 292102
rect 561498 292046 561554 292102
rect 561622 292046 561678 292102
rect 561250 291922 561306 291978
rect 561374 291922 561430 291978
rect 561498 291922 561554 291978
rect 561622 291922 561678 291978
rect 561250 274294 561306 274350
rect 561374 274294 561430 274350
rect 561498 274294 561554 274350
rect 561622 274294 561678 274350
rect 561250 274170 561306 274226
rect 561374 274170 561430 274226
rect 561498 274170 561554 274226
rect 561622 274170 561678 274226
rect 561250 274046 561306 274102
rect 561374 274046 561430 274102
rect 561498 274046 561554 274102
rect 561622 274046 561678 274102
rect 561250 273922 561306 273978
rect 561374 273922 561430 273978
rect 561498 273922 561554 273978
rect 561622 273922 561678 273978
rect 561250 256294 561306 256350
rect 561374 256294 561430 256350
rect 561498 256294 561554 256350
rect 561622 256294 561678 256350
rect 561250 256170 561306 256226
rect 561374 256170 561430 256226
rect 561498 256170 561554 256226
rect 561622 256170 561678 256226
rect 561250 256046 561306 256102
rect 561374 256046 561430 256102
rect 561498 256046 561554 256102
rect 561622 256046 561678 256102
rect 561250 255922 561306 255978
rect 561374 255922 561430 255978
rect 561498 255922 561554 255978
rect 561622 255922 561678 255978
rect 561250 238294 561306 238350
rect 561374 238294 561430 238350
rect 561498 238294 561554 238350
rect 561622 238294 561678 238350
rect 561250 238170 561306 238226
rect 561374 238170 561430 238226
rect 561498 238170 561554 238226
rect 561622 238170 561678 238226
rect 561250 238046 561306 238102
rect 561374 238046 561430 238102
rect 561498 238046 561554 238102
rect 561622 238046 561678 238102
rect 561250 237922 561306 237978
rect 561374 237922 561430 237978
rect 561498 237922 561554 237978
rect 561622 237922 561678 237978
rect 561250 220294 561306 220350
rect 561374 220294 561430 220350
rect 561498 220294 561554 220350
rect 561622 220294 561678 220350
rect 561250 220170 561306 220226
rect 561374 220170 561430 220226
rect 561498 220170 561554 220226
rect 561622 220170 561678 220226
rect 561250 220046 561306 220102
rect 561374 220046 561430 220102
rect 561498 220046 561554 220102
rect 561622 220046 561678 220102
rect 561250 219922 561306 219978
rect 561374 219922 561430 219978
rect 561498 219922 561554 219978
rect 561622 219922 561678 219978
rect 561250 202294 561306 202350
rect 561374 202294 561430 202350
rect 561498 202294 561554 202350
rect 561622 202294 561678 202350
rect 561250 202170 561306 202226
rect 561374 202170 561430 202226
rect 561498 202170 561554 202226
rect 561622 202170 561678 202226
rect 561250 202046 561306 202102
rect 561374 202046 561430 202102
rect 561498 202046 561554 202102
rect 561622 202046 561678 202102
rect 561250 201922 561306 201978
rect 561374 201922 561430 201978
rect 561498 201922 561554 201978
rect 561622 201922 561678 201978
rect 561250 184294 561306 184350
rect 561374 184294 561430 184350
rect 561498 184294 561554 184350
rect 561622 184294 561678 184350
rect 561250 184170 561306 184226
rect 561374 184170 561430 184226
rect 561498 184170 561554 184226
rect 561622 184170 561678 184226
rect 561250 184046 561306 184102
rect 561374 184046 561430 184102
rect 561498 184046 561554 184102
rect 561622 184046 561678 184102
rect 561250 183922 561306 183978
rect 561374 183922 561430 183978
rect 561498 183922 561554 183978
rect 561622 183922 561678 183978
rect 561250 166294 561306 166350
rect 561374 166294 561430 166350
rect 561498 166294 561554 166350
rect 561622 166294 561678 166350
rect 561250 166170 561306 166226
rect 561374 166170 561430 166226
rect 561498 166170 561554 166226
rect 561622 166170 561678 166226
rect 561250 166046 561306 166102
rect 561374 166046 561430 166102
rect 561498 166046 561554 166102
rect 561622 166046 561678 166102
rect 561250 165922 561306 165978
rect 561374 165922 561430 165978
rect 561498 165922 561554 165978
rect 561622 165922 561678 165978
rect 561250 148294 561306 148350
rect 561374 148294 561430 148350
rect 561498 148294 561554 148350
rect 561622 148294 561678 148350
rect 561250 148170 561306 148226
rect 561374 148170 561430 148226
rect 561498 148170 561554 148226
rect 561622 148170 561678 148226
rect 561250 148046 561306 148102
rect 561374 148046 561430 148102
rect 561498 148046 561554 148102
rect 561622 148046 561678 148102
rect 561250 147922 561306 147978
rect 561374 147922 561430 147978
rect 561498 147922 561554 147978
rect 561622 147922 561678 147978
rect 561250 130294 561306 130350
rect 561374 130294 561430 130350
rect 561498 130294 561554 130350
rect 561622 130294 561678 130350
rect 561250 130170 561306 130226
rect 561374 130170 561430 130226
rect 561498 130170 561554 130226
rect 561622 130170 561678 130226
rect 561250 130046 561306 130102
rect 561374 130046 561430 130102
rect 561498 130046 561554 130102
rect 561622 130046 561678 130102
rect 561250 129922 561306 129978
rect 561374 129922 561430 129978
rect 561498 129922 561554 129978
rect 561622 129922 561678 129978
rect 561250 112294 561306 112350
rect 561374 112294 561430 112350
rect 561498 112294 561554 112350
rect 561622 112294 561678 112350
rect 561250 112170 561306 112226
rect 561374 112170 561430 112226
rect 561498 112170 561554 112226
rect 561622 112170 561678 112226
rect 561250 112046 561306 112102
rect 561374 112046 561430 112102
rect 561498 112046 561554 112102
rect 561622 112046 561678 112102
rect 561250 111922 561306 111978
rect 561374 111922 561430 111978
rect 561498 111922 561554 111978
rect 561622 111922 561678 111978
rect 561250 94294 561306 94350
rect 561374 94294 561430 94350
rect 561498 94294 561554 94350
rect 561622 94294 561678 94350
rect 561250 94170 561306 94226
rect 561374 94170 561430 94226
rect 561498 94170 561554 94226
rect 561622 94170 561678 94226
rect 561250 94046 561306 94102
rect 561374 94046 561430 94102
rect 561498 94046 561554 94102
rect 561622 94046 561678 94102
rect 561250 93922 561306 93978
rect 561374 93922 561430 93978
rect 561498 93922 561554 93978
rect 561622 93922 561678 93978
rect 561250 76294 561306 76350
rect 561374 76294 561430 76350
rect 561498 76294 561554 76350
rect 561622 76294 561678 76350
rect 561250 76170 561306 76226
rect 561374 76170 561430 76226
rect 561498 76170 561554 76226
rect 561622 76170 561678 76226
rect 561250 76046 561306 76102
rect 561374 76046 561430 76102
rect 561498 76046 561554 76102
rect 561622 76046 561678 76102
rect 561250 75922 561306 75978
rect 561374 75922 561430 75978
rect 561498 75922 561554 75978
rect 561622 75922 561678 75978
rect 561250 58294 561306 58350
rect 561374 58294 561430 58350
rect 561498 58294 561554 58350
rect 561622 58294 561678 58350
rect 561250 58170 561306 58226
rect 561374 58170 561430 58226
rect 561498 58170 561554 58226
rect 561622 58170 561678 58226
rect 561250 58046 561306 58102
rect 561374 58046 561430 58102
rect 561498 58046 561554 58102
rect 561622 58046 561678 58102
rect 561250 57922 561306 57978
rect 561374 57922 561430 57978
rect 561498 57922 561554 57978
rect 561622 57922 561678 57978
rect 560252 44522 560308 44578
rect 560028 39662 560084 39718
rect 560140 41102 560196 41158
rect 559804 39482 559860 39538
rect 559692 39302 559748 39358
rect 557340 37682 557396 37738
rect 560140 37862 560196 37918
rect 557788 29582 557844 29638
rect 559356 25982 559412 26038
rect 557564 25802 557620 25858
rect 557676 24362 557732 24418
rect 558022 22356 558078 22412
rect 558146 22356 558202 22412
rect 558270 22356 558326 22412
rect 558394 22356 558450 22412
rect 558518 22356 558574 22412
rect 558642 22356 558698 22412
rect 558766 22356 558822 22412
rect 558890 22356 558946 22412
rect 559014 22356 559070 22412
rect 559138 22356 559194 22412
rect 558022 22232 558078 22288
rect 558146 22232 558202 22288
rect 558270 22232 558326 22288
rect 558394 22232 558450 22288
rect 558518 22232 558574 22288
rect 558642 22232 558698 22288
rect 558766 22232 558822 22288
rect 558890 22232 558946 22288
rect 559014 22232 559070 22288
rect 559138 22232 559194 22288
rect 558022 22108 558078 22164
rect 558146 22108 558202 22164
rect 558270 22108 558326 22164
rect 558394 22108 558450 22164
rect 558518 22108 558574 22164
rect 558642 22108 558698 22164
rect 558766 22108 558822 22164
rect 558890 22108 558946 22164
rect 559014 22108 559070 22164
rect 559138 22108 559194 22164
rect 558022 21984 558078 22040
rect 558146 21984 558202 22040
rect 558270 21984 558326 22040
rect 558394 21984 558450 22040
rect 558518 21984 558574 22040
rect 558642 21984 558698 22040
rect 558766 21984 558822 22040
rect 558890 21984 558946 22040
rect 559014 21984 559070 22040
rect 559138 21984 559194 22040
rect 558022 21860 558078 21916
rect 558146 21860 558202 21916
rect 558270 21860 558326 21916
rect 558394 21860 558450 21916
rect 558518 21860 558574 21916
rect 558642 21860 558698 21916
rect 558766 21860 558822 21916
rect 558890 21860 558946 21916
rect 559014 21860 559070 21916
rect 559138 21860 559194 21916
rect 560252 25802 560308 25858
rect 561250 40294 561306 40350
rect 561374 40294 561430 40350
rect 561498 40294 561554 40350
rect 561622 40294 561678 40350
rect 561250 40170 561306 40226
rect 561374 40170 561430 40226
rect 561498 40170 561554 40226
rect 561622 40170 561678 40226
rect 561250 40046 561306 40102
rect 561374 40046 561430 40102
rect 561498 40046 561554 40102
rect 561622 40046 561678 40102
rect 561250 39922 561306 39978
rect 561374 39922 561430 39978
rect 561498 39922 561554 39978
rect 561622 39922 561678 39978
rect 561932 42722 561988 42778
rect 561932 26522 561988 26578
rect 563612 24722 563668 24778
rect 564970 370294 565026 370350
rect 565094 370294 565150 370350
rect 565218 370294 565274 370350
rect 565342 370294 565398 370350
rect 564970 370170 565026 370226
rect 565094 370170 565150 370226
rect 565218 370170 565274 370226
rect 565342 370170 565398 370226
rect 564970 370046 565026 370102
rect 565094 370046 565150 370102
rect 565218 370046 565274 370102
rect 565342 370046 565398 370102
rect 564970 369922 565026 369978
rect 565094 369922 565150 369978
rect 565218 369922 565274 369978
rect 565342 369922 565398 369978
rect 564970 352294 565026 352350
rect 565094 352294 565150 352350
rect 565218 352294 565274 352350
rect 565342 352294 565398 352350
rect 564970 352170 565026 352226
rect 565094 352170 565150 352226
rect 565218 352170 565274 352226
rect 565342 352170 565398 352226
rect 564970 352046 565026 352102
rect 565094 352046 565150 352102
rect 565218 352046 565274 352102
rect 565342 352046 565398 352102
rect 564970 351922 565026 351978
rect 565094 351922 565150 351978
rect 565218 351922 565274 351978
rect 565342 351922 565398 351978
rect 564970 334294 565026 334350
rect 565094 334294 565150 334350
rect 565218 334294 565274 334350
rect 565342 334294 565398 334350
rect 564970 334170 565026 334226
rect 565094 334170 565150 334226
rect 565218 334170 565274 334226
rect 565342 334170 565398 334226
rect 564970 334046 565026 334102
rect 565094 334046 565150 334102
rect 565218 334046 565274 334102
rect 565342 334046 565398 334102
rect 564970 333922 565026 333978
rect 565094 333922 565150 333978
rect 565218 333922 565274 333978
rect 565342 333922 565398 333978
rect 564970 316294 565026 316350
rect 565094 316294 565150 316350
rect 565218 316294 565274 316350
rect 565342 316294 565398 316350
rect 564970 316170 565026 316226
rect 565094 316170 565150 316226
rect 565218 316170 565274 316226
rect 565342 316170 565398 316226
rect 564970 316046 565026 316102
rect 565094 316046 565150 316102
rect 565218 316046 565274 316102
rect 565342 316046 565398 316102
rect 564970 315922 565026 315978
rect 565094 315922 565150 315978
rect 565218 315922 565274 315978
rect 565342 315922 565398 315978
rect 564970 298294 565026 298350
rect 565094 298294 565150 298350
rect 565218 298294 565274 298350
rect 565342 298294 565398 298350
rect 564970 298170 565026 298226
rect 565094 298170 565150 298226
rect 565218 298170 565274 298226
rect 565342 298170 565398 298226
rect 564970 298046 565026 298102
rect 565094 298046 565150 298102
rect 565218 298046 565274 298102
rect 565342 298046 565398 298102
rect 564970 297922 565026 297978
rect 565094 297922 565150 297978
rect 565218 297922 565274 297978
rect 565342 297922 565398 297978
rect 564970 280294 565026 280350
rect 565094 280294 565150 280350
rect 565218 280294 565274 280350
rect 565342 280294 565398 280350
rect 564970 280170 565026 280226
rect 565094 280170 565150 280226
rect 565218 280170 565274 280226
rect 565342 280170 565398 280226
rect 564970 280046 565026 280102
rect 565094 280046 565150 280102
rect 565218 280046 565274 280102
rect 565342 280046 565398 280102
rect 564970 279922 565026 279978
rect 565094 279922 565150 279978
rect 565218 279922 565274 279978
rect 565342 279922 565398 279978
rect 564970 262294 565026 262350
rect 565094 262294 565150 262350
rect 565218 262294 565274 262350
rect 565342 262294 565398 262350
rect 564970 262170 565026 262226
rect 565094 262170 565150 262226
rect 565218 262170 565274 262226
rect 565342 262170 565398 262226
rect 564970 262046 565026 262102
rect 565094 262046 565150 262102
rect 565218 262046 565274 262102
rect 565342 262046 565398 262102
rect 564970 261922 565026 261978
rect 565094 261922 565150 261978
rect 565218 261922 565274 261978
rect 565342 261922 565398 261978
rect 564970 244294 565026 244350
rect 565094 244294 565150 244350
rect 565218 244294 565274 244350
rect 565342 244294 565398 244350
rect 564970 244170 565026 244226
rect 565094 244170 565150 244226
rect 565218 244170 565274 244226
rect 565342 244170 565398 244226
rect 564970 244046 565026 244102
rect 565094 244046 565150 244102
rect 565218 244046 565274 244102
rect 565342 244046 565398 244102
rect 564970 243922 565026 243978
rect 565094 243922 565150 243978
rect 565218 243922 565274 243978
rect 565342 243922 565398 243978
rect 564970 226294 565026 226350
rect 565094 226294 565150 226350
rect 565218 226294 565274 226350
rect 565342 226294 565398 226350
rect 564970 226170 565026 226226
rect 565094 226170 565150 226226
rect 565218 226170 565274 226226
rect 565342 226170 565398 226226
rect 564970 226046 565026 226102
rect 565094 226046 565150 226102
rect 565218 226046 565274 226102
rect 565342 226046 565398 226102
rect 564970 225922 565026 225978
rect 565094 225922 565150 225978
rect 565218 225922 565274 225978
rect 565342 225922 565398 225978
rect 564970 208294 565026 208350
rect 565094 208294 565150 208350
rect 565218 208294 565274 208350
rect 565342 208294 565398 208350
rect 564970 208170 565026 208226
rect 565094 208170 565150 208226
rect 565218 208170 565274 208226
rect 565342 208170 565398 208226
rect 564970 208046 565026 208102
rect 565094 208046 565150 208102
rect 565218 208046 565274 208102
rect 565342 208046 565398 208102
rect 564970 207922 565026 207978
rect 565094 207922 565150 207978
rect 565218 207922 565274 207978
rect 565342 207922 565398 207978
rect 564970 190294 565026 190350
rect 565094 190294 565150 190350
rect 565218 190294 565274 190350
rect 565342 190294 565398 190350
rect 564970 190170 565026 190226
rect 565094 190170 565150 190226
rect 565218 190170 565274 190226
rect 565342 190170 565398 190226
rect 564970 190046 565026 190102
rect 565094 190046 565150 190102
rect 565218 190046 565274 190102
rect 565342 190046 565398 190102
rect 564970 189922 565026 189978
rect 565094 189922 565150 189978
rect 565218 189922 565274 189978
rect 565342 189922 565398 189978
rect 564970 172294 565026 172350
rect 565094 172294 565150 172350
rect 565218 172294 565274 172350
rect 565342 172294 565398 172350
rect 564970 172170 565026 172226
rect 565094 172170 565150 172226
rect 565218 172170 565274 172226
rect 565342 172170 565398 172226
rect 564970 172046 565026 172102
rect 565094 172046 565150 172102
rect 565218 172046 565274 172102
rect 565342 172046 565398 172102
rect 564970 171922 565026 171978
rect 565094 171922 565150 171978
rect 565218 171922 565274 171978
rect 565342 171922 565398 171978
rect 564970 154294 565026 154350
rect 565094 154294 565150 154350
rect 565218 154294 565274 154350
rect 565342 154294 565398 154350
rect 564970 154170 565026 154226
rect 565094 154170 565150 154226
rect 565218 154170 565274 154226
rect 565342 154170 565398 154226
rect 564970 154046 565026 154102
rect 565094 154046 565150 154102
rect 565218 154046 565274 154102
rect 565342 154046 565398 154102
rect 564970 153922 565026 153978
rect 565094 153922 565150 153978
rect 565218 153922 565274 153978
rect 565342 153922 565398 153978
rect 564970 136294 565026 136350
rect 565094 136294 565150 136350
rect 565218 136294 565274 136350
rect 565342 136294 565398 136350
rect 564970 136170 565026 136226
rect 565094 136170 565150 136226
rect 565218 136170 565274 136226
rect 565342 136170 565398 136226
rect 564970 136046 565026 136102
rect 565094 136046 565150 136102
rect 565218 136046 565274 136102
rect 565342 136046 565398 136102
rect 564970 135922 565026 135978
rect 565094 135922 565150 135978
rect 565218 135922 565274 135978
rect 565342 135922 565398 135978
rect 564970 118294 565026 118350
rect 565094 118294 565150 118350
rect 565218 118294 565274 118350
rect 565342 118294 565398 118350
rect 564970 118170 565026 118226
rect 565094 118170 565150 118226
rect 565218 118170 565274 118226
rect 565342 118170 565398 118226
rect 564970 118046 565026 118102
rect 565094 118046 565150 118102
rect 565218 118046 565274 118102
rect 565342 118046 565398 118102
rect 564970 117922 565026 117978
rect 565094 117922 565150 117978
rect 565218 117922 565274 117978
rect 565342 117922 565398 117978
rect 564970 100294 565026 100350
rect 565094 100294 565150 100350
rect 565218 100294 565274 100350
rect 565342 100294 565398 100350
rect 564970 100170 565026 100226
rect 565094 100170 565150 100226
rect 565218 100170 565274 100226
rect 565342 100170 565398 100226
rect 564970 100046 565026 100102
rect 565094 100046 565150 100102
rect 565218 100046 565274 100102
rect 565342 100046 565398 100102
rect 564970 99922 565026 99978
rect 565094 99922 565150 99978
rect 565218 99922 565274 99978
rect 565342 99922 565398 99978
rect 564970 82294 565026 82350
rect 565094 82294 565150 82350
rect 565218 82294 565274 82350
rect 565342 82294 565398 82350
rect 564970 82170 565026 82226
rect 565094 82170 565150 82226
rect 565218 82170 565274 82226
rect 565342 82170 565398 82226
rect 564970 82046 565026 82102
rect 565094 82046 565150 82102
rect 565218 82046 565274 82102
rect 565342 82046 565398 82102
rect 564970 81922 565026 81978
rect 565094 81922 565150 81978
rect 565218 81922 565274 81978
rect 565342 81922 565398 81978
rect 564970 64294 565026 64350
rect 565094 64294 565150 64350
rect 565218 64294 565274 64350
rect 565342 64294 565398 64350
rect 564970 64170 565026 64226
rect 565094 64170 565150 64226
rect 565218 64170 565274 64226
rect 565342 64170 565398 64226
rect 564970 64046 565026 64102
rect 565094 64046 565150 64102
rect 565218 64046 565274 64102
rect 565342 64046 565398 64102
rect 564970 63922 565026 63978
rect 565094 63922 565150 63978
rect 565218 63922 565274 63978
rect 565342 63922 565398 63978
rect 564970 46294 565026 46350
rect 565094 46294 565150 46350
rect 565218 46294 565274 46350
rect 565342 46294 565398 46350
rect 564970 46170 565026 46226
rect 565094 46170 565150 46226
rect 565218 46170 565274 46226
rect 565342 46170 565398 46226
rect 564970 46046 565026 46102
rect 565094 46046 565150 46102
rect 565218 46046 565274 46102
rect 565342 46046 565398 46102
rect 564970 45922 565026 45978
rect 565094 45922 565150 45978
rect 565218 45922 565274 45978
rect 565342 45922 565398 45978
rect 563724 25262 563780 25318
rect 561250 22294 561306 22350
rect 561374 22294 561430 22350
rect 561498 22294 561554 22350
rect 561622 22294 561678 22350
rect 561250 22170 561306 22226
rect 561374 22170 561430 22226
rect 561498 22170 561554 22226
rect 561622 22170 561678 22226
rect 561250 22046 561306 22102
rect 561374 22046 561430 22102
rect 561498 22046 561554 22102
rect 561622 22046 561678 22102
rect 561250 21922 561306 21978
rect 561374 21922 561430 21978
rect 561498 21922 561554 21978
rect 561622 21922 561678 21978
rect 565740 38582 565796 38638
rect 564970 28294 565026 28350
rect 565094 28294 565150 28350
rect 565218 28294 565274 28350
rect 565342 28294 565398 28350
rect 564970 28170 565026 28226
rect 565094 28170 565150 28226
rect 565218 28170 565274 28226
rect 565342 28170 565398 28226
rect 564970 28046 565026 28102
rect 565094 28046 565150 28102
rect 565218 28046 565274 28102
rect 565342 28046 565398 28102
rect 564970 27922 565026 27978
rect 565094 27922 565150 27978
rect 565218 27922 565274 27978
rect 565342 27922 565398 27978
rect 565628 37682 565684 37738
rect 568022 46356 568078 46412
rect 568146 46356 568202 46412
rect 568270 46356 568326 46412
rect 568394 46356 568450 46412
rect 568518 46356 568574 46412
rect 568642 46356 568698 46412
rect 568766 46356 568822 46412
rect 568890 46356 568946 46412
rect 569014 46356 569070 46412
rect 569138 46356 569194 46412
rect 568022 46232 568078 46288
rect 568146 46232 568202 46288
rect 568270 46232 568326 46288
rect 568394 46232 568450 46288
rect 568518 46232 568574 46288
rect 568642 46232 568698 46288
rect 568766 46232 568822 46288
rect 568890 46232 568946 46288
rect 569014 46232 569070 46288
rect 569138 46232 569194 46288
rect 568022 46108 568078 46164
rect 568146 46108 568202 46164
rect 568270 46108 568326 46164
rect 568394 46108 568450 46164
rect 568518 46108 568574 46164
rect 568642 46108 568698 46164
rect 568766 46108 568822 46164
rect 568890 46108 568946 46164
rect 569014 46108 569070 46164
rect 569138 46108 569194 46164
rect 568022 45984 568078 46040
rect 568146 45984 568202 46040
rect 568270 45984 568326 46040
rect 568394 45984 568450 46040
rect 568518 45984 568574 46040
rect 568642 45984 568698 46040
rect 568766 45984 568822 46040
rect 568890 45984 568946 46040
rect 569014 45984 569070 46040
rect 569138 45984 569194 46040
rect 568022 45860 568078 45916
rect 568146 45860 568202 45916
rect 568270 45860 568326 45916
rect 568394 45860 568450 45916
rect 568518 45860 568574 45916
rect 568642 45860 568698 45916
rect 568766 45860 568822 45916
rect 568890 45860 568946 45916
rect 569014 45860 569070 45916
rect 569138 45860 569194 45916
rect 566972 36782 567028 36838
rect 567756 42902 567812 42958
rect 565740 29402 565796 29458
rect 565628 25982 565684 26038
rect 568022 28356 568078 28412
rect 568146 28356 568202 28412
rect 568270 28356 568326 28412
rect 568394 28356 568450 28412
rect 568518 28356 568574 28412
rect 568642 28356 568698 28412
rect 568766 28356 568822 28412
rect 568890 28356 568946 28412
rect 569014 28356 569070 28412
rect 569138 28356 569194 28412
rect 568022 28232 568078 28288
rect 568146 28232 568202 28288
rect 568270 28232 568326 28288
rect 568394 28232 568450 28288
rect 568518 28232 568574 28288
rect 568642 28232 568698 28288
rect 568766 28232 568822 28288
rect 568890 28232 568946 28288
rect 569014 28232 569070 28288
rect 569138 28232 569194 28288
rect 568022 28108 568078 28164
rect 568146 28108 568202 28164
rect 568270 28108 568326 28164
rect 568394 28108 568450 28164
rect 568518 28108 568574 28164
rect 568642 28108 568698 28164
rect 568766 28108 568822 28164
rect 568890 28108 568946 28164
rect 569014 28108 569070 28164
rect 569138 28108 569194 28164
rect 568022 27984 568078 28040
rect 568146 27984 568202 28040
rect 568270 27984 568326 28040
rect 568394 27984 568450 28040
rect 568518 27984 568574 28040
rect 568642 27984 568698 28040
rect 568766 27984 568822 28040
rect 568890 27984 568946 28040
rect 569014 27984 569070 28040
rect 569138 27984 569194 28040
rect 568022 27860 568078 27916
rect 568146 27860 568202 27916
rect 568270 27860 568326 27916
rect 568394 27860 568450 27916
rect 568518 27860 568574 27916
rect 568642 27860 568698 27916
rect 568766 27860 568822 27916
rect 568890 27860 568946 27916
rect 569014 27860 569070 27916
rect 569138 27860 569194 27916
rect 567756 24902 567812 24958
rect 563724 20042 563780 20098
rect 560028 13022 560084 13078
rect 546970 -1176 547026 -1120
rect 547094 -1176 547150 -1120
rect 547218 -1176 547274 -1120
rect 547342 -1176 547398 -1120
rect 546970 -1300 547026 -1244
rect 547094 -1300 547150 -1244
rect 547218 -1300 547274 -1244
rect 547342 -1300 547398 -1244
rect 546970 -1424 547026 -1368
rect 547094 -1424 547150 -1368
rect 547218 -1424 547274 -1368
rect 547342 -1424 547398 -1368
rect 546970 -1548 547026 -1492
rect 547094 -1548 547150 -1492
rect 547218 -1548 547274 -1492
rect 547342 -1548 547398 -1492
rect 561250 4294 561306 4350
rect 561374 4294 561430 4350
rect 561498 4294 561554 4350
rect 561622 4294 561678 4350
rect 561250 4170 561306 4226
rect 561374 4170 561430 4226
rect 561498 4170 561554 4226
rect 561622 4170 561678 4226
rect 561250 4046 561306 4102
rect 561374 4046 561430 4102
rect 561498 4046 561554 4102
rect 561622 4046 561678 4102
rect 561250 3922 561306 3978
rect 561374 3922 561430 3978
rect 561498 3922 561554 3978
rect 561622 3922 561678 3978
rect 561250 -216 561306 -160
rect 561374 -216 561430 -160
rect 561498 -216 561554 -160
rect 561622 -216 561678 -160
rect 561250 -340 561306 -284
rect 561374 -340 561430 -284
rect 561498 -340 561554 -284
rect 561622 -340 561678 -284
rect 561250 -464 561306 -408
rect 561374 -464 561430 -408
rect 561498 -464 561554 -408
rect 561622 -464 561678 -408
rect 561250 -588 561306 -532
rect 561374 -588 561430 -532
rect 561498 -588 561554 -532
rect 561622 -588 561678 -532
rect 564970 10294 565026 10350
rect 565094 10294 565150 10350
rect 565218 10294 565274 10350
rect 565342 10294 565398 10350
rect 564970 10170 565026 10226
rect 565094 10170 565150 10226
rect 565218 10170 565274 10226
rect 565342 10170 565398 10226
rect 564970 10046 565026 10102
rect 565094 10046 565150 10102
rect 565218 10046 565274 10102
rect 565342 10046 565398 10102
rect 564970 9922 565026 9978
rect 565094 9922 565150 9978
rect 565218 9922 565274 9978
rect 565342 9922 565398 9978
rect 570108 24902 570164 24958
rect 571004 7442 571060 7498
rect 572572 7802 572628 7858
rect 572684 7622 572740 7678
rect 572908 36962 572964 37018
rect 572796 7982 572852 8038
rect 573692 38582 573748 38638
rect 579250 364294 579306 364350
rect 579374 364294 579430 364350
rect 579498 364294 579554 364350
rect 579622 364294 579678 364350
rect 579250 364170 579306 364226
rect 579374 364170 579430 364226
rect 579498 364170 579554 364226
rect 579622 364170 579678 364226
rect 579250 364046 579306 364102
rect 579374 364046 579430 364102
rect 579498 364046 579554 364102
rect 579622 364046 579678 364102
rect 579250 363922 579306 363978
rect 579374 363922 579430 363978
rect 579498 363922 579554 363978
rect 579622 363922 579678 363978
rect 579250 346294 579306 346350
rect 579374 346294 579430 346350
rect 579498 346294 579554 346350
rect 579622 346294 579678 346350
rect 579250 346170 579306 346226
rect 579374 346170 579430 346226
rect 579498 346170 579554 346226
rect 579622 346170 579678 346226
rect 579250 346046 579306 346102
rect 579374 346046 579430 346102
rect 579498 346046 579554 346102
rect 579622 346046 579678 346102
rect 579250 345922 579306 345978
rect 579374 345922 579430 345978
rect 579498 345922 579554 345978
rect 579622 345922 579678 345978
rect 579250 328294 579306 328350
rect 579374 328294 579430 328350
rect 579498 328294 579554 328350
rect 579622 328294 579678 328350
rect 579250 328170 579306 328226
rect 579374 328170 579430 328226
rect 579498 328170 579554 328226
rect 579622 328170 579678 328226
rect 579250 328046 579306 328102
rect 579374 328046 579430 328102
rect 579498 328046 579554 328102
rect 579622 328046 579678 328102
rect 579250 327922 579306 327978
rect 579374 327922 579430 327978
rect 579498 327922 579554 327978
rect 579622 327922 579678 327978
rect 579250 310294 579306 310350
rect 579374 310294 579430 310350
rect 579498 310294 579554 310350
rect 579622 310294 579678 310350
rect 579250 310170 579306 310226
rect 579374 310170 579430 310226
rect 579498 310170 579554 310226
rect 579622 310170 579678 310226
rect 579250 310046 579306 310102
rect 579374 310046 579430 310102
rect 579498 310046 579554 310102
rect 579622 310046 579678 310102
rect 579250 309922 579306 309978
rect 579374 309922 579430 309978
rect 579498 309922 579554 309978
rect 579622 309922 579678 309978
rect 579250 292294 579306 292350
rect 579374 292294 579430 292350
rect 579498 292294 579554 292350
rect 579622 292294 579678 292350
rect 579250 292170 579306 292226
rect 579374 292170 579430 292226
rect 579498 292170 579554 292226
rect 579622 292170 579678 292226
rect 579250 292046 579306 292102
rect 579374 292046 579430 292102
rect 579498 292046 579554 292102
rect 579622 292046 579678 292102
rect 579250 291922 579306 291978
rect 579374 291922 579430 291978
rect 579498 291922 579554 291978
rect 579622 291922 579678 291978
rect 579250 274294 579306 274350
rect 579374 274294 579430 274350
rect 579498 274294 579554 274350
rect 579622 274294 579678 274350
rect 579250 274170 579306 274226
rect 579374 274170 579430 274226
rect 579498 274170 579554 274226
rect 579622 274170 579678 274226
rect 579250 274046 579306 274102
rect 579374 274046 579430 274102
rect 579498 274046 579554 274102
rect 579622 274046 579678 274102
rect 579250 273922 579306 273978
rect 579374 273922 579430 273978
rect 579498 273922 579554 273978
rect 579622 273922 579678 273978
rect 579250 256294 579306 256350
rect 579374 256294 579430 256350
rect 579498 256294 579554 256350
rect 579622 256294 579678 256350
rect 579250 256170 579306 256226
rect 579374 256170 579430 256226
rect 579498 256170 579554 256226
rect 579622 256170 579678 256226
rect 579250 256046 579306 256102
rect 579374 256046 579430 256102
rect 579498 256046 579554 256102
rect 579622 256046 579678 256102
rect 579250 255922 579306 255978
rect 579374 255922 579430 255978
rect 579498 255922 579554 255978
rect 579622 255922 579678 255978
rect 579250 238294 579306 238350
rect 579374 238294 579430 238350
rect 579498 238294 579554 238350
rect 579622 238294 579678 238350
rect 579250 238170 579306 238226
rect 579374 238170 579430 238226
rect 579498 238170 579554 238226
rect 579622 238170 579678 238226
rect 579250 238046 579306 238102
rect 579374 238046 579430 238102
rect 579498 238046 579554 238102
rect 579622 238046 579678 238102
rect 579250 237922 579306 237978
rect 579374 237922 579430 237978
rect 579498 237922 579554 237978
rect 579622 237922 579678 237978
rect 579250 220294 579306 220350
rect 579374 220294 579430 220350
rect 579498 220294 579554 220350
rect 579622 220294 579678 220350
rect 579250 220170 579306 220226
rect 579374 220170 579430 220226
rect 579498 220170 579554 220226
rect 579622 220170 579678 220226
rect 579250 220046 579306 220102
rect 579374 220046 579430 220102
rect 579498 220046 579554 220102
rect 579622 220046 579678 220102
rect 579250 219922 579306 219978
rect 579374 219922 579430 219978
rect 579498 219922 579554 219978
rect 579622 219922 579678 219978
rect 579250 202294 579306 202350
rect 579374 202294 579430 202350
rect 579498 202294 579554 202350
rect 579622 202294 579678 202350
rect 579250 202170 579306 202226
rect 579374 202170 579430 202226
rect 579498 202170 579554 202226
rect 579622 202170 579678 202226
rect 579250 202046 579306 202102
rect 579374 202046 579430 202102
rect 579498 202046 579554 202102
rect 579622 202046 579678 202102
rect 579250 201922 579306 201978
rect 579374 201922 579430 201978
rect 579498 201922 579554 201978
rect 579622 201922 579678 201978
rect 579250 184294 579306 184350
rect 579374 184294 579430 184350
rect 579498 184294 579554 184350
rect 579622 184294 579678 184350
rect 579250 184170 579306 184226
rect 579374 184170 579430 184226
rect 579498 184170 579554 184226
rect 579622 184170 579678 184226
rect 579250 184046 579306 184102
rect 579374 184046 579430 184102
rect 579498 184046 579554 184102
rect 579622 184046 579678 184102
rect 579250 183922 579306 183978
rect 579374 183922 579430 183978
rect 579498 183922 579554 183978
rect 579622 183922 579678 183978
rect 579250 166294 579306 166350
rect 579374 166294 579430 166350
rect 579498 166294 579554 166350
rect 579622 166294 579678 166350
rect 579250 166170 579306 166226
rect 579374 166170 579430 166226
rect 579498 166170 579554 166226
rect 579622 166170 579678 166226
rect 579250 166046 579306 166102
rect 579374 166046 579430 166102
rect 579498 166046 579554 166102
rect 579622 166046 579678 166102
rect 579250 165922 579306 165978
rect 579374 165922 579430 165978
rect 579498 165922 579554 165978
rect 579622 165922 579678 165978
rect 579250 148294 579306 148350
rect 579374 148294 579430 148350
rect 579498 148294 579554 148350
rect 579622 148294 579678 148350
rect 579250 148170 579306 148226
rect 579374 148170 579430 148226
rect 579498 148170 579554 148226
rect 579622 148170 579678 148226
rect 579250 148046 579306 148102
rect 579374 148046 579430 148102
rect 579498 148046 579554 148102
rect 579622 148046 579678 148102
rect 579250 147922 579306 147978
rect 579374 147922 579430 147978
rect 579498 147922 579554 147978
rect 579622 147922 579678 147978
rect 579250 130294 579306 130350
rect 579374 130294 579430 130350
rect 579498 130294 579554 130350
rect 579622 130294 579678 130350
rect 579250 130170 579306 130226
rect 579374 130170 579430 130226
rect 579498 130170 579554 130226
rect 579622 130170 579678 130226
rect 579250 130046 579306 130102
rect 579374 130046 579430 130102
rect 579498 130046 579554 130102
rect 579622 130046 579678 130102
rect 579250 129922 579306 129978
rect 579374 129922 579430 129978
rect 579498 129922 579554 129978
rect 579622 129922 579678 129978
rect 579250 112294 579306 112350
rect 579374 112294 579430 112350
rect 579498 112294 579554 112350
rect 579622 112294 579678 112350
rect 579250 112170 579306 112226
rect 579374 112170 579430 112226
rect 579498 112170 579554 112226
rect 579622 112170 579678 112226
rect 579250 112046 579306 112102
rect 579374 112046 579430 112102
rect 579498 112046 579554 112102
rect 579622 112046 579678 112102
rect 579250 111922 579306 111978
rect 579374 111922 579430 111978
rect 579498 111922 579554 111978
rect 579622 111922 579678 111978
rect 579250 94294 579306 94350
rect 579374 94294 579430 94350
rect 579498 94294 579554 94350
rect 579622 94294 579678 94350
rect 579250 94170 579306 94226
rect 579374 94170 579430 94226
rect 579498 94170 579554 94226
rect 579622 94170 579678 94226
rect 579250 94046 579306 94102
rect 579374 94046 579430 94102
rect 579498 94046 579554 94102
rect 579622 94046 579678 94102
rect 579250 93922 579306 93978
rect 579374 93922 579430 93978
rect 579498 93922 579554 93978
rect 579622 93922 579678 93978
rect 579250 76294 579306 76350
rect 579374 76294 579430 76350
rect 579498 76294 579554 76350
rect 579622 76294 579678 76350
rect 579250 76170 579306 76226
rect 579374 76170 579430 76226
rect 579498 76170 579554 76226
rect 579622 76170 579678 76226
rect 579250 76046 579306 76102
rect 579374 76046 579430 76102
rect 579498 76046 579554 76102
rect 579622 76046 579678 76102
rect 579250 75922 579306 75978
rect 579374 75922 579430 75978
rect 579498 75922 579554 75978
rect 579622 75922 579678 75978
rect 577052 42902 577108 42958
rect 578022 40356 578078 40412
rect 578146 40356 578202 40412
rect 578270 40356 578326 40412
rect 578394 40356 578450 40412
rect 578518 40356 578574 40412
rect 578642 40356 578698 40412
rect 578766 40356 578822 40412
rect 578890 40356 578946 40412
rect 579014 40356 579070 40412
rect 579138 40356 579194 40412
rect 578022 40232 578078 40288
rect 578146 40232 578202 40288
rect 578270 40232 578326 40288
rect 578394 40232 578450 40288
rect 578518 40232 578574 40288
rect 578642 40232 578698 40288
rect 578766 40232 578822 40288
rect 578890 40232 578946 40288
rect 579014 40232 579070 40288
rect 579138 40232 579194 40288
rect 578022 40108 578078 40164
rect 578146 40108 578202 40164
rect 578270 40108 578326 40164
rect 578394 40108 578450 40164
rect 578518 40108 578574 40164
rect 578642 40108 578698 40164
rect 578766 40108 578822 40164
rect 578890 40108 578946 40164
rect 579014 40108 579070 40164
rect 579138 40108 579194 40164
rect 578022 39984 578078 40040
rect 578146 39984 578202 40040
rect 578270 39984 578326 40040
rect 578394 39984 578450 40040
rect 578518 39984 578574 40040
rect 578642 39984 578698 40040
rect 578766 39984 578822 40040
rect 578890 39984 578946 40040
rect 579014 39984 579070 40040
rect 579138 39984 579194 40040
rect 578022 39860 578078 39916
rect 578146 39860 578202 39916
rect 578270 39860 578326 39916
rect 578394 39860 578450 39916
rect 578518 39860 578574 39916
rect 578642 39860 578698 39916
rect 578766 39860 578822 39916
rect 578890 39860 578946 39916
rect 579014 39860 579070 39916
rect 579138 39860 579194 39916
rect 577164 36962 577220 37018
rect 577052 25262 577108 25318
rect 578022 22356 578078 22412
rect 578146 22356 578202 22412
rect 578270 22356 578326 22412
rect 578394 22356 578450 22412
rect 578518 22356 578574 22412
rect 578642 22356 578698 22412
rect 578766 22356 578822 22412
rect 578890 22356 578946 22412
rect 579014 22356 579070 22412
rect 579138 22356 579194 22412
rect 578022 22232 578078 22288
rect 578146 22232 578202 22288
rect 578270 22232 578326 22288
rect 578394 22232 578450 22288
rect 578518 22232 578574 22288
rect 578642 22232 578698 22288
rect 578766 22232 578822 22288
rect 578890 22232 578946 22288
rect 579014 22232 579070 22288
rect 579138 22232 579194 22288
rect 578022 22108 578078 22164
rect 578146 22108 578202 22164
rect 578270 22108 578326 22164
rect 578394 22108 578450 22164
rect 578518 22108 578574 22164
rect 578642 22108 578698 22164
rect 578766 22108 578822 22164
rect 578890 22108 578946 22164
rect 579014 22108 579070 22164
rect 579138 22108 579194 22164
rect 578022 21984 578078 22040
rect 578146 21984 578202 22040
rect 578270 21984 578326 22040
rect 578394 21984 578450 22040
rect 578518 21984 578574 22040
rect 578642 21984 578698 22040
rect 578766 21984 578822 22040
rect 578890 21984 578946 22040
rect 579014 21984 579070 22040
rect 579138 21984 579194 22040
rect 578022 21860 578078 21916
rect 578146 21860 578202 21916
rect 578270 21860 578326 21916
rect 578394 21860 578450 21916
rect 578518 21860 578574 21916
rect 578642 21860 578698 21916
rect 578766 21860 578822 21916
rect 578890 21860 578946 21916
rect 579014 21860 579070 21916
rect 579138 21860 579194 21916
rect 577052 7982 577108 8038
rect 577948 7802 578004 7858
rect 578844 7622 578900 7678
rect 582092 44522 582148 44578
rect 582970 370294 583026 370350
rect 583094 370294 583150 370350
rect 583218 370294 583274 370350
rect 583342 370294 583398 370350
rect 582970 370170 583026 370226
rect 583094 370170 583150 370226
rect 583218 370170 583274 370226
rect 583342 370170 583398 370226
rect 582970 370046 583026 370102
rect 583094 370046 583150 370102
rect 583218 370046 583274 370102
rect 583342 370046 583398 370102
rect 582970 369922 583026 369978
rect 583094 369922 583150 369978
rect 583218 369922 583274 369978
rect 583342 369922 583398 369978
rect 582970 352294 583026 352350
rect 583094 352294 583150 352350
rect 583218 352294 583274 352350
rect 583342 352294 583398 352350
rect 582970 352170 583026 352226
rect 583094 352170 583150 352226
rect 583218 352170 583274 352226
rect 583342 352170 583398 352226
rect 582970 352046 583026 352102
rect 583094 352046 583150 352102
rect 583218 352046 583274 352102
rect 583342 352046 583398 352102
rect 582970 351922 583026 351978
rect 583094 351922 583150 351978
rect 583218 351922 583274 351978
rect 583342 351922 583398 351978
rect 582970 334294 583026 334350
rect 583094 334294 583150 334350
rect 583218 334294 583274 334350
rect 583342 334294 583398 334350
rect 582970 334170 583026 334226
rect 583094 334170 583150 334226
rect 583218 334170 583274 334226
rect 583342 334170 583398 334226
rect 582970 334046 583026 334102
rect 583094 334046 583150 334102
rect 583218 334046 583274 334102
rect 583342 334046 583398 334102
rect 582970 333922 583026 333978
rect 583094 333922 583150 333978
rect 583218 333922 583274 333978
rect 583342 333922 583398 333978
rect 582970 316294 583026 316350
rect 583094 316294 583150 316350
rect 583218 316294 583274 316350
rect 583342 316294 583398 316350
rect 582970 316170 583026 316226
rect 583094 316170 583150 316226
rect 583218 316170 583274 316226
rect 583342 316170 583398 316226
rect 582970 316046 583026 316102
rect 583094 316046 583150 316102
rect 583218 316046 583274 316102
rect 583342 316046 583398 316102
rect 582970 315922 583026 315978
rect 583094 315922 583150 315978
rect 583218 315922 583274 315978
rect 583342 315922 583398 315978
rect 582970 298294 583026 298350
rect 583094 298294 583150 298350
rect 583218 298294 583274 298350
rect 583342 298294 583398 298350
rect 582970 298170 583026 298226
rect 583094 298170 583150 298226
rect 583218 298170 583274 298226
rect 583342 298170 583398 298226
rect 582970 298046 583026 298102
rect 583094 298046 583150 298102
rect 583218 298046 583274 298102
rect 583342 298046 583398 298102
rect 582970 297922 583026 297978
rect 583094 297922 583150 297978
rect 583218 297922 583274 297978
rect 583342 297922 583398 297978
rect 582970 280294 583026 280350
rect 583094 280294 583150 280350
rect 583218 280294 583274 280350
rect 583342 280294 583398 280350
rect 582970 280170 583026 280226
rect 583094 280170 583150 280226
rect 583218 280170 583274 280226
rect 583342 280170 583398 280226
rect 582970 280046 583026 280102
rect 583094 280046 583150 280102
rect 583218 280046 583274 280102
rect 583342 280046 583398 280102
rect 582970 279922 583026 279978
rect 583094 279922 583150 279978
rect 583218 279922 583274 279978
rect 583342 279922 583398 279978
rect 582970 262294 583026 262350
rect 583094 262294 583150 262350
rect 583218 262294 583274 262350
rect 583342 262294 583398 262350
rect 582970 262170 583026 262226
rect 583094 262170 583150 262226
rect 583218 262170 583274 262226
rect 583342 262170 583398 262226
rect 582970 262046 583026 262102
rect 583094 262046 583150 262102
rect 583218 262046 583274 262102
rect 583342 262046 583398 262102
rect 582970 261922 583026 261978
rect 583094 261922 583150 261978
rect 583218 261922 583274 261978
rect 583342 261922 583398 261978
rect 582970 244294 583026 244350
rect 583094 244294 583150 244350
rect 583218 244294 583274 244350
rect 583342 244294 583398 244350
rect 582970 244170 583026 244226
rect 583094 244170 583150 244226
rect 583218 244170 583274 244226
rect 583342 244170 583398 244226
rect 582970 244046 583026 244102
rect 583094 244046 583150 244102
rect 583218 244046 583274 244102
rect 583342 244046 583398 244102
rect 582970 243922 583026 243978
rect 583094 243922 583150 243978
rect 583218 243922 583274 243978
rect 583342 243922 583398 243978
rect 582970 226294 583026 226350
rect 583094 226294 583150 226350
rect 583218 226294 583274 226350
rect 583342 226294 583398 226350
rect 582970 226170 583026 226226
rect 583094 226170 583150 226226
rect 583218 226170 583274 226226
rect 583342 226170 583398 226226
rect 582970 226046 583026 226102
rect 583094 226046 583150 226102
rect 583218 226046 583274 226102
rect 583342 226046 583398 226102
rect 582970 225922 583026 225978
rect 583094 225922 583150 225978
rect 583218 225922 583274 225978
rect 583342 225922 583398 225978
rect 582970 208294 583026 208350
rect 583094 208294 583150 208350
rect 583218 208294 583274 208350
rect 583342 208294 583398 208350
rect 582970 208170 583026 208226
rect 583094 208170 583150 208226
rect 583218 208170 583274 208226
rect 583342 208170 583398 208226
rect 582970 208046 583026 208102
rect 583094 208046 583150 208102
rect 583218 208046 583274 208102
rect 583342 208046 583398 208102
rect 582970 207922 583026 207978
rect 583094 207922 583150 207978
rect 583218 207922 583274 207978
rect 583342 207922 583398 207978
rect 582970 190294 583026 190350
rect 583094 190294 583150 190350
rect 583218 190294 583274 190350
rect 583342 190294 583398 190350
rect 582970 190170 583026 190226
rect 583094 190170 583150 190226
rect 583218 190170 583274 190226
rect 583342 190170 583398 190226
rect 582970 190046 583026 190102
rect 583094 190046 583150 190102
rect 583218 190046 583274 190102
rect 583342 190046 583398 190102
rect 582970 189922 583026 189978
rect 583094 189922 583150 189978
rect 583218 189922 583274 189978
rect 583342 189922 583398 189978
rect 582970 172294 583026 172350
rect 583094 172294 583150 172350
rect 583218 172294 583274 172350
rect 583342 172294 583398 172350
rect 582970 172170 583026 172226
rect 583094 172170 583150 172226
rect 583218 172170 583274 172226
rect 583342 172170 583398 172226
rect 582970 172046 583026 172102
rect 583094 172046 583150 172102
rect 583218 172046 583274 172102
rect 583342 172046 583398 172102
rect 582970 171922 583026 171978
rect 583094 171922 583150 171978
rect 583218 171922 583274 171978
rect 583342 171922 583398 171978
rect 582970 154294 583026 154350
rect 583094 154294 583150 154350
rect 583218 154294 583274 154350
rect 583342 154294 583398 154350
rect 582970 154170 583026 154226
rect 583094 154170 583150 154226
rect 583218 154170 583274 154226
rect 583342 154170 583398 154226
rect 582970 154046 583026 154102
rect 583094 154046 583150 154102
rect 583218 154046 583274 154102
rect 583342 154046 583398 154102
rect 582970 153922 583026 153978
rect 583094 153922 583150 153978
rect 583218 153922 583274 153978
rect 583342 153922 583398 153978
rect 582970 136294 583026 136350
rect 583094 136294 583150 136350
rect 583218 136294 583274 136350
rect 583342 136294 583398 136350
rect 582970 136170 583026 136226
rect 583094 136170 583150 136226
rect 583218 136170 583274 136226
rect 583342 136170 583398 136226
rect 582970 136046 583026 136102
rect 583094 136046 583150 136102
rect 583218 136046 583274 136102
rect 583342 136046 583398 136102
rect 582970 135922 583026 135978
rect 583094 135922 583150 135978
rect 583218 135922 583274 135978
rect 583342 135922 583398 135978
rect 582970 118294 583026 118350
rect 583094 118294 583150 118350
rect 583218 118294 583274 118350
rect 583342 118294 583398 118350
rect 582970 118170 583026 118226
rect 583094 118170 583150 118226
rect 583218 118170 583274 118226
rect 583342 118170 583398 118226
rect 582970 118046 583026 118102
rect 583094 118046 583150 118102
rect 583218 118046 583274 118102
rect 583342 118046 583398 118102
rect 582970 117922 583026 117978
rect 583094 117922 583150 117978
rect 583218 117922 583274 117978
rect 583342 117922 583398 117978
rect 582970 100294 583026 100350
rect 583094 100294 583150 100350
rect 583218 100294 583274 100350
rect 583342 100294 583398 100350
rect 582970 100170 583026 100226
rect 583094 100170 583150 100226
rect 583218 100170 583274 100226
rect 583342 100170 583398 100226
rect 582970 100046 583026 100102
rect 583094 100046 583150 100102
rect 583218 100046 583274 100102
rect 583342 100046 583398 100102
rect 582970 99922 583026 99978
rect 583094 99922 583150 99978
rect 583218 99922 583274 99978
rect 583342 99922 583398 99978
rect 582970 82294 583026 82350
rect 583094 82294 583150 82350
rect 583218 82294 583274 82350
rect 583342 82294 583398 82350
rect 582970 82170 583026 82226
rect 583094 82170 583150 82226
rect 583218 82170 583274 82226
rect 583342 82170 583398 82226
rect 582970 82046 583026 82102
rect 583094 82046 583150 82102
rect 583218 82046 583274 82102
rect 583342 82046 583398 82102
rect 582970 81922 583026 81978
rect 583094 81922 583150 81978
rect 583218 81922 583274 81978
rect 583342 81922 583398 81978
rect 582970 64294 583026 64350
rect 583094 64294 583150 64350
rect 583218 64294 583274 64350
rect 583342 64294 583398 64350
rect 582970 64170 583026 64226
rect 583094 64170 583150 64226
rect 583218 64170 583274 64226
rect 583342 64170 583398 64226
rect 582970 64046 583026 64102
rect 583094 64046 583150 64102
rect 583218 64046 583274 64102
rect 583342 64046 583398 64102
rect 582970 63922 583026 63978
rect 583094 63922 583150 63978
rect 583218 63922 583274 63978
rect 583342 63922 583398 63978
rect 582970 46294 583026 46350
rect 583094 46294 583150 46350
rect 583218 46294 583274 46350
rect 583342 46294 583398 46350
rect 582970 46170 583026 46226
rect 583094 46170 583150 46226
rect 583218 46170 583274 46226
rect 583342 46170 583398 46226
rect 582970 46046 583026 46102
rect 583094 46046 583150 46102
rect 583218 46046 583274 46102
rect 583342 46046 583398 46102
rect 582970 45922 583026 45978
rect 583094 45922 583150 45978
rect 583218 45922 583274 45978
rect 583342 45922 583398 45978
rect 581420 37682 581476 37738
rect 582970 28294 583026 28350
rect 583094 28294 583150 28350
rect 583218 28294 583274 28350
rect 583342 28294 583398 28350
rect 582970 28170 583026 28226
rect 583094 28170 583150 28226
rect 583218 28170 583274 28226
rect 583342 28170 583398 28226
rect 582970 28046 583026 28102
rect 583094 28046 583150 28102
rect 583218 28046 583274 28102
rect 583342 28046 583398 28102
rect 582970 27922 583026 27978
rect 583094 27922 583150 27978
rect 583218 27922 583274 27978
rect 583342 27922 583398 27978
rect 582970 10294 583026 10350
rect 583094 10294 583150 10350
rect 583218 10294 583274 10350
rect 583342 10294 583398 10350
rect 582970 10170 583026 10226
rect 583094 10170 583150 10226
rect 583218 10170 583274 10226
rect 583342 10170 583398 10226
rect 582970 10046 583026 10102
rect 583094 10046 583150 10102
rect 583218 10046 583274 10102
rect 583342 10046 583398 10102
rect 582970 9922 583026 9978
rect 583094 9922 583150 9978
rect 583218 9922 583274 9978
rect 583342 9922 583398 9978
rect 579852 7442 579908 7498
rect 579250 4294 579306 4350
rect 579374 4294 579430 4350
rect 579498 4294 579554 4350
rect 579622 4294 579678 4350
rect 579250 4170 579306 4226
rect 579374 4170 579430 4226
rect 579498 4170 579554 4226
rect 579622 4170 579678 4226
rect 579250 4046 579306 4102
rect 579374 4046 579430 4102
rect 579498 4046 579554 4102
rect 579622 4046 579678 4102
rect 579250 3922 579306 3978
rect 579374 3922 579430 3978
rect 579498 3922 579554 3978
rect 579622 3922 579678 3978
rect 564970 -1176 565026 -1120
rect 565094 -1176 565150 -1120
rect 565218 -1176 565274 -1120
rect 565342 -1176 565398 -1120
rect 564970 -1300 565026 -1244
rect 565094 -1300 565150 -1244
rect 565218 -1300 565274 -1244
rect 565342 -1300 565398 -1244
rect 564970 -1424 565026 -1368
rect 565094 -1424 565150 -1368
rect 565218 -1424 565274 -1368
rect 565342 -1424 565398 -1368
rect 564970 -1548 565026 -1492
rect 565094 -1548 565150 -1492
rect 565218 -1548 565274 -1492
rect 565342 -1548 565398 -1492
rect 579250 -216 579306 -160
rect 579374 -216 579430 -160
rect 579498 -216 579554 -160
rect 579622 -216 579678 -160
rect 579250 -340 579306 -284
rect 579374 -340 579430 -284
rect 579498 -340 579554 -284
rect 579622 -340 579678 -284
rect 579250 -464 579306 -408
rect 579374 -464 579430 -408
rect 579498 -464 579554 -408
rect 579622 -464 579678 -408
rect 579250 -588 579306 -532
rect 579374 -588 579430 -532
rect 579498 -588 579554 -532
rect 579622 -588 579678 -532
rect 584892 47762 584948 47818
rect 584780 41102 584836 41158
rect 586012 10682 586068 10738
rect 596496 364294 596552 364350
rect 596620 364294 596676 364350
rect 596744 364294 596800 364350
rect 596868 364294 596924 364350
rect 596496 364170 596552 364226
rect 596620 364170 596676 364226
rect 596744 364170 596800 364226
rect 596868 364170 596924 364226
rect 596496 364046 596552 364102
rect 596620 364046 596676 364102
rect 596744 364046 596800 364102
rect 596868 364046 596924 364102
rect 596496 363922 596552 363978
rect 596620 363922 596676 363978
rect 596744 363922 596800 363978
rect 596868 363922 596924 363978
rect 596496 346294 596552 346350
rect 596620 346294 596676 346350
rect 596744 346294 596800 346350
rect 596868 346294 596924 346350
rect 596496 346170 596552 346226
rect 596620 346170 596676 346226
rect 596744 346170 596800 346226
rect 596868 346170 596924 346226
rect 596496 346046 596552 346102
rect 596620 346046 596676 346102
rect 596744 346046 596800 346102
rect 596868 346046 596924 346102
rect 596496 345922 596552 345978
rect 596620 345922 596676 345978
rect 596744 345922 596800 345978
rect 596868 345922 596924 345978
rect 596496 328294 596552 328350
rect 596620 328294 596676 328350
rect 596744 328294 596800 328350
rect 596868 328294 596924 328350
rect 596496 328170 596552 328226
rect 596620 328170 596676 328226
rect 596744 328170 596800 328226
rect 596868 328170 596924 328226
rect 596496 328046 596552 328102
rect 596620 328046 596676 328102
rect 596744 328046 596800 328102
rect 596868 328046 596924 328102
rect 596496 327922 596552 327978
rect 596620 327922 596676 327978
rect 596744 327922 596800 327978
rect 596868 327922 596924 327978
rect 596496 310294 596552 310350
rect 596620 310294 596676 310350
rect 596744 310294 596800 310350
rect 596868 310294 596924 310350
rect 596496 310170 596552 310226
rect 596620 310170 596676 310226
rect 596744 310170 596800 310226
rect 596868 310170 596924 310226
rect 596496 310046 596552 310102
rect 596620 310046 596676 310102
rect 596744 310046 596800 310102
rect 596868 310046 596924 310102
rect 596496 309922 596552 309978
rect 596620 309922 596676 309978
rect 596744 309922 596800 309978
rect 596868 309922 596924 309978
rect 596496 292294 596552 292350
rect 596620 292294 596676 292350
rect 596744 292294 596800 292350
rect 596868 292294 596924 292350
rect 596496 292170 596552 292226
rect 596620 292170 596676 292226
rect 596744 292170 596800 292226
rect 596868 292170 596924 292226
rect 596496 292046 596552 292102
rect 596620 292046 596676 292102
rect 596744 292046 596800 292102
rect 596868 292046 596924 292102
rect 596496 291922 596552 291978
rect 596620 291922 596676 291978
rect 596744 291922 596800 291978
rect 596868 291922 596924 291978
rect 596496 274294 596552 274350
rect 596620 274294 596676 274350
rect 596744 274294 596800 274350
rect 596868 274294 596924 274350
rect 596496 274170 596552 274226
rect 596620 274170 596676 274226
rect 596744 274170 596800 274226
rect 596868 274170 596924 274226
rect 596496 274046 596552 274102
rect 596620 274046 596676 274102
rect 596744 274046 596800 274102
rect 596868 274046 596924 274102
rect 596496 273922 596552 273978
rect 596620 273922 596676 273978
rect 596744 273922 596800 273978
rect 596868 273922 596924 273978
rect 588022 46356 588078 46412
rect 588146 46356 588202 46412
rect 588270 46356 588326 46412
rect 588394 46356 588450 46412
rect 588518 46356 588574 46412
rect 588642 46356 588698 46412
rect 588766 46356 588822 46412
rect 588890 46356 588946 46412
rect 589014 46356 589070 46412
rect 589138 46356 589194 46412
rect 588022 46232 588078 46288
rect 588146 46232 588202 46288
rect 588270 46232 588326 46288
rect 588394 46232 588450 46288
rect 588518 46232 588574 46288
rect 588642 46232 588698 46288
rect 588766 46232 588822 46288
rect 588890 46232 588946 46288
rect 589014 46232 589070 46288
rect 589138 46232 589194 46288
rect 588022 46108 588078 46164
rect 588146 46108 588202 46164
rect 588270 46108 588326 46164
rect 588394 46108 588450 46164
rect 588518 46108 588574 46164
rect 588642 46108 588698 46164
rect 588766 46108 588822 46164
rect 588890 46108 588946 46164
rect 589014 46108 589070 46164
rect 589138 46108 589194 46164
rect 588022 45984 588078 46040
rect 588146 45984 588202 46040
rect 588270 45984 588326 46040
rect 588394 45984 588450 46040
rect 588518 45984 588574 46040
rect 588642 45984 588698 46040
rect 588766 45984 588822 46040
rect 588890 45984 588946 46040
rect 589014 45984 589070 46040
rect 589138 45984 589194 46040
rect 588022 45860 588078 45916
rect 588146 45860 588202 45916
rect 588270 45860 588326 45916
rect 588394 45860 588450 45916
rect 588518 45860 588574 45916
rect 588642 45860 588698 45916
rect 588766 45860 588822 45916
rect 588890 45860 588946 45916
rect 589014 45860 589070 45916
rect 589138 45860 589194 45916
rect 586460 42722 586516 42778
rect 596496 256294 596552 256350
rect 596620 256294 596676 256350
rect 596744 256294 596800 256350
rect 596868 256294 596924 256350
rect 596496 256170 596552 256226
rect 596620 256170 596676 256226
rect 596744 256170 596800 256226
rect 596868 256170 596924 256226
rect 596496 256046 596552 256102
rect 596620 256046 596676 256102
rect 596744 256046 596800 256102
rect 596868 256046 596924 256102
rect 596496 255922 596552 255978
rect 596620 255922 596676 255978
rect 596744 255922 596800 255978
rect 596868 255922 596924 255978
rect 596496 238294 596552 238350
rect 596620 238294 596676 238350
rect 596744 238294 596800 238350
rect 596868 238294 596924 238350
rect 596496 238170 596552 238226
rect 596620 238170 596676 238226
rect 596744 238170 596800 238226
rect 596868 238170 596924 238226
rect 596496 238046 596552 238102
rect 596620 238046 596676 238102
rect 596744 238046 596800 238102
rect 596868 238046 596924 238102
rect 596496 237922 596552 237978
rect 596620 237922 596676 237978
rect 596744 237922 596800 237978
rect 596868 237922 596924 237978
rect 596496 220294 596552 220350
rect 596620 220294 596676 220350
rect 596744 220294 596800 220350
rect 596868 220294 596924 220350
rect 596496 220170 596552 220226
rect 596620 220170 596676 220226
rect 596744 220170 596800 220226
rect 596868 220170 596924 220226
rect 596496 220046 596552 220102
rect 596620 220046 596676 220102
rect 596744 220046 596800 220102
rect 596868 220046 596924 220102
rect 596496 219922 596552 219978
rect 596620 219922 596676 219978
rect 596744 219922 596800 219978
rect 596868 219922 596924 219978
rect 596496 202294 596552 202350
rect 596620 202294 596676 202350
rect 596744 202294 596800 202350
rect 596868 202294 596924 202350
rect 596496 202170 596552 202226
rect 596620 202170 596676 202226
rect 596744 202170 596800 202226
rect 596868 202170 596924 202226
rect 596496 202046 596552 202102
rect 596620 202046 596676 202102
rect 596744 202046 596800 202102
rect 596868 202046 596924 202102
rect 596496 201922 596552 201978
rect 596620 201922 596676 201978
rect 596744 201922 596800 201978
rect 596868 201922 596924 201978
rect 596496 184294 596552 184350
rect 596620 184294 596676 184350
rect 596744 184294 596800 184350
rect 596868 184294 596924 184350
rect 596496 184170 596552 184226
rect 596620 184170 596676 184226
rect 596744 184170 596800 184226
rect 596868 184170 596924 184226
rect 596496 184046 596552 184102
rect 596620 184046 596676 184102
rect 596744 184046 596800 184102
rect 596868 184046 596924 184102
rect 596496 183922 596552 183978
rect 596620 183922 596676 183978
rect 596744 183922 596800 183978
rect 596868 183922 596924 183978
rect 596496 166294 596552 166350
rect 596620 166294 596676 166350
rect 596744 166294 596800 166350
rect 596868 166294 596924 166350
rect 596496 166170 596552 166226
rect 596620 166170 596676 166226
rect 596744 166170 596800 166226
rect 596868 166170 596924 166226
rect 596496 166046 596552 166102
rect 596620 166046 596676 166102
rect 596744 166046 596800 166102
rect 596868 166046 596924 166102
rect 596496 165922 596552 165978
rect 596620 165922 596676 165978
rect 596744 165922 596800 165978
rect 596868 165922 596924 165978
rect 596496 148294 596552 148350
rect 596620 148294 596676 148350
rect 596744 148294 596800 148350
rect 596868 148294 596924 148350
rect 596496 148170 596552 148226
rect 596620 148170 596676 148226
rect 596744 148170 596800 148226
rect 596868 148170 596924 148226
rect 596496 148046 596552 148102
rect 596620 148046 596676 148102
rect 596744 148046 596800 148102
rect 596868 148046 596924 148102
rect 596496 147922 596552 147978
rect 596620 147922 596676 147978
rect 596744 147922 596800 147978
rect 596868 147922 596924 147978
rect 596496 130294 596552 130350
rect 596620 130294 596676 130350
rect 596744 130294 596800 130350
rect 596868 130294 596924 130350
rect 596496 130170 596552 130226
rect 596620 130170 596676 130226
rect 596744 130170 596800 130226
rect 596868 130170 596924 130226
rect 596496 130046 596552 130102
rect 596620 130046 596676 130102
rect 596744 130046 596800 130102
rect 596868 130046 596924 130102
rect 596496 129922 596552 129978
rect 596620 129922 596676 129978
rect 596744 129922 596800 129978
rect 596868 129922 596924 129978
rect 596496 112294 596552 112350
rect 596620 112294 596676 112350
rect 596744 112294 596800 112350
rect 596868 112294 596924 112350
rect 596496 112170 596552 112226
rect 596620 112170 596676 112226
rect 596744 112170 596800 112226
rect 596868 112170 596924 112226
rect 596496 112046 596552 112102
rect 596620 112046 596676 112102
rect 596744 112046 596800 112102
rect 596868 112046 596924 112102
rect 596496 111922 596552 111978
rect 596620 111922 596676 111978
rect 596744 111922 596800 111978
rect 596868 111922 596924 111978
rect 596496 94294 596552 94350
rect 596620 94294 596676 94350
rect 596744 94294 596800 94350
rect 596868 94294 596924 94350
rect 596496 94170 596552 94226
rect 596620 94170 596676 94226
rect 596744 94170 596800 94226
rect 596868 94170 596924 94226
rect 596496 94046 596552 94102
rect 596620 94046 596676 94102
rect 596744 94046 596800 94102
rect 596868 94046 596924 94102
rect 596496 93922 596552 93978
rect 596620 93922 596676 93978
rect 596744 93922 596800 93978
rect 596868 93922 596924 93978
rect 596496 76294 596552 76350
rect 596620 76294 596676 76350
rect 596744 76294 596800 76350
rect 596868 76294 596924 76350
rect 596496 76170 596552 76226
rect 596620 76170 596676 76226
rect 596744 76170 596800 76226
rect 596868 76170 596924 76226
rect 596496 76046 596552 76102
rect 596620 76046 596676 76102
rect 596744 76046 596800 76102
rect 596868 76046 596924 76102
rect 596496 75922 596552 75978
rect 596620 75922 596676 75978
rect 596744 75922 596800 75978
rect 596868 75922 596924 75978
rect 591276 30122 591332 30178
rect 588022 28356 588078 28412
rect 588146 28356 588202 28412
rect 588270 28356 588326 28412
rect 588394 28356 588450 28412
rect 588518 28356 588574 28412
rect 588642 28356 588698 28412
rect 588766 28356 588822 28412
rect 588890 28356 588946 28412
rect 589014 28356 589070 28412
rect 589138 28356 589194 28412
rect 588022 28232 588078 28288
rect 588146 28232 588202 28288
rect 588270 28232 588326 28288
rect 588394 28232 588450 28288
rect 588518 28232 588574 28288
rect 588642 28232 588698 28288
rect 588766 28232 588822 28288
rect 588890 28232 588946 28288
rect 589014 28232 589070 28288
rect 589138 28232 589194 28288
rect 588022 28108 588078 28164
rect 588146 28108 588202 28164
rect 588270 28108 588326 28164
rect 588394 28108 588450 28164
rect 588518 28108 588574 28164
rect 588642 28108 588698 28164
rect 588766 28108 588822 28164
rect 588890 28108 588946 28164
rect 589014 28108 589070 28164
rect 589138 28108 589194 28164
rect 588022 27984 588078 28040
rect 588146 27984 588202 28040
rect 588270 27984 588326 28040
rect 588394 27984 588450 28040
rect 588518 27984 588574 28040
rect 588642 27984 588698 28040
rect 588766 27984 588822 28040
rect 588890 27984 588946 28040
rect 589014 27984 589070 28040
rect 589138 27984 589194 28040
rect 588022 27860 588078 27916
rect 588146 27860 588202 27916
rect 588270 27860 588326 27916
rect 588394 27860 588450 27916
rect 588518 27860 588574 27916
rect 588642 27860 588698 27916
rect 588766 27860 588822 27916
rect 588890 27860 588946 27916
rect 589014 27860 589070 27916
rect 589138 27860 589194 27916
rect 593292 30122 593348 30178
rect 591388 25082 591444 25138
rect 596496 58294 596552 58350
rect 596620 58294 596676 58350
rect 596744 58294 596800 58350
rect 596868 58294 596924 58350
rect 596496 58170 596552 58226
rect 596620 58170 596676 58226
rect 596744 58170 596800 58226
rect 596868 58170 596924 58226
rect 596496 58046 596552 58102
rect 596620 58046 596676 58102
rect 596744 58046 596800 58102
rect 596868 58046 596924 58102
rect 596496 57922 596552 57978
rect 596620 57922 596676 57978
rect 596744 57922 596800 57978
rect 596868 57922 596924 57978
rect 596496 40294 596552 40350
rect 596620 40294 596676 40350
rect 596744 40294 596800 40350
rect 596868 40294 596924 40350
rect 596496 40170 596552 40226
rect 596620 40170 596676 40226
rect 596744 40170 596800 40226
rect 596868 40170 596924 40226
rect 596496 40046 596552 40102
rect 596620 40046 596676 40102
rect 596744 40046 596800 40102
rect 596868 40046 596924 40102
rect 596496 39922 596552 39978
rect 596620 39922 596676 39978
rect 596744 39922 596800 39978
rect 596868 39922 596924 39978
rect 596496 22294 596552 22350
rect 596620 22294 596676 22350
rect 596744 22294 596800 22350
rect 596868 22294 596924 22350
rect 596496 22170 596552 22226
rect 596620 22170 596676 22226
rect 596744 22170 596800 22226
rect 596868 22170 596924 22226
rect 596496 22046 596552 22102
rect 596620 22046 596676 22102
rect 596744 22046 596800 22102
rect 596868 22046 596924 22102
rect 596496 21922 596552 21978
rect 596620 21922 596676 21978
rect 596744 21922 596800 21978
rect 596868 21922 596924 21978
rect 596496 4294 596552 4350
rect 596620 4294 596676 4350
rect 596744 4294 596800 4350
rect 596868 4294 596924 4350
rect 596496 4170 596552 4226
rect 596620 4170 596676 4226
rect 596744 4170 596800 4226
rect 596868 4170 596924 4226
rect 596496 4046 596552 4102
rect 596620 4046 596676 4102
rect 596744 4046 596800 4102
rect 596868 4046 596924 4102
rect 596496 3922 596552 3978
rect 596620 3922 596676 3978
rect 596744 3922 596800 3978
rect 596868 3922 596924 3978
rect 596496 -216 596552 -160
rect 596620 -216 596676 -160
rect 596744 -216 596800 -160
rect 596868 -216 596924 -160
rect 596496 -340 596552 -284
rect 596620 -340 596676 -284
rect 596744 -340 596800 -284
rect 596868 -340 596924 -284
rect 596496 -464 596552 -408
rect 596620 -464 596676 -408
rect 596744 -464 596800 -408
rect 596868 -464 596924 -408
rect 596496 -588 596552 -532
rect 596620 -588 596676 -532
rect 596744 -588 596800 -532
rect 596868 -588 596924 -532
rect 597456 586294 597512 586350
rect 597580 586294 597636 586350
rect 597704 586294 597760 586350
rect 597828 586294 597884 586350
rect 597456 586170 597512 586226
rect 597580 586170 597636 586226
rect 597704 586170 597760 586226
rect 597828 586170 597884 586226
rect 597456 586046 597512 586102
rect 597580 586046 597636 586102
rect 597704 586046 597760 586102
rect 597828 586046 597884 586102
rect 597456 585922 597512 585978
rect 597580 585922 597636 585978
rect 597704 585922 597760 585978
rect 597828 585922 597884 585978
rect 597456 568294 597512 568350
rect 597580 568294 597636 568350
rect 597704 568294 597760 568350
rect 597828 568294 597884 568350
rect 597456 568170 597512 568226
rect 597580 568170 597636 568226
rect 597704 568170 597760 568226
rect 597828 568170 597884 568226
rect 597456 568046 597512 568102
rect 597580 568046 597636 568102
rect 597704 568046 597760 568102
rect 597828 568046 597884 568102
rect 597456 567922 597512 567978
rect 597580 567922 597636 567978
rect 597704 567922 597760 567978
rect 597828 567922 597884 567978
rect 597456 550294 597512 550350
rect 597580 550294 597636 550350
rect 597704 550294 597760 550350
rect 597828 550294 597884 550350
rect 597456 550170 597512 550226
rect 597580 550170 597636 550226
rect 597704 550170 597760 550226
rect 597828 550170 597884 550226
rect 597456 550046 597512 550102
rect 597580 550046 597636 550102
rect 597704 550046 597760 550102
rect 597828 550046 597884 550102
rect 597456 549922 597512 549978
rect 597580 549922 597636 549978
rect 597704 549922 597760 549978
rect 597828 549922 597884 549978
rect 597456 532294 597512 532350
rect 597580 532294 597636 532350
rect 597704 532294 597760 532350
rect 597828 532294 597884 532350
rect 597456 532170 597512 532226
rect 597580 532170 597636 532226
rect 597704 532170 597760 532226
rect 597828 532170 597884 532226
rect 597456 532046 597512 532102
rect 597580 532046 597636 532102
rect 597704 532046 597760 532102
rect 597828 532046 597884 532102
rect 597456 531922 597512 531978
rect 597580 531922 597636 531978
rect 597704 531922 597760 531978
rect 597828 531922 597884 531978
rect 597456 514294 597512 514350
rect 597580 514294 597636 514350
rect 597704 514294 597760 514350
rect 597828 514294 597884 514350
rect 597456 514170 597512 514226
rect 597580 514170 597636 514226
rect 597704 514170 597760 514226
rect 597828 514170 597884 514226
rect 597456 514046 597512 514102
rect 597580 514046 597636 514102
rect 597704 514046 597760 514102
rect 597828 514046 597884 514102
rect 597456 513922 597512 513978
rect 597580 513922 597636 513978
rect 597704 513922 597760 513978
rect 597828 513922 597884 513978
rect 597456 496294 597512 496350
rect 597580 496294 597636 496350
rect 597704 496294 597760 496350
rect 597828 496294 597884 496350
rect 597456 496170 597512 496226
rect 597580 496170 597636 496226
rect 597704 496170 597760 496226
rect 597828 496170 597884 496226
rect 597456 496046 597512 496102
rect 597580 496046 597636 496102
rect 597704 496046 597760 496102
rect 597828 496046 597884 496102
rect 597456 495922 597512 495978
rect 597580 495922 597636 495978
rect 597704 495922 597760 495978
rect 597828 495922 597884 495978
rect 597456 478294 597512 478350
rect 597580 478294 597636 478350
rect 597704 478294 597760 478350
rect 597828 478294 597884 478350
rect 597456 478170 597512 478226
rect 597580 478170 597636 478226
rect 597704 478170 597760 478226
rect 597828 478170 597884 478226
rect 597456 478046 597512 478102
rect 597580 478046 597636 478102
rect 597704 478046 597760 478102
rect 597828 478046 597884 478102
rect 597456 477922 597512 477978
rect 597580 477922 597636 477978
rect 597704 477922 597760 477978
rect 597828 477922 597884 477978
rect 597456 460294 597512 460350
rect 597580 460294 597636 460350
rect 597704 460294 597760 460350
rect 597828 460294 597884 460350
rect 597456 460170 597512 460226
rect 597580 460170 597636 460226
rect 597704 460170 597760 460226
rect 597828 460170 597884 460226
rect 597456 460046 597512 460102
rect 597580 460046 597636 460102
rect 597704 460046 597760 460102
rect 597828 460046 597884 460102
rect 597456 459922 597512 459978
rect 597580 459922 597636 459978
rect 597704 459922 597760 459978
rect 597828 459922 597884 459978
rect 597456 442294 597512 442350
rect 597580 442294 597636 442350
rect 597704 442294 597760 442350
rect 597828 442294 597884 442350
rect 597456 442170 597512 442226
rect 597580 442170 597636 442226
rect 597704 442170 597760 442226
rect 597828 442170 597884 442226
rect 597456 442046 597512 442102
rect 597580 442046 597636 442102
rect 597704 442046 597760 442102
rect 597828 442046 597884 442102
rect 597456 441922 597512 441978
rect 597580 441922 597636 441978
rect 597704 441922 597760 441978
rect 597828 441922 597884 441978
rect 597456 424294 597512 424350
rect 597580 424294 597636 424350
rect 597704 424294 597760 424350
rect 597828 424294 597884 424350
rect 597456 424170 597512 424226
rect 597580 424170 597636 424226
rect 597704 424170 597760 424226
rect 597828 424170 597884 424226
rect 597456 424046 597512 424102
rect 597580 424046 597636 424102
rect 597704 424046 597760 424102
rect 597828 424046 597884 424102
rect 597456 423922 597512 423978
rect 597580 423922 597636 423978
rect 597704 423922 597760 423978
rect 597828 423922 597884 423978
rect 597456 406294 597512 406350
rect 597580 406294 597636 406350
rect 597704 406294 597760 406350
rect 597828 406294 597884 406350
rect 597456 406170 597512 406226
rect 597580 406170 597636 406226
rect 597704 406170 597760 406226
rect 597828 406170 597884 406226
rect 597456 406046 597512 406102
rect 597580 406046 597636 406102
rect 597704 406046 597760 406102
rect 597828 406046 597884 406102
rect 597456 405922 597512 405978
rect 597580 405922 597636 405978
rect 597704 405922 597760 405978
rect 597828 405922 597884 405978
rect 597456 388294 597512 388350
rect 597580 388294 597636 388350
rect 597704 388294 597760 388350
rect 597828 388294 597884 388350
rect 597456 388170 597512 388226
rect 597580 388170 597636 388226
rect 597704 388170 597760 388226
rect 597828 388170 597884 388226
rect 597456 388046 597512 388102
rect 597580 388046 597636 388102
rect 597704 388046 597760 388102
rect 597828 388046 597884 388102
rect 597456 387922 597512 387978
rect 597580 387922 597636 387978
rect 597704 387922 597760 387978
rect 597828 387922 597884 387978
rect 597456 370294 597512 370350
rect 597580 370294 597636 370350
rect 597704 370294 597760 370350
rect 597828 370294 597884 370350
rect 597456 370170 597512 370226
rect 597580 370170 597636 370226
rect 597704 370170 597760 370226
rect 597828 370170 597884 370226
rect 597456 370046 597512 370102
rect 597580 370046 597636 370102
rect 597704 370046 597760 370102
rect 597828 370046 597884 370102
rect 597456 369922 597512 369978
rect 597580 369922 597636 369978
rect 597704 369922 597760 369978
rect 597828 369922 597884 369978
rect 597456 352294 597512 352350
rect 597580 352294 597636 352350
rect 597704 352294 597760 352350
rect 597828 352294 597884 352350
rect 597456 352170 597512 352226
rect 597580 352170 597636 352226
rect 597704 352170 597760 352226
rect 597828 352170 597884 352226
rect 597456 352046 597512 352102
rect 597580 352046 597636 352102
rect 597704 352046 597760 352102
rect 597828 352046 597884 352102
rect 597456 351922 597512 351978
rect 597580 351922 597636 351978
rect 597704 351922 597760 351978
rect 597828 351922 597884 351978
rect 597456 334294 597512 334350
rect 597580 334294 597636 334350
rect 597704 334294 597760 334350
rect 597828 334294 597884 334350
rect 597456 334170 597512 334226
rect 597580 334170 597636 334226
rect 597704 334170 597760 334226
rect 597828 334170 597884 334226
rect 597456 334046 597512 334102
rect 597580 334046 597636 334102
rect 597704 334046 597760 334102
rect 597828 334046 597884 334102
rect 597456 333922 597512 333978
rect 597580 333922 597636 333978
rect 597704 333922 597760 333978
rect 597828 333922 597884 333978
rect 597456 316294 597512 316350
rect 597580 316294 597636 316350
rect 597704 316294 597760 316350
rect 597828 316294 597884 316350
rect 597456 316170 597512 316226
rect 597580 316170 597636 316226
rect 597704 316170 597760 316226
rect 597828 316170 597884 316226
rect 597456 316046 597512 316102
rect 597580 316046 597636 316102
rect 597704 316046 597760 316102
rect 597828 316046 597884 316102
rect 597456 315922 597512 315978
rect 597580 315922 597636 315978
rect 597704 315922 597760 315978
rect 597828 315922 597884 315978
rect 597456 298294 597512 298350
rect 597580 298294 597636 298350
rect 597704 298294 597760 298350
rect 597828 298294 597884 298350
rect 597456 298170 597512 298226
rect 597580 298170 597636 298226
rect 597704 298170 597760 298226
rect 597828 298170 597884 298226
rect 597456 298046 597512 298102
rect 597580 298046 597636 298102
rect 597704 298046 597760 298102
rect 597828 298046 597884 298102
rect 597456 297922 597512 297978
rect 597580 297922 597636 297978
rect 597704 297922 597760 297978
rect 597828 297922 597884 297978
rect 597456 280294 597512 280350
rect 597580 280294 597636 280350
rect 597704 280294 597760 280350
rect 597828 280294 597884 280350
rect 597456 280170 597512 280226
rect 597580 280170 597636 280226
rect 597704 280170 597760 280226
rect 597828 280170 597884 280226
rect 597456 280046 597512 280102
rect 597580 280046 597636 280102
rect 597704 280046 597760 280102
rect 597828 280046 597884 280102
rect 597456 279922 597512 279978
rect 597580 279922 597636 279978
rect 597704 279922 597760 279978
rect 597828 279922 597884 279978
rect 597456 262294 597512 262350
rect 597580 262294 597636 262350
rect 597704 262294 597760 262350
rect 597828 262294 597884 262350
rect 597456 262170 597512 262226
rect 597580 262170 597636 262226
rect 597704 262170 597760 262226
rect 597828 262170 597884 262226
rect 597456 262046 597512 262102
rect 597580 262046 597636 262102
rect 597704 262046 597760 262102
rect 597828 262046 597884 262102
rect 597456 261922 597512 261978
rect 597580 261922 597636 261978
rect 597704 261922 597760 261978
rect 597828 261922 597884 261978
rect 597456 244294 597512 244350
rect 597580 244294 597636 244350
rect 597704 244294 597760 244350
rect 597828 244294 597884 244350
rect 597456 244170 597512 244226
rect 597580 244170 597636 244226
rect 597704 244170 597760 244226
rect 597828 244170 597884 244226
rect 597456 244046 597512 244102
rect 597580 244046 597636 244102
rect 597704 244046 597760 244102
rect 597828 244046 597884 244102
rect 597456 243922 597512 243978
rect 597580 243922 597636 243978
rect 597704 243922 597760 243978
rect 597828 243922 597884 243978
rect 597456 226294 597512 226350
rect 597580 226294 597636 226350
rect 597704 226294 597760 226350
rect 597828 226294 597884 226350
rect 597456 226170 597512 226226
rect 597580 226170 597636 226226
rect 597704 226170 597760 226226
rect 597828 226170 597884 226226
rect 597456 226046 597512 226102
rect 597580 226046 597636 226102
rect 597704 226046 597760 226102
rect 597828 226046 597884 226102
rect 597456 225922 597512 225978
rect 597580 225922 597636 225978
rect 597704 225922 597760 225978
rect 597828 225922 597884 225978
rect 597456 208294 597512 208350
rect 597580 208294 597636 208350
rect 597704 208294 597760 208350
rect 597828 208294 597884 208350
rect 597456 208170 597512 208226
rect 597580 208170 597636 208226
rect 597704 208170 597760 208226
rect 597828 208170 597884 208226
rect 597456 208046 597512 208102
rect 597580 208046 597636 208102
rect 597704 208046 597760 208102
rect 597828 208046 597884 208102
rect 597456 207922 597512 207978
rect 597580 207922 597636 207978
rect 597704 207922 597760 207978
rect 597828 207922 597884 207978
rect 597456 190294 597512 190350
rect 597580 190294 597636 190350
rect 597704 190294 597760 190350
rect 597828 190294 597884 190350
rect 597456 190170 597512 190226
rect 597580 190170 597636 190226
rect 597704 190170 597760 190226
rect 597828 190170 597884 190226
rect 597456 190046 597512 190102
rect 597580 190046 597636 190102
rect 597704 190046 597760 190102
rect 597828 190046 597884 190102
rect 597456 189922 597512 189978
rect 597580 189922 597636 189978
rect 597704 189922 597760 189978
rect 597828 189922 597884 189978
rect 597456 172294 597512 172350
rect 597580 172294 597636 172350
rect 597704 172294 597760 172350
rect 597828 172294 597884 172350
rect 597456 172170 597512 172226
rect 597580 172170 597636 172226
rect 597704 172170 597760 172226
rect 597828 172170 597884 172226
rect 597456 172046 597512 172102
rect 597580 172046 597636 172102
rect 597704 172046 597760 172102
rect 597828 172046 597884 172102
rect 597456 171922 597512 171978
rect 597580 171922 597636 171978
rect 597704 171922 597760 171978
rect 597828 171922 597884 171978
rect 597456 154294 597512 154350
rect 597580 154294 597636 154350
rect 597704 154294 597760 154350
rect 597828 154294 597884 154350
rect 597456 154170 597512 154226
rect 597580 154170 597636 154226
rect 597704 154170 597760 154226
rect 597828 154170 597884 154226
rect 597456 154046 597512 154102
rect 597580 154046 597636 154102
rect 597704 154046 597760 154102
rect 597828 154046 597884 154102
rect 597456 153922 597512 153978
rect 597580 153922 597636 153978
rect 597704 153922 597760 153978
rect 597828 153922 597884 153978
rect 597456 136294 597512 136350
rect 597580 136294 597636 136350
rect 597704 136294 597760 136350
rect 597828 136294 597884 136350
rect 597456 136170 597512 136226
rect 597580 136170 597636 136226
rect 597704 136170 597760 136226
rect 597828 136170 597884 136226
rect 597456 136046 597512 136102
rect 597580 136046 597636 136102
rect 597704 136046 597760 136102
rect 597828 136046 597884 136102
rect 597456 135922 597512 135978
rect 597580 135922 597636 135978
rect 597704 135922 597760 135978
rect 597828 135922 597884 135978
rect 597456 118294 597512 118350
rect 597580 118294 597636 118350
rect 597704 118294 597760 118350
rect 597828 118294 597884 118350
rect 597456 118170 597512 118226
rect 597580 118170 597636 118226
rect 597704 118170 597760 118226
rect 597828 118170 597884 118226
rect 597456 118046 597512 118102
rect 597580 118046 597636 118102
rect 597704 118046 597760 118102
rect 597828 118046 597884 118102
rect 597456 117922 597512 117978
rect 597580 117922 597636 117978
rect 597704 117922 597760 117978
rect 597828 117922 597884 117978
rect 597456 100294 597512 100350
rect 597580 100294 597636 100350
rect 597704 100294 597760 100350
rect 597828 100294 597884 100350
rect 597456 100170 597512 100226
rect 597580 100170 597636 100226
rect 597704 100170 597760 100226
rect 597828 100170 597884 100226
rect 597456 100046 597512 100102
rect 597580 100046 597636 100102
rect 597704 100046 597760 100102
rect 597828 100046 597884 100102
rect 597456 99922 597512 99978
rect 597580 99922 597636 99978
rect 597704 99922 597760 99978
rect 597828 99922 597884 99978
rect 597456 82294 597512 82350
rect 597580 82294 597636 82350
rect 597704 82294 597760 82350
rect 597828 82294 597884 82350
rect 597456 82170 597512 82226
rect 597580 82170 597636 82226
rect 597704 82170 597760 82226
rect 597828 82170 597884 82226
rect 597456 82046 597512 82102
rect 597580 82046 597636 82102
rect 597704 82046 597760 82102
rect 597828 82046 597884 82102
rect 597456 81922 597512 81978
rect 597580 81922 597636 81978
rect 597704 81922 597760 81978
rect 597828 81922 597884 81978
rect 597456 64294 597512 64350
rect 597580 64294 597636 64350
rect 597704 64294 597760 64350
rect 597828 64294 597884 64350
rect 597456 64170 597512 64226
rect 597580 64170 597636 64226
rect 597704 64170 597760 64226
rect 597828 64170 597884 64226
rect 597456 64046 597512 64102
rect 597580 64046 597636 64102
rect 597704 64046 597760 64102
rect 597828 64046 597884 64102
rect 597456 63922 597512 63978
rect 597580 63922 597636 63978
rect 597704 63922 597760 63978
rect 597828 63922 597884 63978
rect 597456 46294 597512 46350
rect 597580 46294 597636 46350
rect 597704 46294 597760 46350
rect 597828 46294 597884 46350
rect 597456 46170 597512 46226
rect 597580 46170 597636 46226
rect 597704 46170 597760 46226
rect 597828 46170 597884 46226
rect 597456 46046 597512 46102
rect 597580 46046 597636 46102
rect 597704 46046 597760 46102
rect 597828 46046 597884 46102
rect 597456 45922 597512 45978
rect 597580 45922 597636 45978
rect 597704 45922 597760 45978
rect 597828 45922 597884 45978
rect 597456 28294 597512 28350
rect 597580 28294 597636 28350
rect 597704 28294 597760 28350
rect 597828 28294 597884 28350
rect 597456 28170 597512 28226
rect 597580 28170 597636 28226
rect 597704 28170 597760 28226
rect 597828 28170 597884 28226
rect 597456 28046 597512 28102
rect 597580 28046 597636 28102
rect 597704 28046 597760 28102
rect 597828 28046 597884 28102
rect 597456 27922 597512 27978
rect 597580 27922 597636 27978
rect 597704 27922 597760 27978
rect 597828 27922 597884 27978
rect 597456 10294 597512 10350
rect 597580 10294 597636 10350
rect 597704 10294 597760 10350
rect 597828 10294 597884 10350
rect 597456 10170 597512 10226
rect 597580 10170 597636 10226
rect 597704 10170 597760 10226
rect 597828 10170 597884 10226
rect 597456 10046 597512 10102
rect 597580 10046 597636 10102
rect 597704 10046 597760 10102
rect 597828 10046 597884 10102
rect 597456 9922 597512 9978
rect 597580 9922 597636 9978
rect 597704 9922 597760 9978
rect 597828 9922 597884 9978
rect 582970 -1176 583026 -1120
rect 583094 -1176 583150 -1120
rect 583218 -1176 583274 -1120
rect 583342 -1176 583398 -1120
rect 582970 -1300 583026 -1244
rect 583094 -1300 583150 -1244
rect 583218 -1300 583274 -1244
rect 583342 -1300 583398 -1244
rect 582970 -1424 583026 -1368
rect 583094 -1424 583150 -1368
rect 583218 -1424 583274 -1368
rect 583342 -1424 583398 -1368
rect 582970 -1548 583026 -1492
rect 583094 -1548 583150 -1492
rect 583218 -1548 583274 -1492
rect 583342 -1548 583398 -1492
rect 597456 -1176 597512 -1120
rect 597580 -1176 597636 -1120
rect 597704 -1176 597760 -1120
rect 597828 -1176 597884 -1120
rect 597456 -1300 597512 -1244
rect 597580 -1300 597636 -1244
rect 597704 -1300 597760 -1244
rect 597828 -1300 597884 -1244
rect 597456 -1424 597512 -1368
rect 597580 -1424 597636 -1368
rect 597704 -1424 597760 -1368
rect 597828 -1424 597884 -1368
rect 597456 -1548 597512 -1492
rect 597580 -1548 597636 -1492
rect 597704 -1548 597760 -1492
rect 597828 -1548 597884 -1492
<< metal5 >>
rect -1916 598172 597980 598268
rect -1916 598116 -1820 598172
rect -1764 598116 -1696 598172
rect -1640 598116 -1572 598172
rect -1516 598116 -1448 598172
rect -1392 598116 6970 598172
rect 7026 598116 7094 598172
rect 7150 598116 7218 598172
rect 7274 598116 7342 598172
rect 7398 598116 24970 598172
rect 25026 598116 25094 598172
rect 25150 598116 25218 598172
rect 25274 598116 25342 598172
rect 25398 598116 42970 598172
rect 43026 598116 43094 598172
rect 43150 598116 43218 598172
rect 43274 598116 43342 598172
rect 43398 598116 60970 598172
rect 61026 598116 61094 598172
rect 61150 598116 61218 598172
rect 61274 598116 61342 598172
rect 61398 598116 78970 598172
rect 79026 598116 79094 598172
rect 79150 598116 79218 598172
rect 79274 598116 79342 598172
rect 79398 598116 96970 598172
rect 97026 598116 97094 598172
rect 97150 598116 97218 598172
rect 97274 598116 97342 598172
rect 97398 598116 132970 598172
rect 133026 598116 133094 598172
rect 133150 598116 133218 598172
rect 133274 598116 133342 598172
rect 133398 598116 150970 598172
rect 151026 598116 151094 598172
rect 151150 598116 151218 598172
rect 151274 598116 151342 598172
rect 151398 598116 168970 598172
rect 169026 598116 169094 598172
rect 169150 598116 169218 598172
rect 169274 598116 169342 598172
rect 169398 598116 186970 598172
rect 187026 598116 187094 598172
rect 187150 598116 187218 598172
rect 187274 598116 187342 598172
rect 187398 598116 222970 598172
rect 223026 598116 223094 598172
rect 223150 598116 223218 598172
rect 223274 598116 223342 598172
rect 223398 598116 240970 598172
rect 241026 598116 241094 598172
rect 241150 598116 241218 598172
rect 241274 598116 241342 598172
rect 241398 598116 258970 598172
rect 259026 598116 259094 598172
rect 259150 598116 259218 598172
rect 259274 598116 259342 598172
rect 259398 598116 276970 598172
rect 277026 598116 277094 598172
rect 277150 598116 277218 598172
rect 277274 598116 277342 598172
rect 277398 598116 312970 598172
rect 313026 598116 313094 598172
rect 313150 598116 313218 598172
rect 313274 598116 313342 598172
rect 313398 598116 330970 598172
rect 331026 598116 331094 598172
rect 331150 598116 331218 598172
rect 331274 598116 331342 598172
rect 331398 598116 348970 598172
rect 349026 598116 349094 598172
rect 349150 598116 349218 598172
rect 349274 598116 349342 598172
rect 349398 598116 366970 598172
rect 367026 598116 367094 598172
rect 367150 598116 367218 598172
rect 367274 598116 367342 598172
rect 367398 598116 402970 598172
rect 403026 598116 403094 598172
rect 403150 598116 403218 598172
rect 403274 598116 403342 598172
rect 403398 598116 420970 598172
rect 421026 598116 421094 598172
rect 421150 598116 421218 598172
rect 421274 598116 421342 598172
rect 421398 598116 438970 598172
rect 439026 598116 439094 598172
rect 439150 598116 439218 598172
rect 439274 598116 439342 598172
rect 439398 598116 456970 598172
rect 457026 598116 457094 598172
rect 457150 598116 457218 598172
rect 457274 598116 457342 598172
rect 457398 598116 492970 598172
rect 493026 598116 493094 598172
rect 493150 598116 493218 598172
rect 493274 598116 493342 598172
rect 493398 598116 510970 598172
rect 511026 598116 511094 598172
rect 511150 598116 511218 598172
rect 511274 598116 511342 598172
rect 511398 598116 528970 598172
rect 529026 598116 529094 598172
rect 529150 598116 529218 598172
rect 529274 598116 529342 598172
rect 529398 598116 546970 598172
rect 547026 598116 547094 598172
rect 547150 598116 547218 598172
rect 547274 598116 547342 598172
rect 547398 598116 564970 598172
rect 565026 598116 565094 598172
rect 565150 598116 565218 598172
rect 565274 598116 565342 598172
rect 565398 598116 582970 598172
rect 583026 598116 583094 598172
rect 583150 598116 583218 598172
rect 583274 598116 583342 598172
rect 583398 598116 597456 598172
rect 597512 598116 597580 598172
rect 597636 598116 597704 598172
rect 597760 598116 597828 598172
rect 597884 598116 597980 598172
rect -1916 598048 597980 598116
rect -1916 597992 -1820 598048
rect -1764 597992 -1696 598048
rect -1640 597992 -1572 598048
rect -1516 597992 -1448 598048
rect -1392 597992 6970 598048
rect 7026 597992 7094 598048
rect 7150 597992 7218 598048
rect 7274 597992 7342 598048
rect 7398 597992 24970 598048
rect 25026 597992 25094 598048
rect 25150 597992 25218 598048
rect 25274 597992 25342 598048
rect 25398 597992 42970 598048
rect 43026 597992 43094 598048
rect 43150 597992 43218 598048
rect 43274 597992 43342 598048
rect 43398 597992 60970 598048
rect 61026 597992 61094 598048
rect 61150 597992 61218 598048
rect 61274 597992 61342 598048
rect 61398 597992 78970 598048
rect 79026 597992 79094 598048
rect 79150 597992 79218 598048
rect 79274 597992 79342 598048
rect 79398 597992 96970 598048
rect 97026 597992 97094 598048
rect 97150 597992 97218 598048
rect 97274 597992 97342 598048
rect 97398 597992 132970 598048
rect 133026 597992 133094 598048
rect 133150 597992 133218 598048
rect 133274 597992 133342 598048
rect 133398 597992 150970 598048
rect 151026 597992 151094 598048
rect 151150 597992 151218 598048
rect 151274 597992 151342 598048
rect 151398 597992 168970 598048
rect 169026 597992 169094 598048
rect 169150 597992 169218 598048
rect 169274 597992 169342 598048
rect 169398 597992 186970 598048
rect 187026 597992 187094 598048
rect 187150 597992 187218 598048
rect 187274 597992 187342 598048
rect 187398 597992 222970 598048
rect 223026 597992 223094 598048
rect 223150 597992 223218 598048
rect 223274 597992 223342 598048
rect 223398 597992 240970 598048
rect 241026 597992 241094 598048
rect 241150 597992 241218 598048
rect 241274 597992 241342 598048
rect 241398 597992 258970 598048
rect 259026 597992 259094 598048
rect 259150 597992 259218 598048
rect 259274 597992 259342 598048
rect 259398 597992 276970 598048
rect 277026 597992 277094 598048
rect 277150 597992 277218 598048
rect 277274 597992 277342 598048
rect 277398 597992 312970 598048
rect 313026 597992 313094 598048
rect 313150 597992 313218 598048
rect 313274 597992 313342 598048
rect 313398 597992 330970 598048
rect 331026 597992 331094 598048
rect 331150 597992 331218 598048
rect 331274 597992 331342 598048
rect 331398 597992 348970 598048
rect 349026 597992 349094 598048
rect 349150 597992 349218 598048
rect 349274 597992 349342 598048
rect 349398 597992 366970 598048
rect 367026 597992 367094 598048
rect 367150 597992 367218 598048
rect 367274 597992 367342 598048
rect 367398 597992 402970 598048
rect 403026 597992 403094 598048
rect 403150 597992 403218 598048
rect 403274 597992 403342 598048
rect 403398 597992 420970 598048
rect 421026 597992 421094 598048
rect 421150 597992 421218 598048
rect 421274 597992 421342 598048
rect 421398 597992 438970 598048
rect 439026 597992 439094 598048
rect 439150 597992 439218 598048
rect 439274 597992 439342 598048
rect 439398 597992 456970 598048
rect 457026 597992 457094 598048
rect 457150 597992 457218 598048
rect 457274 597992 457342 598048
rect 457398 597992 492970 598048
rect 493026 597992 493094 598048
rect 493150 597992 493218 598048
rect 493274 597992 493342 598048
rect 493398 597992 510970 598048
rect 511026 597992 511094 598048
rect 511150 597992 511218 598048
rect 511274 597992 511342 598048
rect 511398 597992 528970 598048
rect 529026 597992 529094 598048
rect 529150 597992 529218 598048
rect 529274 597992 529342 598048
rect 529398 597992 546970 598048
rect 547026 597992 547094 598048
rect 547150 597992 547218 598048
rect 547274 597992 547342 598048
rect 547398 597992 564970 598048
rect 565026 597992 565094 598048
rect 565150 597992 565218 598048
rect 565274 597992 565342 598048
rect 565398 597992 582970 598048
rect 583026 597992 583094 598048
rect 583150 597992 583218 598048
rect 583274 597992 583342 598048
rect 583398 597992 597456 598048
rect 597512 597992 597580 598048
rect 597636 597992 597704 598048
rect 597760 597992 597828 598048
rect 597884 597992 597980 598048
rect -1916 597924 597980 597992
rect -1916 597868 -1820 597924
rect -1764 597868 -1696 597924
rect -1640 597868 -1572 597924
rect -1516 597868 -1448 597924
rect -1392 597868 6970 597924
rect 7026 597868 7094 597924
rect 7150 597868 7218 597924
rect 7274 597868 7342 597924
rect 7398 597868 24970 597924
rect 25026 597868 25094 597924
rect 25150 597868 25218 597924
rect 25274 597868 25342 597924
rect 25398 597868 42970 597924
rect 43026 597868 43094 597924
rect 43150 597868 43218 597924
rect 43274 597868 43342 597924
rect 43398 597868 60970 597924
rect 61026 597868 61094 597924
rect 61150 597868 61218 597924
rect 61274 597868 61342 597924
rect 61398 597868 78970 597924
rect 79026 597868 79094 597924
rect 79150 597868 79218 597924
rect 79274 597868 79342 597924
rect 79398 597868 96970 597924
rect 97026 597868 97094 597924
rect 97150 597868 97218 597924
rect 97274 597868 97342 597924
rect 97398 597868 132970 597924
rect 133026 597868 133094 597924
rect 133150 597868 133218 597924
rect 133274 597868 133342 597924
rect 133398 597868 150970 597924
rect 151026 597868 151094 597924
rect 151150 597868 151218 597924
rect 151274 597868 151342 597924
rect 151398 597868 168970 597924
rect 169026 597868 169094 597924
rect 169150 597868 169218 597924
rect 169274 597868 169342 597924
rect 169398 597868 186970 597924
rect 187026 597868 187094 597924
rect 187150 597868 187218 597924
rect 187274 597868 187342 597924
rect 187398 597868 222970 597924
rect 223026 597868 223094 597924
rect 223150 597868 223218 597924
rect 223274 597868 223342 597924
rect 223398 597868 240970 597924
rect 241026 597868 241094 597924
rect 241150 597868 241218 597924
rect 241274 597868 241342 597924
rect 241398 597868 258970 597924
rect 259026 597868 259094 597924
rect 259150 597868 259218 597924
rect 259274 597868 259342 597924
rect 259398 597868 276970 597924
rect 277026 597868 277094 597924
rect 277150 597868 277218 597924
rect 277274 597868 277342 597924
rect 277398 597868 312970 597924
rect 313026 597868 313094 597924
rect 313150 597868 313218 597924
rect 313274 597868 313342 597924
rect 313398 597868 330970 597924
rect 331026 597868 331094 597924
rect 331150 597868 331218 597924
rect 331274 597868 331342 597924
rect 331398 597868 348970 597924
rect 349026 597868 349094 597924
rect 349150 597868 349218 597924
rect 349274 597868 349342 597924
rect 349398 597868 366970 597924
rect 367026 597868 367094 597924
rect 367150 597868 367218 597924
rect 367274 597868 367342 597924
rect 367398 597868 402970 597924
rect 403026 597868 403094 597924
rect 403150 597868 403218 597924
rect 403274 597868 403342 597924
rect 403398 597868 420970 597924
rect 421026 597868 421094 597924
rect 421150 597868 421218 597924
rect 421274 597868 421342 597924
rect 421398 597868 438970 597924
rect 439026 597868 439094 597924
rect 439150 597868 439218 597924
rect 439274 597868 439342 597924
rect 439398 597868 456970 597924
rect 457026 597868 457094 597924
rect 457150 597868 457218 597924
rect 457274 597868 457342 597924
rect 457398 597868 492970 597924
rect 493026 597868 493094 597924
rect 493150 597868 493218 597924
rect 493274 597868 493342 597924
rect 493398 597868 510970 597924
rect 511026 597868 511094 597924
rect 511150 597868 511218 597924
rect 511274 597868 511342 597924
rect 511398 597868 528970 597924
rect 529026 597868 529094 597924
rect 529150 597868 529218 597924
rect 529274 597868 529342 597924
rect 529398 597868 546970 597924
rect 547026 597868 547094 597924
rect 547150 597868 547218 597924
rect 547274 597868 547342 597924
rect 547398 597868 564970 597924
rect 565026 597868 565094 597924
rect 565150 597868 565218 597924
rect 565274 597868 565342 597924
rect 565398 597868 582970 597924
rect 583026 597868 583094 597924
rect 583150 597868 583218 597924
rect 583274 597868 583342 597924
rect 583398 597868 597456 597924
rect 597512 597868 597580 597924
rect 597636 597868 597704 597924
rect 597760 597868 597828 597924
rect 597884 597868 597980 597924
rect -1916 597800 597980 597868
rect -1916 597744 -1820 597800
rect -1764 597744 -1696 597800
rect -1640 597744 -1572 597800
rect -1516 597744 -1448 597800
rect -1392 597744 6970 597800
rect 7026 597744 7094 597800
rect 7150 597744 7218 597800
rect 7274 597744 7342 597800
rect 7398 597744 24970 597800
rect 25026 597744 25094 597800
rect 25150 597744 25218 597800
rect 25274 597744 25342 597800
rect 25398 597744 42970 597800
rect 43026 597744 43094 597800
rect 43150 597744 43218 597800
rect 43274 597744 43342 597800
rect 43398 597744 60970 597800
rect 61026 597744 61094 597800
rect 61150 597744 61218 597800
rect 61274 597744 61342 597800
rect 61398 597744 78970 597800
rect 79026 597744 79094 597800
rect 79150 597744 79218 597800
rect 79274 597744 79342 597800
rect 79398 597744 96970 597800
rect 97026 597744 97094 597800
rect 97150 597744 97218 597800
rect 97274 597744 97342 597800
rect 97398 597744 132970 597800
rect 133026 597744 133094 597800
rect 133150 597744 133218 597800
rect 133274 597744 133342 597800
rect 133398 597744 150970 597800
rect 151026 597744 151094 597800
rect 151150 597744 151218 597800
rect 151274 597744 151342 597800
rect 151398 597744 168970 597800
rect 169026 597744 169094 597800
rect 169150 597744 169218 597800
rect 169274 597744 169342 597800
rect 169398 597744 186970 597800
rect 187026 597744 187094 597800
rect 187150 597744 187218 597800
rect 187274 597744 187342 597800
rect 187398 597744 222970 597800
rect 223026 597744 223094 597800
rect 223150 597744 223218 597800
rect 223274 597744 223342 597800
rect 223398 597744 240970 597800
rect 241026 597744 241094 597800
rect 241150 597744 241218 597800
rect 241274 597744 241342 597800
rect 241398 597744 258970 597800
rect 259026 597744 259094 597800
rect 259150 597744 259218 597800
rect 259274 597744 259342 597800
rect 259398 597744 276970 597800
rect 277026 597744 277094 597800
rect 277150 597744 277218 597800
rect 277274 597744 277342 597800
rect 277398 597744 312970 597800
rect 313026 597744 313094 597800
rect 313150 597744 313218 597800
rect 313274 597744 313342 597800
rect 313398 597744 330970 597800
rect 331026 597744 331094 597800
rect 331150 597744 331218 597800
rect 331274 597744 331342 597800
rect 331398 597744 348970 597800
rect 349026 597744 349094 597800
rect 349150 597744 349218 597800
rect 349274 597744 349342 597800
rect 349398 597744 366970 597800
rect 367026 597744 367094 597800
rect 367150 597744 367218 597800
rect 367274 597744 367342 597800
rect 367398 597744 402970 597800
rect 403026 597744 403094 597800
rect 403150 597744 403218 597800
rect 403274 597744 403342 597800
rect 403398 597744 420970 597800
rect 421026 597744 421094 597800
rect 421150 597744 421218 597800
rect 421274 597744 421342 597800
rect 421398 597744 438970 597800
rect 439026 597744 439094 597800
rect 439150 597744 439218 597800
rect 439274 597744 439342 597800
rect 439398 597744 456970 597800
rect 457026 597744 457094 597800
rect 457150 597744 457218 597800
rect 457274 597744 457342 597800
rect 457398 597744 492970 597800
rect 493026 597744 493094 597800
rect 493150 597744 493218 597800
rect 493274 597744 493342 597800
rect 493398 597744 510970 597800
rect 511026 597744 511094 597800
rect 511150 597744 511218 597800
rect 511274 597744 511342 597800
rect 511398 597744 528970 597800
rect 529026 597744 529094 597800
rect 529150 597744 529218 597800
rect 529274 597744 529342 597800
rect 529398 597744 546970 597800
rect 547026 597744 547094 597800
rect 547150 597744 547218 597800
rect 547274 597744 547342 597800
rect 547398 597744 564970 597800
rect 565026 597744 565094 597800
rect 565150 597744 565218 597800
rect 565274 597744 565342 597800
rect 565398 597744 582970 597800
rect 583026 597744 583094 597800
rect 583150 597744 583218 597800
rect 583274 597744 583342 597800
rect 583398 597744 597456 597800
rect 597512 597744 597580 597800
rect 597636 597744 597704 597800
rect 597760 597744 597828 597800
rect 597884 597744 597980 597800
rect -1916 597648 597980 597744
rect -956 597212 597020 597308
rect -956 597156 -860 597212
rect -804 597156 -736 597212
rect -680 597156 -612 597212
rect -556 597156 -488 597212
rect -432 597156 3250 597212
rect 3306 597156 3374 597212
rect 3430 597156 3498 597212
rect 3554 597156 3622 597212
rect 3678 597156 21250 597212
rect 21306 597156 21374 597212
rect 21430 597156 21498 597212
rect 21554 597156 21622 597212
rect 21678 597156 39250 597212
rect 39306 597156 39374 597212
rect 39430 597156 39498 597212
rect 39554 597156 39622 597212
rect 39678 597156 57250 597212
rect 57306 597156 57374 597212
rect 57430 597156 57498 597212
rect 57554 597156 57622 597212
rect 57678 597156 93250 597212
rect 93306 597156 93374 597212
rect 93430 597156 93498 597212
rect 93554 597156 93622 597212
rect 93678 597156 111250 597212
rect 111306 597156 111374 597212
rect 111430 597156 111498 597212
rect 111554 597156 111622 597212
rect 111678 597156 129250 597212
rect 129306 597156 129374 597212
rect 129430 597156 129498 597212
rect 129554 597156 129622 597212
rect 129678 597156 147250 597212
rect 147306 597156 147374 597212
rect 147430 597156 147498 597212
rect 147554 597156 147622 597212
rect 147678 597156 183250 597212
rect 183306 597156 183374 597212
rect 183430 597156 183498 597212
rect 183554 597156 183622 597212
rect 183678 597156 201250 597212
rect 201306 597156 201374 597212
rect 201430 597156 201498 597212
rect 201554 597156 201622 597212
rect 201678 597156 219250 597212
rect 219306 597156 219374 597212
rect 219430 597156 219498 597212
rect 219554 597156 219622 597212
rect 219678 597156 237250 597212
rect 237306 597156 237374 597212
rect 237430 597156 237498 597212
rect 237554 597156 237622 597212
rect 237678 597156 273250 597212
rect 273306 597156 273374 597212
rect 273430 597156 273498 597212
rect 273554 597156 273622 597212
rect 273678 597156 291250 597212
rect 291306 597156 291374 597212
rect 291430 597156 291498 597212
rect 291554 597156 291622 597212
rect 291678 597156 309250 597212
rect 309306 597156 309374 597212
rect 309430 597156 309498 597212
rect 309554 597156 309622 597212
rect 309678 597156 327250 597212
rect 327306 597156 327374 597212
rect 327430 597156 327498 597212
rect 327554 597156 327622 597212
rect 327678 597156 363250 597212
rect 363306 597156 363374 597212
rect 363430 597156 363498 597212
rect 363554 597156 363622 597212
rect 363678 597156 381250 597212
rect 381306 597156 381374 597212
rect 381430 597156 381498 597212
rect 381554 597156 381622 597212
rect 381678 597156 399250 597212
rect 399306 597156 399374 597212
rect 399430 597156 399498 597212
rect 399554 597156 399622 597212
rect 399678 597156 417250 597212
rect 417306 597156 417374 597212
rect 417430 597156 417498 597212
rect 417554 597156 417622 597212
rect 417678 597156 453250 597212
rect 453306 597156 453374 597212
rect 453430 597156 453498 597212
rect 453554 597156 453622 597212
rect 453678 597156 471250 597212
rect 471306 597156 471374 597212
rect 471430 597156 471498 597212
rect 471554 597156 471622 597212
rect 471678 597156 489250 597212
rect 489306 597156 489374 597212
rect 489430 597156 489498 597212
rect 489554 597156 489622 597212
rect 489678 597156 507250 597212
rect 507306 597156 507374 597212
rect 507430 597156 507498 597212
rect 507554 597156 507622 597212
rect 507678 597156 543250 597212
rect 543306 597156 543374 597212
rect 543430 597156 543498 597212
rect 543554 597156 543622 597212
rect 543678 597156 561250 597212
rect 561306 597156 561374 597212
rect 561430 597156 561498 597212
rect 561554 597156 561622 597212
rect 561678 597156 579250 597212
rect 579306 597156 579374 597212
rect 579430 597156 579498 597212
rect 579554 597156 579622 597212
rect 579678 597156 596496 597212
rect 596552 597156 596620 597212
rect 596676 597156 596744 597212
rect 596800 597156 596868 597212
rect 596924 597156 597020 597212
rect -956 597088 597020 597156
rect -956 597032 -860 597088
rect -804 597032 -736 597088
rect -680 597032 -612 597088
rect -556 597032 -488 597088
rect -432 597032 3250 597088
rect 3306 597032 3374 597088
rect 3430 597032 3498 597088
rect 3554 597032 3622 597088
rect 3678 597032 21250 597088
rect 21306 597032 21374 597088
rect 21430 597032 21498 597088
rect 21554 597032 21622 597088
rect 21678 597032 39250 597088
rect 39306 597032 39374 597088
rect 39430 597032 39498 597088
rect 39554 597032 39622 597088
rect 39678 597032 57250 597088
rect 57306 597032 57374 597088
rect 57430 597032 57498 597088
rect 57554 597032 57622 597088
rect 57678 597032 93250 597088
rect 93306 597032 93374 597088
rect 93430 597032 93498 597088
rect 93554 597032 93622 597088
rect 93678 597032 111250 597088
rect 111306 597032 111374 597088
rect 111430 597032 111498 597088
rect 111554 597032 111622 597088
rect 111678 597032 129250 597088
rect 129306 597032 129374 597088
rect 129430 597032 129498 597088
rect 129554 597032 129622 597088
rect 129678 597032 147250 597088
rect 147306 597032 147374 597088
rect 147430 597032 147498 597088
rect 147554 597032 147622 597088
rect 147678 597032 183250 597088
rect 183306 597032 183374 597088
rect 183430 597032 183498 597088
rect 183554 597032 183622 597088
rect 183678 597032 201250 597088
rect 201306 597032 201374 597088
rect 201430 597032 201498 597088
rect 201554 597032 201622 597088
rect 201678 597032 219250 597088
rect 219306 597032 219374 597088
rect 219430 597032 219498 597088
rect 219554 597032 219622 597088
rect 219678 597032 237250 597088
rect 237306 597032 237374 597088
rect 237430 597032 237498 597088
rect 237554 597032 237622 597088
rect 237678 597032 273250 597088
rect 273306 597032 273374 597088
rect 273430 597032 273498 597088
rect 273554 597032 273622 597088
rect 273678 597032 291250 597088
rect 291306 597032 291374 597088
rect 291430 597032 291498 597088
rect 291554 597032 291622 597088
rect 291678 597032 309250 597088
rect 309306 597032 309374 597088
rect 309430 597032 309498 597088
rect 309554 597032 309622 597088
rect 309678 597032 327250 597088
rect 327306 597032 327374 597088
rect 327430 597032 327498 597088
rect 327554 597032 327622 597088
rect 327678 597032 363250 597088
rect 363306 597032 363374 597088
rect 363430 597032 363498 597088
rect 363554 597032 363622 597088
rect 363678 597032 381250 597088
rect 381306 597032 381374 597088
rect 381430 597032 381498 597088
rect 381554 597032 381622 597088
rect 381678 597032 399250 597088
rect 399306 597032 399374 597088
rect 399430 597032 399498 597088
rect 399554 597032 399622 597088
rect 399678 597032 417250 597088
rect 417306 597032 417374 597088
rect 417430 597032 417498 597088
rect 417554 597032 417622 597088
rect 417678 597032 453250 597088
rect 453306 597032 453374 597088
rect 453430 597032 453498 597088
rect 453554 597032 453622 597088
rect 453678 597032 471250 597088
rect 471306 597032 471374 597088
rect 471430 597032 471498 597088
rect 471554 597032 471622 597088
rect 471678 597032 489250 597088
rect 489306 597032 489374 597088
rect 489430 597032 489498 597088
rect 489554 597032 489622 597088
rect 489678 597032 507250 597088
rect 507306 597032 507374 597088
rect 507430 597032 507498 597088
rect 507554 597032 507622 597088
rect 507678 597032 543250 597088
rect 543306 597032 543374 597088
rect 543430 597032 543498 597088
rect 543554 597032 543622 597088
rect 543678 597032 561250 597088
rect 561306 597032 561374 597088
rect 561430 597032 561498 597088
rect 561554 597032 561622 597088
rect 561678 597032 579250 597088
rect 579306 597032 579374 597088
rect 579430 597032 579498 597088
rect 579554 597032 579622 597088
rect 579678 597032 596496 597088
rect 596552 597032 596620 597088
rect 596676 597032 596744 597088
rect 596800 597032 596868 597088
rect 596924 597032 597020 597088
rect -956 596964 597020 597032
rect -956 596908 -860 596964
rect -804 596908 -736 596964
rect -680 596908 -612 596964
rect -556 596908 -488 596964
rect -432 596908 3250 596964
rect 3306 596908 3374 596964
rect 3430 596908 3498 596964
rect 3554 596908 3622 596964
rect 3678 596908 21250 596964
rect 21306 596908 21374 596964
rect 21430 596908 21498 596964
rect 21554 596908 21622 596964
rect 21678 596908 39250 596964
rect 39306 596908 39374 596964
rect 39430 596908 39498 596964
rect 39554 596908 39622 596964
rect 39678 596908 57250 596964
rect 57306 596908 57374 596964
rect 57430 596908 57498 596964
rect 57554 596908 57622 596964
rect 57678 596908 93250 596964
rect 93306 596908 93374 596964
rect 93430 596908 93498 596964
rect 93554 596908 93622 596964
rect 93678 596908 111250 596964
rect 111306 596908 111374 596964
rect 111430 596908 111498 596964
rect 111554 596908 111622 596964
rect 111678 596908 129250 596964
rect 129306 596908 129374 596964
rect 129430 596908 129498 596964
rect 129554 596908 129622 596964
rect 129678 596908 147250 596964
rect 147306 596908 147374 596964
rect 147430 596908 147498 596964
rect 147554 596908 147622 596964
rect 147678 596908 183250 596964
rect 183306 596908 183374 596964
rect 183430 596908 183498 596964
rect 183554 596908 183622 596964
rect 183678 596908 201250 596964
rect 201306 596908 201374 596964
rect 201430 596908 201498 596964
rect 201554 596908 201622 596964
rect 201678 596908 219250 596964
rect 219306 596908 219374 596964
rect 219430 596908 219498 596964
rect 219554 596908 219622 596964
rect 219678 596908 237250 596964
rect 237306 596908 237374 596964
rect 237430 596908 237498 596964
rect 237554 596908 237622 596964
rect 237678 596908 273250 596964
rect 273306 596908 273374 596964
rect 273430 596908 273498 596964
rect 273554 596908 273622 596964
rect 273678 596908 291250 596964
rect 291306 596908 291374 596964
rect 291430 596908 291498 596964
rect 291554 596908 291622 596964
rect 291678 596908 309250 596964
rect 309306 596908 309374 596964
rect 309430 596908 309498 596964
rect 309554 596908 309622 596964
rect 309678 596908 327250 596964
rect 327306 596908 327374 596964
rect 327430 596908 327498 596964
rect 327554 596908 327622 596964
rect 327678 596908 363250 596964
rect 363306 596908 363374 596964
rect 363430 596908 363498 596964
rect 363554 596908 363622 596964
rect 363678 596908 381250 596964
rect 381306 596908 381374 596964
rect 381430 596908 381498 596964
rect 381554 596908 381622 596964
rect 381678 596908 399250 596964
rect 399306 596908 399374 596964
rect 399430 596908 399498 596964
rect 399554 596908 399622 596964
rect 399678 596908 417250 596964
rect 417306 596908 417374 596964
rect 417430 596908 417498 596964
rect 417554 596908 417622 596964
rect 417678 596908 453250 596964
rect 453306 596908 453374 596964
rect 453430 596908 453498 596964
rect 453554 596908 453622 596964
rect 453678 596908 471250 596964
rect 471306 596908 471374 596964
rect 471430 596908 471498 596964
rect 471554 596908 471622 596964
rect 471678 596908 489250 596964
rect 489306 596908 489374 596964
rect 489430 596908 489498 596964
rect 489554 596908 489622 596964
rect 489678 596908 507250 596964
rect 507306 596908 507374 596964
rect 507430 596908 507498 596964
rect 507554 596908 507622 596964
rect 507678 596908 543250 596964
rect 543306 596908 543374 596964
rect 543430 596908 543498 596964
rect 543554 596908 543622 596964
rect 543678 596908 561250 596964
rect 561306 596908 561374 596964
rect 561430 596908 561498 596964
rect 561554 596908 561622 596964
rect 561678 596908 579250 596964
rect 579306 596908 579374 596964
rect 579430 596908 579498 596964
rect 579554 596908 579622 596964
rect 579678 596908 596496 596964
rect 596552 596908 596620 596964
rect 596676 596908 596744 596964
rect 596800 596908 596868 596964
rect 596924 596908 597020 596964
rect -956 596840 597020 596908
rect -956 596784 -860 596840
rect -804 596784 -736 596840
rect -680 596784 -612 596840
rect -556 596784 -488 596840
rect -432 596784 3250 596840
rect 3306 596784 3374 596840
rect 3430 596784 3498 596840
rect 3554 596784 3622 596840
rect 3678 596784 21250 596840
rect 21306 596784 21374 596840
rect 21430 596784 21498 596840
rect 21554 596784 21622 596840
rect 21678 596784 39250 596840
rect 39306 596784 39374 596840
rect 39430 596784 39498 596840
rect 39554 596784 39622 596840
rect 39678 596784 57250 596840
rect 57306 596784 57374 596840
rect 57430 596784 57498 596840
rect 57554 596784 57622 596840
rect 57678 596784 93250 596840
rect 93306 596784 93374 596840
rect 93430 596784 93498 596840
rect 93554 596784 93622 596840
rect 93678 596784 111250 596840
rect 111306 596784 111374 596840
rect 111430 596784 111498 596840
rect 111554 596784 111622 596840
rect 111678 596784 129250 596840
rect 129306 596784 129374 596840
rect 129430 596784 129498 596840
rect 129554 596784 129622 596840
rect 129678 596784 147250 596840
rect 147306 596784 147374 596840
rect 147430 596784 147498 596840
rect 147554 596784 147622 596840
rect 147678 596784 183250 596840
rect 183306 596784 183374 596840
rect 183430 596784 183498 596840
rect 183554 596784 183622 596840
rect 183678 596784 201250 596840
rect 201306 596784 201374 596840
rect 201430 596784 201498 596840
rect 201554 596784 201622 596840
rect 201678 596784 219250 596840
rect 219306 596784 219374 596840
rect 219430 596784 219498 596840
rect 219554 596784 219622 596840
rect 219678 596784 237250 596840
rect 237306 596784 237374 596840
rect 237430 596784 237498 596840
rect 237554 596784 237622 596840
rect 237678 596784 273250 596840
rect 273306 596784 273374 596840
rect 273430 596784 273498 596840
rect 273554 596784 273622 596840
rect 273678 596784 291250 596840
rect 291306 596784 291374 596840
rect 291430 596784 291498 596840
rect 291554 596784 291622 596840
rect 291678 596784 309250 596840
rect 309306 596784 309374 596840
rect 309430 596784 309498 596840
rect 309554 596784 309622 596840
rect 309678 596784 327250 596840
rect 327306 596784 327374 596840
rect 327430 596784 327498 596840
rect 327554 596784 327622 596840
rect 327678 596784 363250 596840
rect 363306 596784 363374 596840
rect 363430 596784 363498 596840
rect 363554 596784 363622 596840
rect 363678 596784 381250 596840
rect 381306 596784 381374 596840
rect 381430 596784 381498 596840
rect 381554 596784 381622 596840
rect 381678 596784 399250 596840
rect 399306 596784 399374 596840
rect 399430 596784 399498 596840
rect 399554 596784 399622 596840
rect 399678 596784 417250 596840
rect 417306 596784 417374 596840
rect 417430 596784 417498 596840
rect 417554 596784 417622 596840
rect 417678 596784 453250 596840
rect 453306 596784 453374 596840
rect 453430 596784 453498 596840
rect 453554 596784 453622 596840
rect 453678 596784 471250 596840
rect 471306 596784 471374 596840
rect 471430 596784 471498 596840
rect 471554 596784 471622 596840
rect 471678 596784 489250 596840
rect 489306 596784 489374 596840
rect 489430 596784 489498 596840
rect 489554 596784 489622 596840
rect 489678 596784 507250 596840
rect 507306 596784 507374 596840
rect 507430 596784 507498 596840
rect 507554 596784 507622 596840
rect 507678 596784 543250 596840
rect 543306 596784 543374 596840
rect 543430 596784 543498 596840
rect 543554 596784 543622 596840
rect 543678 596784 561250 596840
rect 561306 596784 561374 596840
rect 561430 596784 561498 596840
rect 561554 596784 561622 596840
rect 561678 596784 579250 596840
rect 579306 596784 579374 596840
rect 579430 596784 579498 596840
rect 579554 596784 579622 596840
rect 579678 596784 596496 596840
rect 596552 596784 596620 596840
rect 596676 596784 596744 596840
rect 596800 596784 596868 596840
rect 596924 596784 597020 596840
rect -956 596688 597020 596784
rect -1916 586350 597980 586446
rect -1916 586294 -1820 586350
rect -1764 586294 -1696 586350
rect -1640 586294 -1572 586350
rect -1516 586294 -1448 586350
rect -1392 586294 6970 586350
rect 7026 586294 7094 586350
rect 7150 586294 7218 586350
rect 7274 586294 7342 586350
rect 7398 586294 24970 586350
rect 25026 586294 25094 586350
rect 25150 586294 25218 586350
rect 25274 586294 25342 586350
rect 25398 586294 42970 586350
rect 43026 586294 43094 586350
rect 43150 586294 43218 586350
rect 43274 586294 43342 586350
rect 43398 586294 60970 586350
rect 61026 586294 61094 586350
rect 61150 586294 61218 586350
rect 61274 586294 61342 586350
rect 61398 586294 78970 586350
rect 79026 586294 79094 586350
rect 79150 586294 79218 586350
rect 79274 586294 79342 586350
rect 79398 586294 96970 586350
rect 97026 586294 97094 586350
rect 97150 586294 97218 586350
rect 97274 586294 97342 586350
rect 97398 586294 132970 586350
rect 133026 586294 133094 586350
rect 133150 586294 133218 586350
rect 133274 586294 133342 586350
rect 133398 586294 150970 586350
rect 151026 586294 151094 586350
rect 151150 586294 151218 586350
rect 151274 586294 151342 586350
rect 151398 586294 168970 586350
rect 169026 586294 169094 586350
rect 169150 586294 169218 586350
rect 169274 586294 169342 586350
rect 169398 586294 186970 586350
rect 187026 586294 187094 586350
rect 187150 586294 187218 586350
rect 187274 586294 187342 586350
rect 187398 586294 222970 586350
rect 223026 586294 223094 586350
rect 223150 586294 223218 586350
rect 223274 586294 223342 586350
rect 223398 586294 240970 586350
rect 241026 586294 241094 586350
rect 241150 586294 241218 586350
rect 241274 586294 241342 586350
rect 241398 586294 258970 586350
rect 259026 586294 259094 586350
rect 259150 586294 259218 586350
rect 259274 586294 259342 586350
rect 259398 586294 276970 586350
rect 277026 586294 277094 586350
rect 277150 586294 277218 586350
rect 277274 586294 277342 586350
rect 277398 586294 312970 586350
rect 313026 586294 313094 586350
rect 313150 586294 313218 586350
rect 313274 586294 313342 586350
rect 313398 586294 330970 586350
rect 331026 586294 331094 586350
rect 331150 586294 331218 586350
rect 331274 586294 331342 586350
rect 331398 586294 348970 586350
rect 349026 586294 349094 586350
rect 349150 586294 349218 586350
rect 349274 586294 349342 586350
rect 349398 586294 366970 586350
rect 367026 586294 367094 586350
rect 367150 586294 367218 586350
rect 367274 586294 367342 586350
rect 367398 586294 402970 586350
rect 403026 586294 403094 586350
rect 403150 586294 403218 586350
rect 403274 586294 403342 586350
rect 403398 586294 420970 586350
rect 421026 586294 421094 586350
rect 421150 586294 421218 586350
rect 421274 586294 421342 586350
rect 421398 586294 438970 586350
rect 439026 586294 439094 586350
rect 439150 586294 439218 586350
rect 439274 586294 439342 586350
rect 439398 586294 456970 586350
rect 457026 586294 457094 586350
rect 457150 586294 457218 586350
rect 457274 586294 457342 586350
rect 457398 586294 492970 586350
rect 493026 586294 493094 586350
rect 493150 586294 493218 586350
rect 493274 586294 493342 586350
rect 493398 586294 510970 586350
rect 511026 586294 511094 586350
rect 511150 586294 511218 586350
rect 511274 586294 511342 586350
rect 511398 586294 528970 586350
rect 529026 586294 529094 586350
rect 529150 586294 529218 586350
rect 529274 586294 529342 586350
rect 529398 586294 546970 586350
rect 547026 586294 547094 586350
rect 547150 586294 547218 586350
rect 547274 586294 547342 586350
rect 547398 586294 564970 586350
rect 565026 586294 565094 586350
rect 565150 586294 565218 586350
rect 565274 586294 565342 586350
rect 565398 586294 582970 586350
rect 583026 586294 583094 586350
rect 583150 586294 583218 586350
rect 583274 586294 583342 586350
rect 583398 586294 597456 586350
rect 597512 586294 597580 586350
rect 597636 586294 597704 586350
rect 597760 586294 597828 586350
rect 597884 586294 597980 586350
rect -1916 586226 597980 586294
rect -1916 586170 -1820 586226
rect -1764 586170 -1696 586226
rect -1640 586170 -1572 586226
rect -1516 586170 -1448 586226
rect -1392 586170 6970 586226
rect 7026 586170 7094 586226
rect 7150 586170 7218 586226
rect 7274 586170 7342 586226
rect 7398 586170 24970 586226
rect 25026 586170 25094 586226
rect 25150 586170 25218 586226
rect 25274 586170 25342 586226
rect 25398 586170 42970 586226
rect 43026 586170 43094 586226
rect 43150 586170 43218 586226
rect 43274 586170 43342 586226
rect 43398 586170 60970 586226
rect 61026 586170 61094 586226
rect 61150 586170 61218 586226
rect 61274 586170 61342 586226
rect 61398 586170 78970 586226
rect 79026 586170 79094 586226
rect 79150 586170 79218 586226
rect 79274 586170 79342 586226
rect 79398 586170 96970 586226
rect 97026 586170 97094 586226
rect 97150 586170 97218 586226
rect 97274 586170 97342 586226
rect 97398 586170 132970 586226
rect 133026 586170 133094 586226
rect 133150 586170 133218 586226
rect 133274 586170 133342 586226
rect 133398 586170 150970 586226
rect 151026 586170 151094 586226
rect 151150 586170 151218 586226
rect 151274 586170 151342 586226
rect 151398 586170 168970 586226
rect 169026 586170 169094 586226
rect 169150 586170 169218 586226
rect 169274 586170 169342 586226
rect 169398 586170 186970 586226
rect 187026 586170 187094 586226
rect 187150 586170 187218 586226
rect 187274 586170 187342 586226
rect 187398 586170 222970 586226
rect 223026 586170 223094 586226
rect 223150 586170 223218 586226
rect 223274 586170 223342 586226
rect 223398 586170 240970 586226
rect 241026 586170 241094 586226
rect 241150 586170 241218 586226
rect 241274 586170 241342 586226
rect 241398 586170 258970 586226
rect 259026 586170 259094 586226
rect 259150 586170 259218 586226
rect 259274 586170 259342 586226
rect 259398 586170 276970 586226
rect 277026 586170 277094 586226
rect 277150 586170 277218 586226
rect 277274 586170 277342 586226
rect 277398 586170 312970 586226
rect 313026 586170 313094 586226
rect 313150 586170 313218 586226
rect 313274 586170 313342 586226
rect 313398 586170 330970 586226
rect 331026 586170 331094 586226
rect 331150 586170 331218 586226
rect 331274 586170 331342 586226
rect 331398 586170 348970 586226
rect 349026 586170 349094 586226
rect 349150 586170 349218 586226
rect 349274 586170 349342 586226
rect 349398 586170 366970 586226
rect 367026 586170 367094 586226
rect 367150 586170 367218 586226
rect 367274 586170 367342 586226
rect 367398 586170 402970 586226
rect 403026 586170 403094 586226
rect 403150 586170 403218 586226
rect 403274 586170 403342 586226
rect 403398 586170 420970 586226
rect 421026 586170 421094 586226
rect 421150 586170 421218 586226
rect 421274 586170 421342 586226
rect 421398 586170 438970 586226
rect 439026 586170 439094 586226
rect 439150 586170 439218 586226
rect 439274 586170 439342 586226
rect 439398 586170 456970 586226
rect 457026 586170 457094 586226
rect 457150 586170 457218 586226
rect 457274 586170 457342 586226
rect 457398 586170 492970 586226
rect 493026 586170 493094 586226
rect 493150 586170 493218 586226
rect 493274 586170 493342 586226
rect 493398 586170 510970 586226
rect 511026 586170 511094 586226
rect 511150 586170 511218 586226
rect 511274 586170 511342 586226
rect 511398 586170 528970 586226
rect 529026 586170 529094 586226
rect 529150 586170 529218 586226
rect 529274 586170 529342 586226
rect 529398 586170 546970 586226
rect 547026 586170 547094 586226
rect 547150 586170 547218 586226
rect 547274 586170 547342 586226
rect 547398 586170 564970 586226
rect 565026 586170 565094 586226
rect 565150 586170 565218 586226
rect 565274 586170 565342 586226
rect 565398 586170 582970 586226
rect 583026 586170 583094 586226
rect 583150 586170 583218 586226
rect 583274 586170 583342 586226
rect 583398 586170 597456 586226
rect 597512 586170 597580 586226
rect 597636 586170 597704 586226
rect 597760 586170 597828 586226
rect 597884 586170 597980 586226
rect -1916 586102 597980 586170
rect -1916 586046 -1820 586102
rect -1764 586046 -1696 586102
rect -1640 586046 -1572 586102
rect -1516 586046 -1448 586102
rect -1392 586046 6970 586102
rect 7026 586046 7094 586102
rect 7150 586046 7218 586102
rect 7274 586046 7342 586102
rect 7398 586046 24970 586102
rect 25026 586046 25094 586102
rect 25150 586046 25218 586102
rect 25274 586046 25342 586102
rect 25398 586046 42970 586102
rect 43026 586046 43094 586102
rect 43150 586046 43218 586102
rect 43274 586046 43342 586102
rect 43398 586046 60970 586102
rect 61026 586046 61094 586102
rect 61150 586046 61218 586102
rect 61274 586046 61342 586102
rect 61398 586046 78970 586102
rect 79026 586046 79094 586102
rect 79150 586046 79218 586102
rect 79274 586046 79342 586102
rect 79398 586046 96970 586102
rect 97026 586046 97094 586102
rect 97150 586046 97218 586102
rect 97274 586046 97342 586102
rect 97398 586046 132970 586102
rect 133026 586046 133094 586102
rect 133150 586046 133218 586102
rect 133274 586046 133342 586102
rect 133398 586046 150970 586102
rect 151026 586046 151094 586102
rect 151150 586046 151218 586102
rect 151274 586046 151342 586102
rect 151398 586046 168970 586102
rect 169026 586046 169094 586102
rect 169150 586046 169218 586102
rect 169274 586046 169342 586102
rect 169398 586046 186970 586102
rect 187026 586046 187094 586102
rect 187150 586046 187218 586102
rect 187274 586046 187342 586102
rect 187398 586046 222970 586102
rect 223026 586046 223094 586102
rect 223150 586046 223218 586102
rect 223274 586046 223342 586102
rect 223398 586046 240970 586102
rect 241026 586046 241094 586102
rect 241150 586046 241218 586102
rect 241274 586046 241342 586102
rect 241398 586046 258970 586102
rect 259026 586046 259094 586102
rect 259150 586046 259218 586102
rect 259274 586046 259342 586102
rect 259398 586046 276970 586102
rect 277026 586046 277094 586102
rect 277150 586046 277218 586102
rect 277274 586046 277342 586102
rect 277398 586046 312970 586102
rect 313026 586046 313094 586102
rect 313150 586046 313218 586102
rect 313274 586046 313342 586102
rect 313398 586046 330970 586102
rect 331026 586046 331094 586102
rect 331150 586046 331218 586102
rect 331274 586046 331342 586102
rect 331398 586046 348970 586102
rect 349026 586046 349094 586102
rect 349150 586046 349218 586102
rect 349274 586046 349342 586102
rect 349398 586046 366970 586102
rect 367026 586046 367094 586102
rect 367150 586046 367218 586102
rect 367274 586046 367342 586102
rect 367398 586046 402970 586102
rect 403026 586046 403094 586102
rect 403150 586046 403218 586102
rect 403274 586046 403342 586102
rect 403398 586046 420970 586102
rect 421026 586046 421094 586102
rect 421150 586046 421218 586102
rect 421274 586046 421342 586102
rect 421398 586046 438970 586102
rect 439026 586046 439094 586102
rect 439150 586046 439218 586102
rect 439274 586046 439342 586102
rect 439398 586046 456970 586102
rect 457026 586046 457094 586102
rect 457150 586046 457218 586102
rect 457274 586046 457342 586102
rect 457398 586046 492970 586102
rect 493026 586046 493094 586102
rect 493150 586046 493218 586102
rect 493274 586046 493342 586102
rect 493398 586046 510970 586102
rect 511026 586046 511094 586102
rect 511150 586046 511218 586102
rect 511274 586046 511342 586102
rect 511398 586046 528970 586102
rect 529026 586046 529094 586102
rect 529150 586046 529218 586102
rect 529274 586046 529342 586102
rect 529398 586046 546970 586102
rect 547026 586046 547094 586102
rect 547150 586046 547218 586102
rect 547274 586046 547342 586102
rect 547398 586046 564970 586102
rect 565026 586046 565094 586102
rect 565150 586046 565218 586102
rect 565274 586046 565342 586102
rect 565398 586046 582970 586102
rect 583026 586046 583094 586102
rect 583150 586046 583218 586102
rect 583274 586046 583342 586102
rect 583398 586046 597456 586102
rect 597512 586046 597580 586102
rect 597636 586046 597704 586102
rect 597760 586046 597828 586102
rect 597884 586046 597980 586102
rect -1916 585978 597980 586046
rect -1916 585922 -1820 585978
rect -1764 585922 -1696 585978
rect -1640 585922 -1572 585978
rect -1516 585922 -1448 585978
rect -1392 585922 6970 585978
rect 7026 585922 7094 585978
rect 7150 585922 7218 585978
rect 7274 585922 7342 585978
rect 7398 585922 24970 585978
rect 25026 585922 25094 585978
rect 25150 585922 25218 585978
rect 25274 585922 25342 585978
rect 25398 585922 42970 585978
rect 43026 585922 43094 585978
rect 43150 585922 43218 585978
rect 43274 585922 43342 585978
rect 43398 585922 60970 585978
rect 61026 585922 61094 585978
rect 61150 585922 61218 585978
rect 61274 585922 61342 585978
rect 61398 585922 78970 585978
rect 79026 585922 79094 585978
rect 79150 585922 79218 585978
rect 79274 585922 79342 585978
rect 79398 585922 96970 585978
rect 97026 585922 97094 585978
rect 97150 585922 97218 585978
rect 97274 585922 97342 585978
rect 97398 585922 132970 585978
rect 133026 585922 133094 585978
rect 133150 585922 133218 585978
rect 133274 585922 133342 585978
rect 133398 585922 150970 585978
rect 151026 585922 151094 585978
rect 151150 585922 151218 585978
rect 151274 585922 151342 585978
rect 151398 585922 168970 585978
rect 169026 585922 169094 585978
rect 169150 585922 169218 585978
rect 169274 585922 169342 585978
rect 169398 585922 186970 585978
rect 187026 585922 187094 585978
rect 187150 585922 187218 585978
rect 187274 585922 187342 585978
rect 187398 585922 222970 585978
rect 223026 585922 223094 585978
rect 223150 585922 223218 585978
rect 223274 585922 223342 585978
rect 223398 585922 240970 585978
rect 241026 585922 241094 585978
rect 241150 585922 241218 585978
rect 241274 585922 241342 585978
rect 241398 585922 258970 585978
rect 259026 585922 259094 585978
rect 259150 585922 259218 585978
rect 259274 585922 259342 585978
rect 259398 585922 276970 585978
rect 277026 585922 277094 585978
rect 277150 585922 277218 585978
rect 277274 585922 277342 585978
rect 277398 585922 312970 585978
rect 313026 585922 313094 585978
rect 313150 585922 313218 585978
rect 313274 585922 313342 585978
rect 313398 585922 330970 585978
rect 331026 585922 331094 585978
rect 331150 585922 331218 585978
rect 331274 585922 331342 585978
rect 331398 585922 348970 585978
rect 349026 585922 349094 585978
rect 349150 585922 349218 585978
rect 349274 585922 349342 585978
rect 349398 585922 366970 585978
rect 367026 585922 367094 585978
rect 367150 585922 367218 585978
rect 367274 585922 367342 585978
rect 367398 585922 402970 585978
rect 403026 585922 403094 585978
rect 403150 585922 403218 585978
rect 403274 585922 403342 585978
rect 403398 585922 420970 585978
rect 421026 585922 421094 585978
rect 421150 585922 421218 585978
rect 421274 585922 421342 585978
rect 421398 585922 438970 585978
rect 439026 585922 439094 585978
rect 439150 585922 439218 585978
rect 439274 585922 439342 585978
rect 439398 585922 456970 585978
rect 457026 585922 457094 585978
rect 457150 585922 457218 585978
rect 457274 585922 457342 585978
rect 457398 585922 492970 585978
rect 493026 585922 493094 585978
rect 493150 585922 493218 585978
rect 493274 585922 493342 585978
rect 493398 585922 510970 585978
rect 511026 585922 511094 585978
rect 511150 585922 511218 585978
rect 511274 585922 511342 585978
rect 511398 585922 528970 585978
rect 529026 585922 529094 585978
rect 529150 585922 529218 585978
rect 529274 585922 529342 585978
rect 529398 585922 546970 585978
rect 547026 585922 547094 585978
rect 547150 585922 547218 585978
rect 547274 585922 547342 585978
rect 547398 585922 564970 585978
rect 565026 585922 565094 585978
rect 565150 585922 565218 585978
rect 565274 585922 565342 585978
rect 565398 585922 582970 585978
rect 583026 585922 583094 585978
rect 583150 585922 583218 585978
rect 583274 585922 583342 585978
rect 583398 585922 597456 585978
rect 597512 585922 597580 585978
rect 597636 585922 597704 585978
rect 597760 585922 597828 585978
rect 597884 585922 597980 585978
rect -1916 585826 597980 585922
rect -1916 580350 597980 580446
rect -1916 580294 -860 580350
rect -804 580294 -736 580350
rect -680 580294 -612 580350
rect -556 580294 -488 580350
rect -432 580294 3250 580350
rect 3306 580294 3374 580350
rect 3430 580294 3498 580350
rect 3554 580294 3622 580350
rect 3678 580294 21250 580350
rect 21306 580294 21374 580350
rect 21430 580294 21498 580350
rect 21554 580294 21622 580350
rect 21678 580294 39250 580350
rect 39306 580294 39374 580350
rect 39430 580294 39498 580350
rect 39554 580294 39622 580350
rect 39678 580294 57250 580350
rect 57306 580294 57374 580350
rect 57430 580294 57498 580350
rect 57554 580294 57622 580350
rect 57678 580294 93250 580350
rect 93306 580294 93374 580350
rect 93430 580294 93498 580350
rect 93554 580294 93622 580350
rect 93678 580294 111250 580350
rect 111306 580294 111374 580350
rect 111430 580294 111498 580350
rect 111554 580294 111622 580350
rect 111678 580294 129250 580350
rect 129306 580294 129374 580350
rect 129430 580294 129498 580350
rect 129554 580294 129622 580350
rect 129678 580294 147250 580350
rect 147306 580294 147374 580350
rect 147430 580294 147498 580350
rect 147554 580294 147622 580350
rect 147678 580294 183250 580350
rect 183306 580294 183374 580350
rect 183430 580294 183498 580350
rect 183554 580294 183622 580350
rect 183678 580294 201250 580350
rect 201306 580294 201374 580350
rect 201430 580294 201498 580350
rect 201554 580294 201622 580350
rect 201678 580294 219250 580350
rect 219306 580294 219374 580350
rect 219430 580294 219498 580350
rect 219554 580294 219622 580350
rect 219678 580294 237250 580350
rect 237306 580294 237374 580350
rect 237430 580294 237498 580350
rect 237554 580294 237622 580350
rect 237678 580294 273250 580350
rect 273306 580294 273374 580350
rect 273430 580294 273498 580350
rect 273554 580294 273622 580350
rect 273678 580294 291250 580350
rect 291306 580294 291374 580350
rect 291430 580294 291498 580350
rect 291554 580294 291622 580350
rect 291678 580294 309250 580350
rect 309306 580294 309374 580350
rect 309430 580294 309498 580350
rect 309554 580294 309622 580350
rect 309678 580294 327250 580350
rect 327306 580294 327374 580350
rect 327430 580294 327498 580350
rect 327554 580294 327622 580350
rect 327678 580294 363250 580350
rect 363306 580294 363374 580350
rect 363430 580294 363498 580350
rect 363554 580294 363622 580350
rect 363678 580294 381250 580350
rect 381306 580294 381374 580350
rect 381430 580294 381498 580350
rect 381554 580294 381622 580350
rect 381678 580294 399250 580350
rect 399306 580294 399374 580350
rect 399430 580294 399498 580350
rect 399554 580294 399622 580350
rect 399678 580294 417250 580350
rect 417306 580294 417374 580350
rect 417430 580294 417498 580350
rect 417554 580294 417622 580350
rect 417678 580294 453250 580350
rect 453306 580294 453374 580350
rect 453430 580294 453498 580350
rect 453554 580294 453622 580350
rect 453678 580294 471250 580350
rect 471306 580294 471374 580350
rect 471430 580294 471498 580350
rect 471554 580294 471622 580350
rect 471678 580294 489250 580350
rect 489306 580294 489374 580350
rect 489430 580294 489498 580350
rect 489554 580294 489622 580350
rect 489678 580294 507250 580350
rect 507306 580294 507374 580350
rect 507430 580294 507498 580350
rect 507554 580294 507622 580350
rect 507678 580294 543250 580350
rect 543306 580294 543374 580350
rect 543430 580294 543498 580350
rect 543554 580294 543622 580350
rect 543678 580294 561250 580350
rect 561306 580294 561374 580350
rect 561430 580294 561498 580350
rect 561554 580294 561622 580350
rect 561678 580294 579250 580350
rect 579306 580294 579374 580350
rect 579430 580294 579498 580350
rect 579554 580294 579622 580350
rect 579678 580294 596496 580350
rect 596552 580294 596620 580350
rect 596676 580294 596744 580350
rect 596800 580294 596868 580350
rect 596924 580294 597980 580350
rect -1916 580226 597980 580294
rect -1916 580170 -860 580226
rect -804 580170 -736 580226
rect -680 580170 -612 580226
rect -556 580170 -488 580226
rect -432 580170 3250 580226
rect 3306 580170 3374 580226
rect 3430 580170 3498 580226
rect 3554 580170 3622 580226
rect 3678 580170 21250 580226
rect 21306 580170 21374 580226
rect 21430 580170 21498 580226
rect 21554 580170 21622 580226
rect 21678 580170 39250 580226
rect 39306 580170 39374 580226
rect 39430 580170 39498 580226
rect 39554 580170 39622 580226
rect 39678 580170 57250 580226
rect 57306 580170 57374 580226
rect 57430 580170 57498 580226
rect 57554 580170 57622 580226
rect 57678 580170 93250 580226
rect 93306 580170 93374 580226
rect 93430 580170 93498 580226
rect 93554 580170 93622 580226
rect 93678 580170 111250 580226
rect 111306 580170 111374 580226
rect 111430 580170 111498 580226
rect 111554 580170 111622 580226
rect 111678 580170 129250 580226
rect 129306 580170 129374 580226
rect 129430 580170 129498 580226
rect 129554 580170 129622 580226
rect 129678 580170 147250 580226
rect 147306 580170 147374 580226
rect 147430 580170 147498 580226
rect 147554 580170 147622 580226
rect 147678 580170 183250 580226
rect 183306 580170 183374 580226
rect 183430 580170 183498 580226
rect 183554 580170 183622 580226
rect 183678 580170 201250 580226
rect 201306 580170 201374 580226
rect 201430 580170 201498 580226
rect 201554 580170 201622 580226
rect 201678 580170 219250 580226
rect 219306 580170 219374 580226
rect 219430 580170 219498 580226
rect 219554 580170 219622 580226
rect 219678 580170 237250 580226
rect 237306 580170 237374 580226
rect 237430 580170 237498 580226
rect 237554 580170 237622 580226
rect 237678 580170 273250 580226
rect 273306 580170 273374 580226
rect 273430 580170 273498 580226
rect 273554 580170 273622 580226
rect 273678 580170 291250 580226
rect 291306 580170 291374 580226
rect 291430 580170 291498 580226
rect 291554 580170 291622 580226
rect 291678 580170 309250 580226
rect 309306 580170 309374 580226
rect 309430 580170 309498 580226
rect 309554 580170 309622 580226
rect 309678 580170 327250 580226
rect 327306 580170 327374 580226
rect 327430 580170 327498 580226
rect 327554 580170 327622 580226
rect 327678 580170 363250 580226
rect 363306 580170 363374 580226
rect 363430 580170 363498 580226
rect 363554 580170 363622 580226
rect 363678 580170 381250 580226
rect 381306 580170 381374 580226
rect 381430 580170 381498 580226
rect 381554 580170 381622 580226
rect 381678 580170 399250 580226
rect 399306 580170 399374 580226
rect 399430 580170 399498 580226
rect 399554 580170 399622 580226
rect 399678 580170 417250 580226
rect 417306 580170 417374 580226
rect 417430 580170 417498 580226
rect 417554 580170 417622 580226
rect 417678 580170 453250 580226
rect 453306 580170 453374 580226
rect 453430 580170 453498 580226
rect 453554 580170 453622 580226
rect 453678 580170 471250 580226
rect 471306 580170 471374 580226
rect 471430 580170 471498 580226
rect 471554 580170 471622 580226
rect 471678 580170 489250 580226
rect 489306 580170 489374 580226
rect 489430 580170 489498 580226
rect 489554 580170 489622 580226
rect 489678 580170 507250 580226
rect 507306 580170 507374 580226
rect 507430 580170 507498 580226
rect 507554 580170 507622 580226
rect 507678 580170 543250 580226
rect 543306 580170 543374 580226
rect 543430 580170 543498 580226
rect 543554 580170 543622 580226
rect 543678 580170 561250 580226
rect 561306 580170 561374 580226
rect 561430 580170 561498 580226
rect 561554 580170 561622 580226
rect 561678 580170 579250 580226
rect 579306 580170 579374 580226
rect 579430 580170 579498 580226
rect 579554 580170 579622 580226
rect 579678 580170 596496 580226
rect 596552 580170 596620 580226
rect 596676 580170 596744 580226
rect 596800 580170 596868 580226
rect 596924 580170 597980 580226
rect -1916 580102 597980 580170
rect -1916 580046 -860 580102
rect -804 580046 -736 580102
rect -680 580046 -612 580102
rect -556 580046 -488 580102
rect -432 580046 3250 580102
rect 3306 580046 3374 580102
rect 3430 580046 3498 580102
rect 3554 580046 3622 580102
rect 3678 580046 21250 580102
rect 21306 580046 21374 580102
rect 21430 580046 21498 580102
rect 21554 580046 21622 580102
rect 21678 580046 39250 580102
rect 39306 580046 39374 580102
rect 39430 580046 39498 580102
rect 39554 580046 39622 580102
rect 39678 580046 57250 580102
rect 57306 580046 57374 580102
rect 57430 580046 57498 580102
rect 57554 580046 57622 580102
rect 57678 580046 93250 580102
rect 93306 580046 93374 580102
rect 93430 580046 93498 580102
rect 93554 580046 93622 580102
rect 93678 580046 111250 580102
rect 111306 580046 111374 580102
rect 111430 580046 111498 580102
rect 111554 580046 111622 580102
rect 111678 580046 129250 580102
rect 129306 580046 129374 580102
rect 129430 580046 129498 580102
rect 129554 580046 129622 580102
rect 129678 580046 147250 580102
rect 147306 580046 147374 580102
rect 147430 580046 147498 580102
rect 147554 580046 147622 580102
rect 147678 580046 183250 580102
rect 183306 580046 183374 580102
rect 183430 580046 183498 580102
rect 183554 580046 183622 580102
rect 183678 580046 201250 580102
rect 201306 580046 201374 580102
rect 201430 580046 201498 580102
rect 201554 580046 201622 580102
rect 201678 580046 219250 580102
rect 219306 580046 219374 580102
rect 219430 580046 219498 580102
rect 219554 580046 219622 580102
rect 219678 580046 237250 580102
rect 237306 580046 237374 580102
rect 237430 580046 237498 580102
rect 237554 580046 237622 580102
rect 237678 580046 273250 580102
rect 273306 580046 273374 580102
rect 273430 580046 273498 580102
rect 273554 580046 273622 580102
rect 273678 580046 291250 580102
rect 291306 580046 291374 580102
rect 291430 580046 291498 580102
rect 291554 580046 291622 580102
rect 291678 580046 309250 580102
rect 309306 580046 309374 580102
rect 309430 580046 309498 580102
rect 309554 580046 309622 580102
rect 309678 580046 327250 580102
rect 327306 580046 327374 580102
rect 327430 580046 327498 580102
rect 327554 580046 327622 580102
rect 327678 580046 363250 580102
rect 363306 580046 363374 580102
rect 363430 580046 363498 580102
rect 363554 580046 363622 580102
rect 363678 580046 381250 580102
rect 381306 580046 381374 580102
rect 381430 580046 381498 580102
rect 381554 580046 381622 580102
rect 381678 580046 399250 580102
rect 399306 580046 399374 580102
rect 399430 580046 399498 580102
rect 399554 580046 399622 580102
rect 399678 580046 417250 580102
rect 417306 580046 417374 580102
rect 417430 580046 417498 580102
rect 417554 580046 417622 580102
rect 417678 580046 453250 580102
rect 453306 580046 453374 580102
rect 453430 580046 453498 580102
rect 453554 580046 453622 580102
rect 453678 580046 471250 580102
rect 471306 580046 471374 580102
rect 471430 580046 471498 580102
rect 471554 580046 471622 580102
rect 471678 580046 489250 580102
rect 489306 580046 489374 580102
rect 489430 580046 489498 580102
rect 489554 580046 489622 580102
rect 489678 580046 507250 580102
rect 507306 580046 507374 580102
rect 507430 580046 507498 580102
rect 507554 580046 507622 580102
rect 507678 580046 543250 580102
rect 543306 580046 543374 580102
rect 543430 580046 543498 580102
rect 543554 580046 543622 580102
rect 543678 580046 561250 580102
rect 561306 580046 561374 580102
rect 561430 580046 561498 580102
rect 561554 580046 561622 580102
rect 561678 580046 579250 580102
rect 579306 580046 579374 580102
rect 579430 580046 579498 580102
rect 579554 580046 579622 580102
rect 579678 580046 596496 580102
rect 596552 580046 596620 580102
rect 596676 580046 596744 580102
rect 596800 580046 596868 580102
rect 596924 580046 597980 580102
rect -1916 579978 597980 580046
rect -1916 579922 -860 579978
rect -804 579922 -736 579978
rect -680 579922 -612 579978
rect -556 579922 -488 579978
rect -432 579922 3250 579978
rect 3306 579922 3374 579978
rect 3430 579922 3498 579978
rect 3554 579922 3622 579978
rect 3678 579922 21250 579978
rect 21306 579922 21374 579978
rect 21430 579922 21498 579978
rect 21554 579922 21622 579978
rect 21678 579922 39250 579978
rect 39306 579922 39374 579978
rect 39430 579922 39498 579978
rect 39554 579922 39622 579978
rect 39678 579922 57250 579978
rect 57306 579922 57374 579978
rect 57430 579922 57498 579978
rect 57554 579922 57622 579978
rect 57678 579922 93250 579978
rect 93306 579922 93374 579978
rect 93430 579922 93498 579978
rect 93554 579922 93622 579978
rect 93678 579922 111250 579978
rect 111306 579922 111374 579978
rect 111430 579922 111498 579978
rect 111554 579922 111622 579978
rect 111678 579922 129250 579978
rect 129306 579922 129374 579978
rect 129430 579922 129498 579978
rect 129554 579922 129622 579978
rect 129678 579922 147250 579978
rect 147306 579922 147374 579978
rect 147430 579922 147498 579978
rect 147554 579922 147622 579978
rect 147678 579922 183250 579978
rect 183306 579922 183374 579978
rect 183430 579922 183498 579978
rect 183554 579922 183622 579978
rect 183678 579922 201250 579978
rect 201306 579922 201374 579978
rect 201430 579922 201498 579978
rect 201554 579922 201622 579978
rect 201678 579922 219250 579978
rect 219306 579922 219374 579978
rect 219430 579922 219498 579978
rect 219554 579922 219622 579978
rect 219678 579922 237250 579978
rect 237306 579922 237374 579978
rect 237430 579922 237498 579978
rect 237554 579922 237622 579978
rect 237678 579922 273250 579978
rect 273306 579922 273374 579978
rect 273430 579922 273498 579978
rect 273554 579922 273622 579978
rect 273678 579922 291250 579978
rect 291306 579922 291374 579978
rect 291430 579922 291498 579978
rect 291554 579922 291622 579978
rect 291678 579922 309250 579978
rect 309306 579922 309374 579978
rect 309430 579922 309498 579978
rect 309554 579922 309622 579978
rect 309678 579922 327250 579978
rect 327306 579922 327374 579978
rect 327430 579922 327498 579978
rect 327554 579922 327622 579978
rect 327678 579922 363250 579978
rect 363306 579922 363374 579978
rect 363430 579922 363498 579978
rect 363554 579922 363622 579978
rect 363678 579922 381250 579978
rect 381306 579922 381374 579978
rect 381430 579922 381498 579978
rect 381554 579922 381622 579978
rect 381678 579922 399250 579978
rect 399306 579922 399374 579978
rect 399430 579922 399498 579978
rect 399554 579922 399622 579978
rect 399678 579922 417250 579978
rect 417306 579922 417374 579978
rect 417430 579922 417498 579978
rect 417554 579922 417622 579978
rect 417678 579922 453250 579978
rect 453306 579922 453374 579978
rect 453430 579922 453498 579978
rect 453554 579922 453622 579978
rect 453678 579922 471250 579978
rect 471306 579922 471374 579978
rect 471430 579922 471498 579978
rect 471554 579922 471622 579978
rect 471678 579922 489250 579978
rect 489306 579922 489374 579978
rect 489430 579922 489498 579978
rect 489554 579922 489622 579978
rect 489678 579922 507250 579978
rect 507306 579922 507374 579978
rect 507430 579922 507498 579978
rect 507554 579922 507622 579978
rect 507678 579922 543250 579978
rect 543306 579922 543374 579978
rect 543430 579922 543498 579978
rect 543554 579922 543622 579978
rect 543678 579922 561250 579978
rect 561306 579922 561374 579978
rect 561430 579922 561498 579978
rect 561554 579922 561622 579978
rect 561678 579922 579250 579978
rect 579306 579922 579374 579978
rect 579430 579922 579498 579978
rect 579554 579922 579622 579978
rect 579678 579922 596496 579978
rect 596552 579922 596620 579978
rect 596676 579922 596744 579978
rect 596800 579922 596868 579978
rect 596924 579922 597980 579978
rect -1916 579826 597980 579922
rect -1916 568350 597980 568446
rect -1916 568294 -1820 568350
rect -1764 568294 -1696 568350
rect -1640 568294 -1572 568350
rect -1516 568294 -1448 568350
rect -1392 568294 6970 568350
rect 7026 568294 7094 568350
rect 7150 568294 7218 568350
rect 7274 568294 7342 568350
rect 7398 568294 24970 568350
rect 25026 568294 25094 568350
rect 25150 568294 25218 568350
rect 25274 568294 25342 568350
rect 25398 568294 42970 568350
rect 43026 568294 43094 568350
rect 43150 568294 43218 568350
rect 43274 568294 43342 568350
rect 43398 568294 60970 568350
rect 61026 568294 61094 568350
rect 61150 568294 61218 568350
rect 61274 568294 61342 568350
rect 61398 568294 78970 568350
rect 79026 568294 79094 568350
rect 79150 568294 79218 568350
rect 79274 568294 79342 568350
rect 79398 568294 96970 568350
rect 97026 568294 97094 568350
rect 97150 568294 97218 568350
rect 97274 568294 97342 568350
rect 97398 568294 132970 568350
rect 133026 568294 133094 568350
rect 133150 568294 133218 568350
rect 133274 568294 133342 568350
rect 133398 568294 150970 568350
rect 151026 568294 151094 568350
rect 151150 568294 151218 568350
rect 151274 568294 151342 568350
rect 151398 568294 168970 568350
rect 169026 568294 169094 568350
rect 169150 568294 169218 568350
rect 169274 568294 169342 568350
rect 169398 568294 186970 568350
rect 187026 568294 187094 568350
rect 187150 568294 187218 568350
rect 187274 568294 187342 568350
rect 187398 568294 222970 568350
rect 223026 568294 223094 568350
rect 223150 568294 223218 568350
rect 223274 568294 223342 568350
rect 223398 568294 240970 568350
rect 241026 568294 241094 568350
rect 241150 568294 241218 568350
rect 241274 568294 241342 568350
rect 241398 568294 258970 568350
rect 259026 568294 259094 568350
rect 259150 568294 259218 568350
rect 259274 568294 259342 568350
rect 259398 568294 276970 568350
rect 277026 568294 277094 568350
rect 277150 568294 277218 568350
rect 277274 568294 277342 568350
rect 277398 568294 312970 568350
rect 313026 568294 313094 568350
rect 313150 568294 313218 568350
rect 313274 568294 313342 568350
rect 313398 568294 330970 568350
rect 331026 568294 331094 568350
rect 331150 568294 331218 568350
rect 331274 568294 331342 568350
rect 331398 568294 348970 568350
rect 349026 568294 349094 568350
rect 349150 568294 349218 568350
rect 349274 568294 349342 568350
rect 349398 568294 366970 568350
rect 367026 568294 367094 568350
rect 367150 568294 367218 568350
rect 367274 568294 367342 568350
rect 367398 568294 402970 568350
rect 403026 568294 403094 568350
rect 403150 568294 403218 568350
rect 403274 568294 403342 568350
rect 403398 568294 420970 568350
rect 421026 568294 421094 568350
rect 421150 568294 421218 568350
rect 421274 568294 421342 568350
rect 421398 568294 438970 568350
rect 439026 568294 439094 568350
rect 439150 568294 439218 568350
rect 439274 568294 439342 568350
rect 439398 568294 456970 568350
rect 457026 568294 457094 568350
rect 457150 568294 457218 568350
rect 457274 568294 457342 568350
rect 457398 568294 492970 568350
rect 493026 568294 493094 568350
rect 493150 568294 493218 568350
rect 493274 568294 493342 568350
rect 493398 568294 510970 568350
rect 511026 568294 511094 568350
rect 511150 568294 511218 568350
rect 511274 568294 511342 568350
rect 511398 568294 528970 568350
rect 529026 568294 529094 568350
rect 529150 568294 529218 568350
rect 529274 568294 529342 568350
rect 529398 568294 546970 568350
rect 547026 568294 547094 568350
rect 547150 568294 547218 568350
rect 547274 568294 547342 568350
rect 547398 568294 564970 568350
rect 565026 568294 565094 568350
rect 565150 568294 565218 568350
rect 565274 568294 565342 568350
rect 565398 568294 582970 568350
rect 583026 568294 583094 568350
rect 583150 568294 583218 568350
rect 583274 568294 583342 568350
rect 583398 568294 597456 568350
rect 597512 568294 597580 568350
rect 597636 568294 597704 568350
rect 597760 568294 597828 568350
rect 597884 568294 597980 568350
rect -1916 568226 597980 568294
rect -1916 568170 -1820 568226
rect -1764 568170 -1696 568226
rect -1640 568170 -1572 568226
rect -1516 568170 -1448 568226
rect -1392 568170 6970 568226
rect 7026 568170 7094 568226
rect 7150 568170 7218 568226
rect 7274 568170 7342 568226
rect 7398 568170 24970 568226
rect 25026 568170 25094 568226
rect 25150 568170 25218 568226
rect 25274 568170 25342 568226
rect 25398 568170 42970 568226
rect 43026 568170 43094 568226
rect 43150 568170 43218 568226
rect 43274 568170 43342 568226
rect 43398 568170 60970 568226
rect 61026 568170 61094 568226
rect 61150 568170 61218 568226
rect 61274 568170 61342 568226
rect 61398 568170 78970 568226
rect 79026 568170 79094 568226
rect 79150 568170 79218 568226
rect 79274 568170 79342 568226
rect 79398 568170 96970 568226
rect 97026 568170 97094 568226
rect 97150 568170 97218 568226
rect 97274 568170 97342 568226
rect 97398 568170 132970 568226
rect 133026 568170 133094 568226
rect 133150 568170 133218 568226
rect 133274 568170 133342 568226
rect 133398 568170 150970 568226
rect 151026 568170 151094 568226
rect 151150 568170 151218 568226
rect 151274 568170 151342 568226
rect 151398 568170 168970 568226
rect 169026 568170 169094 568226
rect 169150 568170 169218 568226
rect 169274 568170 169342 568226
rect 169398 568170 186970 568226
rect 187026 568170 187094 568226
rect 187150 568170 187218 568226
rect 187274 568170 187342 568226
rect 187398 568170 222970 568226
rect 223026 568170 223094 568226
rect 223150 568170 223218 568226
rect 223274 568170 223342 568226
rect 223398 568170 240970 568226
rect 241026 568170 241094 568226
rect 241150 568170 241218 568226
rect 241274 568170 241342 568226
rect 241398 568170 258970 568226
rect 259026 568170 259094 568226
rect 259150 568170 259218 568226
rect 259274 568170 259342 568226
rect 259398 568170 276970 568226
rect 277026 568170 277094 568226
rect 277150 568170 277218 568226
rect 277274 568170 277342 568226
rect 277398 568170 312970 568226
rect 313026 568170 313094 568226
rect 313150 568170 313218 568226
rect 313274 568170 313342 568226
rect 313398 568170 330970 568226
rect 331026 568170 331094 568226
rect 331150 568170 331218 568226
rect 331274 568170 331342 568226
rect 331398 568170 348970 568226
rect 349026 568170 349094 568226
rect 349150 568170 349218 568226
rect 349274 568170 349342 568226
rect 349398 568170 366970 568226
rect 367026 568170 367094 568226
rect 367150 568170 367218 568226
rect 367274 568170 367342 568226
rect 367398 568170 402970 568226
rect 403026 568170 403094 568226
rect 403150 568170 403218 568226
rect 403274 568170 403342 568226
rect 403398 568170 420970 568226
rect 421026 568170 421094 568226
rect 421150 568170 421218 568226
rect 421274 568170 421342 568226
rect 421398 568170 438970 568226
rect 439026 568170 439094 568226
rect 439150 568170 439218 568226
rect 439274 568170 439342 568226
rect 439398 568170 456970 568226
rect 457026 568170 457094 568226
rect 457150 568170 457218 568226
rect 457274 568170 457342 568226
rect 457398 568170 492970 568226
rect 493026 568170 493094 568226
rect 493150 568170 493218 568226
rect 493274 568170 493342 568226
rect 493398 568170 510970 568226
rect 511026 568170 511094 568226
rect 511150 568170 511218 568226
rect 511274 568170 511342 568226
rect 511398 568170 528970 568226
rect 529026 568170 529094 568226
rect 529150 568170 529218 568226
rect 529274 568170 529342 568226
rect 529398 568170 546970 568226
rect 547026 568170 547094 568226
rect 547150 568170 547218 568226
rect 547274 568170 547342 568226
rect 547398 568170 564970 568226
rect 565026 568170 565094 568226
rect 565150 568170 565218 568226
rect 565274 568170 565342 568226
rect 565398 568170 582970 568226
rect 583026 568170 583094 568226
rect 583150 568170 583218 568226
rect 583274 568170 583342 568226
rect 583398 568170 597456 568226
rect 597512 568170 597580 568226
rect 597636 568170 597704 568226
rect 597760 568170 597828 568226
rect 597884 568170 597980 568226
rect -1916 568102 597980 568170
rect -1916 568046 -1820 568102
rect -1764 568046 -1696 568102
rect -1640 568046 -1572 568102
rect -1516 568046 -1448 568102
rect -1392 568046 6970 568102
rect 7026 568046 7094 568102
rect 7150 568046 7218 568102
rect 7274 568046 7342 568102
rect 7398 568046 24970 568102
rect 25026 568046 25094 568102
rect 25150 568046 25218 568102
rect 25274 568046 25342 568102
rect 25398 568046 42970 568102
rect 43026 568046 43094 568102
rect 43150 568046 43218 568102
rect 43274 568046 43342 568102
rect 43398 568046 60970 568102
rect 61026 568046 61094 568102
rect 61150 568046 61218 568102
rect 61274 568046 61342 568102
rect 61398 568046 78970 568102
rect 79026 568046 79094 568102
rect 79150 568046 79218 568102
rect 79274 568046 79342 568102
rect 79398 568046 96970 568102
rect 97026 568046 97094 568102
rect 97150 568046 97218 568102
rect 97274 568046 97342 568102
rect 97398 568046 132970 568102
rect 133026 568046 133094 568102
rect 133150 568046 133218 568102
rect 133274 568046 133342 568102
rect 133398 568046 150970 568102
rect 151026 568046 151094 568102
rect 151150 568046 151218 568102
rect 151274 568046 151342 568102
rect 151398 568046 168970 568102
rect 169026 568046 169094 568102
rect 169150 568046 169218 568102
rect 169274 568046 169342 568102
rect 169398 568046 186970 568102
rect 187026 568046 187094 568102
rect 187150 568046 187218 568102
rect 187274 568046 187342 568102
rect 187398 568046 222970 568102
rect 223026 568046 223094 568102
rect 223150 568046 223218 568102
rect 223274 568046 223342 568102
rect 223398 568046 240970 568102
rect 241026 568046 241094 568102
rect 241150 568046 241218 568102
rect 241274 568046 241342 568102
rect 241398 568046 258970 568102
rect 259026 568046 259094 568102
rect 259150 568046 259218 568102
rect 259274 568046 259342 568102
rect 259398 568046 276970 568102
rect 277026 568046 277094 568102
rect 277150 568046 277218 568102
rect 277274 568046 277342 568102
rect 277398 568046 312970 568102
rect 313026 568046 313094 568102
rect 313150 568046 313218 568102
rect 313274 568046 313342 568102
rect 313398 568046 330970 568102
rect 331026 568046 331094 568102
rect 331150 568046 331218 568102
rect 331274 568046 331342 568102
rect 331398 568046 348970 568102
rect 349026 568046 349094 568102
rect 349150 568046 349218 568102
rect 349274 568046 349342 568102
rect 349398 568046 366970 568102
rect 367026 568046 367094 568102
rect 367150 568046 367218 568102
rect 367274 568046 367342 568102
rect 367398 568046 402970 568102
rect 403026 568046 403094 568102
rect 403150 568046 403218 568102
rect 403274 568046 403342 568102
rect 403398 568046 420970 568102
rect 421026 568046 421094 568102
rect 421150 568046 421218 568102
rect 421274 568046 421342 568102
rect 421398 568046 438970 568102
rect 439026 568046 439094 568102
rect 439150 568046 439218 568102
rect 439274 568046 439342 568102
rect 439398 568046 456970 568102
rect 457026 568046 457094 568102
rect 457150 568046 457218 568102
rect 457274 568046 457342 568102
rect 457398 568046 492970 568102
rect 493026 568046 493094 568102
rect 493150 568046 493218 568102
rect 493274 568046 493342 568102
rect 493398 568046 510970 568102
rect 511026 568046 511094 568102
rect 511150 568046 511218 568102
rect 511274 568046 511342 568102
rect 511398 568046 528970 568102
rect 529026 568046 529094 568102
rect 529150 568046 529218 568102
rect 529274 568046 529342 568102
rect 529398 568046 546970 568102
rect 547026 568046 547094 568102
rect 547150 568046 547218 568102
rect 547274 568046 547342 568102
rect 547398 568046 564970 568102
rect 565026 568046 565094 568102
rect 565150 568046 565218 568102
rect 565274 568046 565342 568102
rect 565398 568046 582970 568102
rect 583026 568046 583094 568102
rect 583150 568046 583218 568102
rect 583274 568046 583342 568102
rect 583398 568046 597456 568102
rect 597512 568046 597580 568102
rect 597636 568046 597704 568102
rect 597760 568046 597828 568102
rect 597884 568046 597980 568102
rect -1916 567978 597980 568046
rect -1916 567922 -1820 567978
rect -1764 567922 -1696 567978
rect -1640 567922 -1572 567978
rect -1516 567922 -1448 567978
rect -1392 567922 6970 567978
rect 7026 567922 7094 567978
rect 7150 567922 7218 567978
rect 7274 567922 7342 567978
rect 7398 567922 24970 567978
rect 25026 567922 25094 567978
rect 25150 567922 25218 567978
rect 25274 567922 25342 567978
rect 25398 567922 42970 567978
rect 43026 567922 43094 567978
rect 43150 567922 43218 567978
rect 43274 567922 43342 567978
rect 43398 567922 60970 567978
rect 61026 567922 61094 567978
rect 61150 567922 61218 567978
rect 61274 567922 61342 567978
rect 61398 567922 78970 567978
rect 79026 567922 79094 567978
rect 79150 567922 79218 567978
rect 79274 567922 79342 567978
rect 79398 567922 96970 567978
rect 97026 567922 97094 567978
rect 97150 567922 97218 567978
rect 97274 567922 97342 567978
rect 97398 567922 132970 567978
rect 133026 567922 133094 567978
rect 133150 567922 133218 567978
rect 133274 567922 133342 567978
rect 133398 567922 150970 567978
rect 151026 567922 151094 567978
rect 151150 567922 151218 567978
rect 151274 567922 151342 567978
rect 151398 567922 168970 567978
rect 169026 567922 169094 567978
rect 169150 567922 169218 567978
rect 169274 567922 169342 567978
rect 169398 567922 186970 567978
rect 187026 567922 187094 567978
rect 187150 567922 187218 567978
rect 187274 567922 187342 567978
rect 187398 567922 222970 567978
rect 223026 567922 223094 567978
rect 223150 567922 223218 567978
rect 223274 567922 223342 567978
rect 223398 567922 240970 567978
rect 241026 567922 241094 567978
rect 241150 567922 241218 567978
rect 241274 567922 241342 567978
rect 241398 567922 258970 567978
rect 259026 567922 259094 567978
rect 259150 567922 259218 567978
rect 259274 567922 259342 567978
rect 259398 567922 276970 567978
rect 277026 567922 277094 567978
rect 277150 567922 277218 567978
rect 277274 567922 277342 567978
rect 277398 567922 312970 567978
rect 313026 567922 313094 567978
rect 313150 567922 313218 567978
rect 313274 567922 313342 567978
rect 313398 567922 330970 567978
rect 331026 567922 331094 567978
rect 331150 567922 331218 567978
rect 331274 567922 331342 567978
rect 331398 567922 348970 567978
rect 349026 567922 349094 567978
rect 349150 567922 349218 567978
rect 349274 567922 349342 567978
rect 349398 567922 366970 567978
rect 367026 567922 367094 567978
rect 367150 567922 367218 567978
rect 367274 567922 367342 567978
rect 367398 567922 402970 567978
rect 403026 567922 403094 567978
rect 403150 567922 403218 567978
rect 403274 567922 403342 567978
rect 403398 567922 420970 567978
rect 421026 567922 421094 567978
rect 421150 567922 421218 567978
rect 421274 567922 421342 567978
rect 421398 567922 438970 567978
rect 439026 567922 439094 567978
rect 439150 567922 439218 567978
rect 439274 567922 439342 567978
rect 439398 567922 456970 567978
rect 457026 567922 457094 567978
rect 457150 567922 457218 567978
rect 457274 567922 457342 567978
rect 457398 567922 492970 567978
rect 493026 567922 493094 567978
rect 493150 567922 493218 567978
rect 493274 567922 493342 567978
rect 493398 567922 510970 567978
rect 511026 567922 511094 567978
rect 511150 567922 511218 567978
rect 511274 567922 511342 567978
rect 511398 567922 528970 567978
rect 529026 567922 529094 567978
rect 529150 567922 529218 567978
rect 529274 567922 529342 567978
rect 529398 567922 546970 567978
rect 547026 567922 547094 567978
rect 547150 567922 547218 567978
rect 547274 567922 547342 567978
rect 547398 567922 564970 567978
rect 565026 567922 565094 567978
rect 565150 567922 565218 567978
rect 565274 567922 565342 567978
rect 565398 567922 582970 567978
rect 583026 567922 583094 567978
rect 583150 567922 583218 567978
rect 583274 567922 583342 567978
rect 583398 567922 597456 567978
rect 597512 567922 597580 567978
rect 597636 567922 597704 567978
rect 597760 567922 597828 567978
rect 597884 567922 597980 567978
rect -1916 567826 597980 567922
rect -1916 562350 597980 562446
rect -1916 562294 -860 562350
rect -804 562294 -736 562350
rect -680 562294 -612 562350
rect -556 562294 -488 562350
rect -432 562294 3250 562350
rect 3306 562294 3374 562350
rect 3430 562294 3498 562350
rect 3554 562294 3622 562350
rect 3678 562294 21250 562350
rect 21306 562294 21374 562350
rect 21430 562294 21498 562350
rect 21554 562294 21622 562350
rect 21678 562294 39250 562350
rect 39306 562294 39374 562350
rect 39430 562294 39498 562350
rect 39554 562294 39622 562350
rect 39678 562294 57250 562350
rect 57306 562294 57374 562350
rect 57430 562294 57498 562350
rect 57554 562294 57622 562350
rect 57678 562294 93250 562350
rect 93306 562294 93374 562350
rect 93430 562294 93498 562350
rect 93554 562294 93622 562350
rect 93678 562294 111250 562350
rect 111306 562294 111374 562350
rect 111430 562294 111498 562350
rect 111554 562294 111622 562350
rect 111678 562294 129250 562350
rect 129306 562294 129374 562350
rect 129430 562294 129498 562350
rect 129554 562294 129622 562350
rect 129678 562294 147250 562350
rect 147306 562294 147374 562350
rect 147430 562294 147498 562350
rect 147554 562294 147622 562350
rect 147678 562294 183250 562350
rect 183306 562294 183374 562350
rect 183430 562294 183498 562350
rect 183554 562294 183622 562350
rect 183678 562294 201250 562350
rect 201306 562294 201374 562350
rect 201430 562294 201498 562350
rect 201554 562294 201622 562350
rect 201678 562294 219250 562350
rect 219306 562294 219374 562350
rect 219430 562294 219498 562350
rect 219554 562294 219622 562350
rect 219678 562294 237250 562350
rect 237306 562294 237374 562350
rect 237430 562294 237498 562350
rect 237554 562294 237622 562350
rect 237678 562294 273250 562350
rect 273306 562294 273374 562350
rect 273430 562294 273498 562350
rect 273554 562294 273622 562350
rect 273678 562294 291250 562350
rect 291306 562294 291374 562350
rect 291430 562294 291498 562350
rect 291554 562294 291622 562350
rect 291678 562294 309250 562350
rect 309306 562294 309374 562350
rect 309430 562294 309498 562350
rect 309554 562294 309622 562350
rect 309678 562294 327250 562350
rect 327306 562294 327374 562350
rect 327430 562294 327498 562350
rect 327554 562294 327622 562350
rect 327678 562294 363250 562350
rect 363306 562294 363374 562350
rect 363430 562294 363498 562350
rect 363554 562294 363622 562350
rect 363678 562294 381250 562350
rect 381306 562294 381374 562350
rect 381430 562294 381498 562350
rect 381554 562294 381622 562350
rect 381678 562294 399250 562350
rect 399306 562294 399374 562350
rect 399430 562294 399498 562350
rect 399554 562294 399622 562350
rect 399678 562294 417250 562350
rect 417306 562294 417374 562350
rect 417430 562294 417498 562350
rect 417554 562294 417622 562350
rect 417678 562294 453250 562350
rect 453306 562294 453374 562350
rect 453430 562294 453498 562350
rect 453554 562294 453622 562350
rect 453678 562294 471250 562350
rect 471306 562294 471374 562350
rect 471430 562294 471498 562350
rect 471554 562294 471622 562350
rect 471678 562294 489250 562350
rect 489306 562294 489374 562350
rect 489430 562294 489498 562350
rect 489554 562294 489622 562350
rect 489678 562294 507250 562350
rect 507306 562294 507374 562350
rect 507430 562294 507498 562350
rect 507554 562294 507622 562350
rect 507678 562294 543250 562350
rect 543306 562294 543374 562350
rect 543430 562294 543498 562350
rect 543554 562294 543622 562350
rect 543678 562294 561250 562350
rect 561306 562294 561374 562350
rect 561430 562294 561498 562350
rect 561554 562294 561622 562350
rect 561678 562294 579250 562350
rect 579306 562294 579374 562350
rect 579430 562294 579498 562350
rect 579554 562294 579622 562350
rect 579678 562294 596496 562350
rect 596552 562294 596620 562350
rect 596676 562294 596744 562350
rect 596800 562294 596868 562350
rect 596924 562294 597980 562350
rect -1916 562226 597980 562294
rect -1916 562170 -860 562226
rect -804 562170 -736 562226
rect -680 562170 -612 562226
rect -556 562170 -488 562226
rect -432 562170 3250 562226
rect 3306 562170 3374 562226
rect 3430 562170 3498 562226
rect 3554 562170 3622 562226
rect 3678 562170 21250 562226
rect 21306 562170 21374 562226
rect 21430 562170 21498 562226
rect 21554 562170 21622 562226
rect 21678 562170 39250 562226
rect 39306 562170 39374 562226
rect 39430 562170 39498 562226
rect 39554 562170 39622 562226
rect 39678 562170 57250 562226
rect 57306 562170 57374 562226
rect 57430 562170 57498 562226
rect 57554 562170 57622 562226
rect 57678 562170 93250 562226
rect 93306 562170 93374 562226
rect 93430 562170 93498 562226
rect 93554 562170 93622 562226
rect 93678 562170 111250 562226
rect 111306 562170 111374 562226
rect 111430 562170 111498 562226
rect 111554 562170 111622 562226
rect 111678 562170 129250 562226
rect 129306 562170 129374 562226
rect 129430 562170 129498 562226
rect 129554 562170 129622 562226
rect 129678 562170 147250 562226
rect 147306 562170 147374 562226
rect 147430 562170 147498 562226
rect 147554 562170 147622 562226
rect 147678 562170 183250 562226
rect 183306 562170 183374 562226
rect 183430 562170 183498 562226
rect 183554 562170 183622 562226
rect 183678 562170 201250 562226
rect 201306 562170 201374 562226
rect 201430 562170 201498 562226
rect 201554 562170 201622 562226
rect 201678 562170 219250 562226
rect 219306 562170 219374 562226
rect 219430 562170 219498 562226
rect 219554 562170 219622 562226
rect 219678 562170 237250 562226
rect 237306 562170 237374 562226
rect 237430 562170 237498 562226
rect 237554 562170 237622 562226
rect 237678 562170 273250 562226
rect 273306 562170 273374 562226
rect 273430 562170 273498 562226
rect 273554 562170 273622 562226
rect 273678 562170 291250 562226
rect 291306 562170 291374 562226
rect 291430 562170 291498 562226
rect 291554 562170 291622 562226
rect 291678 562170 309250 562226
rect 309306 562170 309374 562226
rect 309430 562170 309498 562226
rect 309554 562170 309622 562226
rect 309678 562170 327250 562226
rect 327306 562170 327374 562226
rect 327430 562170 327498 562226
rect 327554 562170 327622 562226
rect 327678 562170 363250 562226
rect 363306 562170 363374 562226
rect 363430 562170 363498 562226
rect 363554 562170 363622 562226
rect 363678 562170 381250 562226
rect 381306 562170 381374 562226
rect 381430 562170 381498 562226
rect 381554 562170 381622 562226
rect 381678 562170 399250 562226
rect 399306 562170 399374 562226
rect 399430 562170 399498 562226
rect 399554 562170 399622 562226
rect 399678 562170 417250 562226
rect 417306 562170 417374 562226
rect 417430 562170 417498 562226
rect 417554 562170 417622 562226
rect 417678 562170 453250 562226
rect 453306 562170 453374 562226
rect 453430 562170 453498 562226
rect 453554 562170 453622 562226
rect 453678 562170 471250 562226
rect 471306 562170 471374 562226
rect 471430 562170 471498 562226
rect 471554 562170 471622 562226
rect 471678 562170 489250 562226
rect 489306 562170 489374 562226
rect 489430 562170 489498 562226
rect 489554 562170 489622 562226
rect 489678 562170 507250 562226
rect 507306 562170 507374 562226
rect 507430 562170 507498 562226
rect 507554 562170 507622 562226
rect 507678 562170 543250 562226
rect 543306 562170 543374 562226
rect 543430 562170 543498 562226
rect 543554 562170 543622 562226
rect 543678 562170 561250 562226
rect 561306 562170 561374 562226
rect 561430 562170 561498 562226
rect 561554 562170 561622 562226
rect 561678 562170 579250 562226
rect 579306 562170 579374 562226
rect 579430 562170 579498 562226
rect 579554 562170 579622 562226
rect 579678 562170 596496 562226
rect 596552 562170 596620 562226
rect 596676 562170 596744 562226
rect 596800 562170 596868 562226
rect 596924 562170 597980 562226
rect -1916 562102 597980 562170
rect -1916 562046 -860 562102
rect -804 562046 -736 562102
rect -680 562046 -612 562102
rect -556 562046 -488 562102
rect -432 562046 3250 562102
rect 3306 562046 3374 562102
rect 3430 562046 3498 562102
rect 3554 562046 3622 562102
rect 3678 562046 21250 562102
rect 21306 562046 21374 562102
rect 21430 562046 21498 562102
rect 21554 562046 21622 562102
rect 21678 562046 39250 562102
rect 39306 562046 39374 562102
rect 39430 562046 39498 562102
rect 39554 562046 39622 562102
rect 39678 562046 57250 562102
rect 57306 562046 57374 562102
rect 57430 562046 57498 562102
rect 57554 562046 57622 562102
rect 57678 562046 93250 562102
rect 93306 562046 93374 562102
rect 93430 562046 93498 562102
rect 93554 562046 93622 562102
rect 93678 562046 111250 562102
rect 111306 562046 111374 562102
rect 111430 562046 111498 562102
rect 111554 562046 111622 562102
rect 111678 562046 129250 562102
rect 129306 562046 129374 562102
rect 129430 562046 129498 562102
rect 129554 562046 129622 562102
rect 129678 562046 147250 562102
rect 147306 562046 147374 562102
rect 147430 562046 147498 562102
rect 147554 562046 147622 562102
rect 147678 562046 183250 562102
rect 183306 562046 183374 562102
rect 183430 562046 183498 562102
rect 183554 562046 183622 562102
rect 183678 562046 201250 562102
rect 201306 562046 201374 562102
rect 201430 562046 201498 562102
rect 201554 562046 201622 562102
rect 201678 562046 219250 562102
rect 219306 562046 219374 562102
rect 219430 562046 219498 562102
rect 219554 562046 219622 562102
rect 219678 562046 237250 562102
rect 237306 562046 237374 562102
rect 237430 562046 237498 562102
rect 237554 562046 237622 562102
rect 237678 562046 273250 562102
rect 273306 562046 273374 562102
rect 273430 562046 273498 562102
rect 273554 562046 273622 562102
rect 273678 562046 291250 562102
rect 291306 562046 291374 562102
rect 291430 562046 291498 562102
rect 291554 562046 291622 562102
rect 291678 562046 309250 562102
rect 309306 562046 309374 562102
rect 309430 562046 309498 562102
rect 309554 562046 309622 562102
rect 309678 562046 327250 562102
rect 327306 562046 327374 562102
rect 327430 562046 327498 562102
rect 327554 562046 327622 562102
rect 327678 562046 363250 562102
rect 363306 562046 363374 562102
rect 363430 562046 363498 562102
rect 363554 562046 363622 562102
rect 363678 562046 381250 562102
rect 381306 562046 381374 562102
rect 381430 562046 381498 562102
rect 381554 562046 381622 562102
rect 381678 562046 399250 562102
rect 399306 562046 399374 562102
rect 399430 562046 399498 562102
rect 399554 562046 399622 562102
rect 399678 562046 417250 562102
rect 417306 562046 417374 562102
rect 417430 562046 417498 562102
rect 417554 562046 417622 562102
rect 417678 562046 453250 562102
rect 453306 562046 453374 562102
rect 453430 562046 453498 562102
rect 453554 562046 453622 562102
rect 453678 562046 471250 562102
rect 471306 562046 471374 562102
rect 471430 562046 471498 562102
rect 471554 562046 471622 562102
rect 471678 562046 489250 562102
rect 489306 562046 489374 562102
rect 489430 562046 489498 562102
rect 489554 562046 489622 562102
rect 489678 562046 507250 562102
rect 507306 562046 507374 562102
rect 507430 562046 507498 562102
rect 507554 562046 507622 562102
rect 507678 562046 543250 562102
rect 543306 562046 543374 562102
rect 543430 562046 543498 562102
rect 543554 562046 543622 562102
rect 543678 562046 561250 562102
rect 561306 562046 561374 562102
rect 561430 562046 561498 562102
rect 561554 562046 561622 562102
rect 561678 562046 579250 562102
rect 579306 562046 579374 562102
rect 579430 562046 579498 562102
rect 579554 562046 579622 562102
rect 579678 562046 596496 562102
rect 596552 562046 596620 562102
rect 596676 562046 596744 562102
rect 596800 562046 596868 562102
rect 596924 562046 597980 562102
rect -1916 561978 597980 562046
rect -1916 561922 -860 561978
rect -804 561922 -736 561978
rect -680 561922 -612 561978
rect -556 561922 -488 561978
rect -432 561922 3250 561978
rect 3306 561922 3374 561978
rect 3430 561922 3498 561978
rect 3554 561922 3622 561978
rect 3678 561922 21250 561978
rect 21306 561922 21374 561978
rect 21430 561922 21498 561978
rect 21554 561922 21622 561978
rect 21678 561922 39250 561978
rect 39306 561922 39374 561978
rect 39430 561922 39498 561978
rect 39554 561922 39622 561978
rect 39678 561922 57250 561978
rect 57306 561922 57374 561978
rect 57430 561922 57498 561978
rect 57554 561922 57622 561978
rect 57678 561922 93250 561978
rect 93306 561922 93374 561978
rect 93430 561922 93498 561978
rect 93554 561922 93622 561978
rect 93678 561922 111250 561978
rect 111306 561922 111374 561978
rect 111430 561922 111498 561978
rect 111554 561922 111622 561978
rect 111678 561922 129250 561978
rect 129306 561922 129374 561978
rect 129430 561922 129498 561978
rect 129554 561922 129622 561978
rect 129678 561922 147250 561978
rect 147306 561922 147374 561978
rect 147430 561922 147498 561978
rect 147554 561922 147622 561978
rect 147678 561922 183250 561978
rect 183306 561922 183374 561978
rect 183430 561922 183498 561978
rect 183554 561922 183622 561978
rect 183678 561922 201250 561978
rect 201306 561922 201374 561978
rect 201430 561922 201498 561978
rect 201554 561922 201622 561978
rect 201678 561922 219250 561978
rect 219306 561922 219374 561978
rect 219430 561922 219498 561978
rect 219554 561922 219622 561978
rect 219678 561922 237250 561978
rect 237306 561922 237374 561978
rect 237430 561922 237498 561978
rect 237554 561922 237622 561978
rect 237678 561922 273250 561978
rect 273306 561922 273374 561978
rect 273430 561922 273498 561978
rect 273554 561922 273622 561978
rect 273678 561922 291250 561978
rect 291306 561922 291374 561978
rect 291430 561922 291498 561978
rect 291554 561922 291622 561978
rect 291678 561922 309250 561978
rect 309306 561922 309374 561978
rect 309430 561922 309498 561978
rect 309554 561922 309622 561978
rect 309678 561922 327250 561978
rect 327306 561922 327374 561978
rect 327430 561922 327498 561978
rect 327554 561922 327622 561978
rect 327678 561922 363250 561978
rect 363306 561922 363374 561978
rect 363430 561922 363498 561978
rect 363554 561922 363622 561978
rect 363678 561922 381250 561978
rect 381306 561922 381374 561978
rect 381430 561922 381498 561978
rect 381554 561922 381622 561978
rect 381678 561922 399250 561978
rect 399306 561922 399374 561978
rect 399430 561922 399498 561978
rect 399554 561922 399622 561978
rect 399678 561922 417250 561978
rect 417306 561922 417374 561978
rect 417430 561922 417498 561978
rect 417554 561922 417622 561978
rect 417678 561922 453250 561978
rect 453306 561922 453374 561978
rect 453430 561922 453498 561978
rect 453554 561922 453622 561978
rect 453678 561922 471250 561978
rect 471306 561922 471374 561978
rect 471430 561922 471498 561978
rect 471554 561922 471622 561978
rect 471678 561922 489250 561978
rect 489306 561922 489374 561978
rect 489430 561922 489498 561978
rect 489554 561922 489622 561978
rect 489678 561922 507250 561978
rect 507306 561922 507374 561978
rect 507430 561922 507498 561978
rect 507554 561922 507622 561978
rect 507678 561922 543250 561978
rect 543306 561922 543374 561978
rect 543430 561922 543498 561978
rect 543554 561922 543622 561978
rect 543678 561922 561250 561978
rect 561306 561922 561374 561978
rect 561430 561922 561498 561978
rect 561554 561922 561622 561978
rect 561678 561922 579250 561978
rect 579306 561922 579374 561978
rect 579430 561922 579498 561978
rect 579554 561922 579622 561978
rect 579678 561922 596496 561978
rect 596552 561922 596620 561978
rect 596676 561922 596744 561978
rect 596800 561922 596868 561978
rect 596924 561922 597980 561978
rect -1916 561826 597980 561922
rect -1916 550350 597980 550446
rect -1916 550294 -1820 550350
rect -1764 550294 -1696 550350
rect -1640 550294 -1572 550350
rect -1516 550294 -1448 550350
rect -1392 550294 6970 550350
rect 7026 550294 7094 550350
rect 7150 550294 7218 550350
rect 7274 550294 7342 550350
rect 7398 550294 24970 550350
rect 25026 550294 25094 550350
rect 25150 550294 25218 550350
rect 25274 550294 25342 550350
rect 25398 550294 42970 550350
rect 43026 550294 43094 550350
rect 43150 550294 43218 550350
rect 43274 550294 43342 550350
rect 43398 550294 60970 550350
rect 61026 550294 61094 550350
rect 61150 550294 61218 550350
rect 61274 550294 61342 550350
rect 61398 550294 78970 550350
rect 79026 550294 79094 550350
rect 79150 550294 79218 550350
rect 79274 550294 79342 550350
rect 79398 550294 96970 550350
rect 97026 550294 97094 550350
rect 97150 550294 97218 550350
rect 97274 550294 97342 550350
rect 97398 550294 132970 550350
rect 133026 550294 133094 550350
rect 133150 550294 133218 550350
rect 133274 550294 133342 550350
rect 133398 550294 150970 550350
rect 151026 550294 151094 550350
rect 151150 550294 151218 550350
rect 151274 550294 151342 550350
rect 151398 550294 168970 550350
rect 169026 550294 169094 550350
rect 169150 550294 169218 550350
rect 169274 550294 169342 550350
rect 169398 550294 186970 550350
rect 187026 550294 187094 550350
rect 187150 550294 187218 550350
rect 187274 550294 187342 550350
rect 187398 550294 222970 550350
rect 223026 550294 223094 550350
rect 223150 550294 223218 550350
rect 223274 550294 223342 550350
rect 223398 550294 240970 550350
rect 241026 550294 241094 550350
rect 241150 550294 241218 550350
rect 241274 550294 241342 550350
rect 241398 550294 258970 550350
rect 259026 550294 259094 550350
rect 259150 550294 259218 550350
rect 259274 550294 259342 550350
rect 259398 550294 276970 550350
rect 277026 550294 277094 550350
rect 277150 550294 277218 550350
rect 277274 550294 277342 550350
rect 277398 550294 312970 550350
rect 313026 550294 313094 550350
rect 313150 550294 313218 550350
rect 313274 550294 313342 550350
rect 313398 550294 330970 550350
rect 331026 550294 331094 550350
rect 331150 550294 331218 550350
rect 331274 550294 331342 550350
rect 331398 550294 348970 550350
rect 349026 550294 349094 550350
rect 349150 550294 349218 550350
rect 349274 550294 349342 550350
rect 349398 550294 366970 550350
rect 367026 550294 367094 550350
rect 367150 550294 367218 550350
rect 367274 550294 367342 550350
rect 367398 550294 402970 550350
rect 403026 550294 403094 550350
rect 403150 550294 403218 550350
rect 403274 550294 403342 550350
rect 403398 550294 420970 550350
rect 421026 550294 421094 550350
rect 421150 550294 421218 550350
rect 421274 550294 421342 550350
rect 421398 550294 438970 550350
rect 439026 550294 439094 550350
rect 439150 550294 439218 550350
rect 439274 550294 439342 550350
rect 439398 550294 456970 550350
rect 457026 550294 457094 550350
rect 457150 550294 457218 550350
rect 457274 550294 457342 550350
rect 457398 550294 492970 550350
rect 493026 550294 493094 550350
rect 493150 550294 493218 550350
rect 493274 550294 493342 550350
rect 493398 550294 510970 550350
rect 511026 550294 511094 550350
rect 511150 550294 511218 550350
rect 511274 550294 511342 550350
rect 511398 550294 528970 550350
rect 529026 550294 529094 550350
rect 529150 550294 529218 550350
rect 529274 550294 529342 550350
rect 529398 550294 546970 550350
rect 547026 550294 547094 550350
rect 547150 550294 547218 550350
rect 547274 550294 547342 550350
rect 547398 550294 564970 550350
rect 565026 550294 565094 550350
rect 565150 550294 565218 550350
rect 565274 550294 565342 550350
rect 565398 550294 582970 550350
rect 583026 550294 583094 550350
rect 583150 550294 583218 550350
rect 583274 550294 583342 550350
rect 583398 550294 597456 550350
rect 597512 550294 597580 550350
rect 597636 550294 597704 550350
rect 597760 550294 597828 550350
rect 597884 550294 597980 550350
rect -1916 550226 597980 550294
rect -1916 550170 -1820 550226
rect -1764 550170 -1696 550226
rect -1640 550170 -1572 550226
rect -1516 550170 -1448 550226
rect -1392 550170 6970 550226
rect 7026 550170 7094 550226
rect 7150 550170 7218 550226
rect 7274 550170 7342 550226
rect 7398 550170 24970 550226
rect 25026 550170 25094 550226
rect 25150 550170 25218 550226
rect 25274 550170 25342 550226
rect 25398 550170 42970 550226
rect 43026 550170 43094 550226
rect 43150 550170 43218 550226
rect 43274 550170 43342 550226
rect 43398 550170 60970 550226
rect 61026 550170 61094 550226
rect 61150 550170 61218 550226
rect 61274 550170 61342 550226
rect 61398 550170 78970 550226
rect 79026 550170 79094 550226
rect 79150 550170 79218 550226
rect 79274 550170 79342 550226
rect 79398 550170 96970 550226
rect 97026 550170 97094 550226
rect 97150 550170 97218 550226
rect 97274 550170 97342 550226
rect 97398 550170 132970 550226
rect 133026 550170 133094 550226
rect 133150 550170 133218 550226
rect 133274 550170 133342 550226
rect 133398 550170 150970 550226
rect 151026 550170 151094 550226
rect 151150 550170 151218 550226
rect 151274 550170 151342 550226
rect 151398 550170 168970 550226
rect 169026 550170 169094 550226
rect 169150 550170 169218 550226
rect 169274 550170 169342 550226
rect 169398 550170 186970 550226
rect 187026 550170 187094 550226
rect 187150 550170 187218 550226
rect 187274 550170 187342 550226
rect 187398 550170 222970 550226
rect 223026 550170 223094 550226
rect 223150 550170 223218 550226
rect 223274 550170 223342 550226
rect 223398 550170 240970 550226
rect 241026 550170 241094 550226
rect 241150 550170 241218 550226
rect 241274 550170 241342 550226
rect 241398 550170 258970 550226
rect 259026 550170 259094 550226
rect 259150 550170 259218 550226
rect 259274 550170 259342 550226
rect 259398 550170 276970 550226
rect 277026 550170 277094 550226
rect 277150 550170 277218 550226
rect 277274 550170 277342 550226
rect 277398 550170 312970 550226
rect 313026 550170 313094 550226
rect 313150 550170 313218 550226
rect 313274 550170 313342 550226
rect 313398 550170 330970 550226
rect 331026 550170 331094 550226
rect 331150 550170 331218 550226
rect 331274 550170 331342 550226
rect 331398 550170 348970 550226
rect 349026 550170 349094 550226
rect 349150 550170 349218 550226
rect 349274 550170 349342 550226
rect 349398 550170 366970 550226
rect 367026 550170 367094 550226
rect 367150 550170 367218 550226
rect 367274 550170 367342 550226
rect 367398 550170 402970 550226
rect 403026 550170 403094 550226
rect 403150 550170 403218 550226
rect 403274 550170 403342 550226
rect 403398 550170 420970 550226
rect 421026 550170 421094 550226
rect 421150 550170 421218 550226
rect 421274 550170 421342 550226
rect 421398 550170 438970 550226
rect 439026 550170 439094 550226
rect 439150 550170 439218 550226
rect 439274 550170 439342 550226
rect 439398 550170 456970 550226
rect 457026 550170 457094 550226
rect 457150 550170 457218 550226
rect 457274 550170 457342 550226
rect 457398 550170 492970 550226
rect 493026 550170 493094 550226
rect 493150 550170 493218 550226
rect 493274 550170 493342 550226
rect 493398 550170 510970 550226
rect 511026 550170 511094 550226
rect 511150 550170 511218 550226
rect 511274 550170 511342 550226
rect 511398 550170 528970 550226
rect 529026 550170 529094 550226
rect 529150 550170 529218 550226
rect 529274 550170 529342 550226
rect 529398 550170 546970 550226
rect 547026 550170 547094 550226
rect 547150 550170 547218 550226
rect 547274 550170 547342 550226
rect 547398 550170 564970 550226
rect 565026 550170 565094 550226
rect 565150 550170 565218 550226
rect 565274 550170 565342 550226
rect 565398 550170 582970 550226
rect 583026 550170 583094 550226
rect 583150 550170 583218 550226
rect 583274 550170 583342 550226
rect 583398 550170 597456 550226
rect 597512 550170 597580 550226
rect 597636 550170 597704 550226
rect 597760 550170 597828 550226
rect 597884 550170 597980 550226
rect -1916 550102 597980 550170
rect -1916 550046 -1820 550102
rect -1764 550046 -1696 550102
rect -1640 550046 -1572 550102
rect -1516 550046 -1448 550102
rect -1392 550046 6970 550102
rect 7026 550046 7094 550102
rect 7150 550046 7218 550102
rect 7274 550046 7342 550102
rect 7398 550046 24970 550102
rect 25026 550046 25094 550102
rect 25150 550046 25218 550102
rect 25274 550046 25342 550102
rect 25398 550046 42970 550102
rect 43026 550046 43094 550102
rect 43150 550046 43218 550102
rect 43274 550046 43342 550102
rect 43398 550046 60970 550102
rect 61026 550046 61094 550102
rect 61150 550046 61218 550102
rect 61274 550046 61342 550102
rect 61398 550046 78970 550102
rect 79026 550046 79094 550102
rect 79150 550046 79218 550102
rect 79274 550046 79342 550102
rect 79398 550046 96970 550102
rect 97026 550046 97094 550102
rect 97150 550046 97218 550102
rect 97274 550046 97342 550102
rect 97398 550046 132970 550102
rect 133026 550046 133094 550102
rect 133150 550046 133218 550102
rect 133274 550046 133342 550102
rect 133398 550046 150970 550102
rect 151026 550046 151094 550102
rect 151150 550046 151218 550102
rect 151274 550046 151342 550102
rect 151398 550046 168970 550102
rect 169026 550046 169094 550102
rect 169150 550046 169218 550102
rect 169274 550046 169342 550102
rect 169398 550046 186970 550102
rect 187026 550046 187094 550102
rect 187150 550046 187218 550102
rect 187274 550046 187342 550102
rect 187398 550046 222970 550102
rect 223026 550046 223094 550102
rect 223150 550046 223218 550102
rect 223274 550046 223342 550102
rect 223398 550046 240970 550102
rect 241026 550046 241094 550102
rect 241150 550046 241218 550102
rect 241274 550046 241342 550102
rect 241398 550046 258970 550102
rect 259026 550046 259094 550102
rect 259150 550046 259218 550102
rect 259274 550046 259342 550102
rect 259398 550046 276970 550102
rect 277026 550046 277094 550102
rect 277150 550046 277218 550102
rect 277274 550046 277342 550102
rect 277398 550046 312970 550102
rect 313026 550046 313094 550102
rect 313150 550046 313218 550102
rect 313274 550046 313342 550102
rect 313398 550046 330970 550102
rect 331026 550046 331094 550102
rect 331150 550046 331218 550102
rect 331274 550046 331342 550102
rect 331398 550046 348970 550102
rect 349026 550046 349094 550102
rect 349150 550046 349218 550102
rect 349274 550046 349342 550102
rect 349398 550046 366970 550102
rect 367026 550046 367094 550102
rect 367150 550046 367218 550102
rect 367274 550046 367342 550102
rect 367398 550046 402970 550102
rect 403026 550046 403094 550102
rect 403150 550046 403218 550102
rect 403274 550046 403342 550102
rect 403398 550046 420970 550102
rect 421026 550046 421094 550102
rect 421150 550046 421218 550102
rect 421274 550046 421342 550102
rect 421398 550046 438970 550102
rect 439026 550046 439094 550102
rect 439150 550046 439218 550102
rect 439274 550046 439342 550102
rect 439398 550046 456970 550102
rect 457026 550046 457094 550102
rect 457150 550046 457218 550102
rect 457274 550046 457342 550102
rect 457398 550046 492970 550102
rect 493026 550046 493094 550102
rect 493150 550046 493218 550102
rect 493274 550046 493342 550102
rect 493398 550046 510970 550102
rect 511026 550046 511094 550102
rect 511150 550046 511218 550102
rect 511274 550046 511342 550102
rect 511398 550046 528970 550102
rect 529026 550046 529094 550102
rect 529150 550046 529218 550102
rect 529274 550046 529342 550102
rect 529398 550046 546970 550102
rect 547026 550046 547094 550102
rect 547150 550046 547218 550102
rect 547274 550046 547342 550102
rect 547398 550046 564970 550102
rect 565026 550046 565094 550102
rect 565150 550046 565218 550102
rect 565274 550046 565342 550102
rect 565398 550046 582970 550102
rect 583026 550046 583094 550102
rect 583150 550046 583218 550102
rect 583274 550046 583342 550102
rect 583398 550046 597456 550102
rect 597512 550046 597580 550102
rect 597636 550046 597704 550102
rect 597760 550046 597828 550102
rect 597884 550046 597980 550102
rect -1916 549978 597980 550046
rect -1916 549922 -1820 549978
rect -1764 549922 -1696 549978
rect -1640 549922 -1572 549978
rect -1516 549922 -1448 549978
rect -1392 549922 6970 549978
rect 7026 549922 7094 549978
rect 7150 549922 7218 549978
rect 7274 549922 7342 549978
rect 7398 549922 24970 549978
rect 25026 549922 25094 549978
rect 25150 549922 25218 549978
rect 25274 549922 25342 549978
rect 25398 549922 42970 549978
rect 43026 549922 43094 549978
rect 43150 549922 43218 549978
rect 43274 549922 43342 549978
rect 43398 549922 60970 549978
rect 61026 549922 61094 549978
rect 61150 549922 61218 549978
rect 61274 549922 61342 549978
rect 61398 549922 78970 549978
rect 79026 549922 79094 549978
rect 79150 549922 79218 549978
rect 79274 549922 79342 549978
rect 79398 549922 96970 549978
rect 97026 549922 97094 549978
rect 97150 549922 97218 549978
rect 97274 549922 97342 549978
rect 97398 549922 132970 549978
rect 133026 549922 133094 549978
rect 133150 549922 133218 549978
rect 133274 549922 133342 549978
rect 133398 549922 150970 549978
rect 151026 549922 151094 549978
rect 151150 549922 151218 549978
rect 151274 549922 151342 549978
rect 151398 549922 168970 549978
rect 169026 549922 169094 549978
rect 169150 549922 169218 549978
rect 169274 549922 169342 549978
rect 169398 549922 186970 549978
rect 187026 549922 187094 549978
rect 187150 549922 187218 549978
rect 187274 549922 187342 549978
rect 187398 549922 222970 549978
rect 223026 549922 223094 549978
rect 223150 549922 223218 549978
rect 223274 549922 223342 549978
rect 223398 549922 240970 549978
rect 241026 549922 241094 549978
rect 241150 549922 241218 549978
rect 241274 549922 241342 549978
rect 241398 549922 258970 549978
rect 259026 549922 259094 549978
rect 259150 549922 259218 549978
rect 259274 549922 259342 549978
rect 259398 549922 276970 549978
rect 277026 549922 277094 549978
rect 277150 549922 277218 549978
rect 277274 549922 277342 549978
rect 277398 549922 312970 549978
rect 313026 549922 313094 549978
rect 313150 549922 313218 549978
rect 313274 549922 313342 549978
rect 313398 549922 330970 549978
rect 331026 549922 331094 549978
rect 331150 549922 331218 549978
rect 331274 549922 331342 549978
rect 331398 549922 348970 549978
rect 349026 549922 349094 549978
rect 349150 549922 349218 549978
rect 349274 549922 349342 549978
rect 349398 549922 366970 549978
rect 367026 549922 367094 549978
rect 367150 549922 367218 549978
rect 367274 549922 367342 549978
rect 367398 549922 402970 549978
rect 403026 549922 403094 549978
rect 403150 549922 403218 549978
rect 403274 549922 403342 549978
rect 403398 549922 420970 549978
rect 421026 549922 421094 549978
rect 421150 549922 421218 549978
rect 421274 549922 421342 549978
rect 421398 549922 438970 549978
rect 439026 549922 439094 549978
rect 439150 549922 439218 549978
rect 439274 549922 439342 549978
rect 439398 549922 456970 549978
rect 457026 549922 457094 549978
rect 457150 549922 457218 549978
rect 457274 549922 457342 549978
rect 457398 549922 492970 549978
rect 493026 549922 493094 549978
rect 493150 549922 493218 549978
rect 493274 549922 493342 549978
rect 493398 549922 510970 549978
rect 511026 549922 511094 549978
rect 511150 549922 511218 549978
rect 511274 549922 511342 549978
rect 511398 549922 528970 549978
rect 529026 549922 529094 549978
rect 529150 549922 529218 549978
rect 529274 549922 529342 549978
rect 529398 549922 546970 549978
rect 547026 549922 547094 549978
rect 547150 549922 547218 549978
rect 547274 549922 547342 549978
rect 547398 549922 564970 549978
rect 565026 549922 565094 549978
rect 565150 549922 565218 549978
rect 565274 549922 565342 549978
rect 565398 549922 582970 549978
rect 583026 549922 583094 549978
rect 583150 549922 583218 549978
rect 583274 549922 583342 549978
rect 583398 549922 597456 549978
rect 597512 549922 597580 549978
rect 597636 549922 597704 549978
rect 597760 549922 597828 549978
rect 597884 549922 597980 549978
rect -1916 549826 597980 549922
rect -1916 544350 597980 544446
rect -1916 544294 -860 544350
rect -804 544294 -736 544350
rect -680 544294 -612 544350
rect -556 544294 -488 544350
rect -432 544294 3250 544350
rect 3306 544294 3374 544350
rect 3430 544294 3498 544350
rect 3554 544294 3622 544350
rect 3678 544294 21250 544350
rect 21306 544294 21374 544350
rect 21430 544294 21498 544350
rect 21554 544294 21622 544350
rect 21678 544294 39250 544350
rect 39306 544294 39374 544350
rect 39430 544294 39498 544350
rect 39554 544294 39622 544350
rect 39678 544294 57250 544350
rect 57306 544294 57374 544350
rect 57430 544294 57498 544350
rect 57554 544294 57622 544350
rect 57678 544294 93250 544350
rect 93306 544294 93374 544350
rect 93430 544294 93498 544350
rect 93554 544294 93622 544350
rect 93678 544294 111250 544350
rect 111306 544294 111374 544350
rect 111430 544294 111498 544350
rect 111554 544294 111622 544350
rect 111678 544294 129250 544350
rect 129306 544294 129374 544350
rect 129430 544294 129498 544350
rect 129554 544294 129622 544350
rect 129678 544294 147250 544350
rect 147306 544294 147374 544350
rect 147430 544294 147498 544350
rect 147554 544294 147622 544350
rect 147678 544294 183250 544350
rect 183306 544294 183374 544350
rect 183430 544294 183498 544350
rect 183554 544294 183622 544350
rect 183678 544294 201250 544350
rect 201306 544294 201374 544350
rect 201430 544294 201498 544350
rect 201554 544294 201622 544350
rect 201678 544294 219250 544350
rect 219306 544294 219374 544350
rect 219430 544294 219498 544350
rect 219554 544294 219622 544350
rect 219678 544294 237250 544350
rect 237306 544294 237374 544350
rect 237430 544294 237498 544350
rect 237554 544294 237622 544350
rect 237678 544294 273250 544350
rect 273306 544294 273374 544350
rect 273430 544294 273498 544350
rect 273554 544294 273622 544350
rect 273678 544294 291250 544350
rect 291306 544294 291374 544350
rect 291430 544294 291498 544350
rect 291554 544294 291622 544350
rect 291678 544294 309250 544350
rect 309306 544294 309374 544350
rect 309430 544294 309498 544350
rect 309554 544294 309622 544350
rect 309678 544294 327250 544350
rect 327306 544294 327374 544350
rect 327430 544294 327498 544350
rect 327554 544294 327622 544350
rect 327678 544294 363250 544350
rect 363306 544294 363374 544350
rect 363430 544294 363498 544350
rect 363554 544294 363622 544350
rect 363678 544294 381250 544350
rect 381306 544294 381374 544350
rect 381430 544294 381498 544350
rect 381554 544294 381622 544350
rect 381678 544294 399250 544350
rect 399306 544294 399374 544350
rect 399430 544294 399498 544350
rect 399554 544294 399622 544350
rect 399678 544294 417250 544350
rect 417306 544294 417374 544350
rect 417430 544294 417498 544350
rect 417554 544294 417622 544350
rect 417678 544294 453250 544350
rect 453306 544294 453374 544350
rect 453430 544294 453498 544350
rect 453554 544294 453622 544350
rect 453678 544294 471250 544350
rect 471306 544294 471374 544350
rect 471430 544294 471498 544350
rect 471554 544294 471622 544350
rect 471678 544294 489250 544350
rect 489306 544294 489374 544350
rect 489430 544294 489498 544350
rect 489554 544294 489622 544350
rect 489678 544294 507250 544350
rect 507306 544294 507374 544350
rect 507430 544294 507498 544350
rect 507554 544294 507622 544350
rect 507678 544294 543250 544350
rect 543306 544294 543374 544350
rect 543430 544294 543498 544350
rect 543554 544294 543622 544350
rect 543678 544294 561250 544350
rect 561306 544294 561374 544350
rect 561430 544294 561498 544350
rect 561554 544294 561622 544350
rect 561678 544294 579250 544350
rect 579306 544294 579374 544350
rect 579430 544294 579498 544350
rect 579554 544294 579622 544350
rect 579678 544294 596496 544350
rect 596552 544294 596620 544350
rect 596676 544294 596744 544350
rect 596800 544294 596868 544350
rect 596924 544294 597980 544350
rect -1916 544226 597980 544294
rect -1916 544170 -860 544226
rect -804 544170 -736 544226
rect -680 544170 -612 544226
rect -556 544170 -488 544226
rect -432 544170 3250 544226
rect 3306 544170 3374 544226
rect 3430 544170 3498 544226
rect 3554 544170 3622 544226
rect 3678 544170 21250 544226
rect 21306 544170 21374 544226
rect 21430 544170 21498 544226
rect 21554 544170 21622 544226
rect 21678 544170 39250 544226
rect 39306 544170 39374 544226
rect 39430 544170 39498 544226
rect 39554 544170 39622 544226
rect 39678 544170 57250 544226
rect 57306 544170 57374 544226
rect 57430 544170 57498 544226
rect 57554 544170 57622 544226
rect 57678 544170 93250 544226
rect 93306 544170 93374 544226
rect 93430 544170 93498 544226
rect 93554 544170 93622 544226
rect 93678 544170 111250 544226
rect 111306 544170 111374 544226
rect 111430 544170 111498 544226
rect 111554 544170 111622 544226
rect 111678 544170 129250 544226
rect 129306 544170 129374 544226
rect 129430 544170 129498 544226
rect 129554 544170 129622 544226
rect 129678 544170 147250 544226
rect 147306 544170 147374 544226
rect 147430 544170 147498 544226
rect 147554 544170 147622 544226
rect 147678 544170 183250 544226
rect 183306 544170 183374 544226
rect 183430 544170 183498 544226
rect 183554 544170 183622 544226
rect 183678 544170 201250 544226
rect 201306 544170 201374 544226
rect 201430 544170 201498 544226
rect 201554 544170 201622 544226
rect 201678 544170 219250 544226
rect 219306 544170 219374 544226
rect 219430 544170 219498 544226
rect 219554 544170 219622 544226
rect 219678 544170 237250 544226
rect 237306 544170 237374 544226
rect 237430 544170 237498 544226
rect 237554 544170 237622 544226
rect 237678 544170 273250 544226
rect 273306 544170 273374 544226
rect 273430 544170 273498 544226
rect 273554 544170 273622 544226
rect 273678 544170 291250 544226
rect 291306 544170 291374 544226
rect 291430 544170 291498 544226
rect 291554 544170 291622 544226
rect 291678 544170 309250 544226
rect 309306 544170 309374 544226
rect 309430 544170 309498 544226
rect 309554 544170 309622 544226
rect 309678 544170 327250 544226
rect 327306 544170 327374 544226
rect 327430 544170 327498 544226
rect 327554 544170 327622 544226
rect 327678 544170 363250 544226
rect 363306 544170 363374 544226
rect 363430 544170 363498 544226
rect 363554 544170 363622 544226
rect 363678 544170 381250 544226
rect 381306 544170 381374 544226
rect 381430 544170 381498 544226
rect 381554 544170 381622 544226
rect 381678 544170 399250 544226
rect 399306 544170 399374 544226
rect 399430 544170 399498 544226
rect 399554 544170 399622 544226
rect 399678 544170 417250 544226
rect 417306 544170 417374 544226
rect 417430 544170 417498 544226
rect 417554 544170 417622 544226
rect 417678 544170 453250 544226
rect 453306 544170 453374 544226
rect 453430 544170 453498 544226
rect 453554 544170 453622 544226
rect 453678 544170 471250 544226
rect 471306 544170 471374 544226
rect 471430 544170 471498 544226
rect 471554 544170 471622 544226
rect 471678 544170 489250 544226
rect 489306 544170 489374 544226
rect 489430 544170 489498 544226
rect 489554 544170 489622 544226
rect 489678 544170 507250 544226
rect 507306 544170 507374 544226
rect 507430 544170 507498 544226
rect 507554 544170 507622 544226
rect 507678 544170 543250 544226
rect 543306 544170 543374 544226
rect 543430 544170 543498 544226
rect 543554 544170 543622 544226
rect 543678 544170 561250 544226
rect 561306 544170 561374 544226
rect 561430 544170 561498 544226
rect 561554 544170 561622 544226
rect 561678 544170 579250 544226
rect 579306 544170 579374 544226
rect 579430 544170 579498 544226
rect 579554 544170 579622 544226
rect 579678 544170 596496 544226
rect 596552 544170 596620 544226
rect 596676 544170 596744 544226
rect 596800 544170 596868 544226
rect 596924 544170 597980 544226
rect -1916 544102 597980 544170
rect -1916 544046 -860 544102
rect -804 544046 -736 544102
rect -680 544046 -612 544102
rect -556 544046 -488 544102
rect -432 544046 3250 544102
rect 3306 544046 3374 544102
rect 3430 544046 3498 544102
rect 3554 544046 3622 544102
rect 3678 544046 21250 544102
rect 21306 544046 21374 544102
rect 21430 544046 21498 544102
rect 21554 544046 21622 544102
rect 21678 544046 39250 544102
rect 39306 544046 39374 544102
rect 39430 544046 39498 544102
rect 39554 544046 39622 544102
rect 39678 544046 57250 544102
rect 57306 544046 57374 544102
rect 57430 544046 57498 544102
rect 57554 544046 57622 544102
rect 57678 544046 93250 544102
rect 93306 544046 93374 544102
rect 93430 544046 93498 544102
rect 93554 544046 93622 544102
rect 93678 544046 111250 544102
rect 111306 544046 111374 544102
rect 111430 544046 111498 544102
rect 111554 544046 111622 544102
rect 111678 544046 129250 544102
rect 129306 544046 129374 544102
rect 129430 544046 129498 544102
rect 129554 544046 129622 544102
rect 129678 544046 147250 544102
rect 147306 544046 147374 544102
rect 147430 544046 147498 544102
rect 147554 544046 147622 544102
rect 147678 544046 183250 544102
rect 183306 544046 183374 544102
rect 183430 544046 183498 544102
rect 183554 544046 183622 544102
rect 183678 544046 201250 544102
rect 201306 544046 201374 544102
rect 201430 544046 201498 544102
rect 201554 544046 201622 544102
rect 201678 544046 219250 544102
rect 219306 544046 219374 544102
rect 219430 544046 219498 544102
rect 219554 544046 219622 544102
rect 219678 544046 237250 544102
rect 237306 544046 237374 544102
rect 237430 544046 237498 544102
rect 237554 544046 237622 544102
rect 237678 544046 273250 544102
rect 273306 544046 273374 544102
rect 273430 544046 273498 544102
rect 273554 544046 273622 544102
rect 273678 544046 291250 544102
rect 291306 544046 291374 544102
rect 291430 544046 291498 544102
rect 291554 544046 291622 544102
rect 291678 544046 309250 544102
rect 309306 544046 309374 544102
rect 309430 544046 309498 544102
rect 309554 544046 309622 544102
rect 309678 544046 327250 544102
rect 327306 544046 327374 544102
rect 327430 544046 327498 544102
rect 327554 544046 327622 544102
rect 327678 544046 363250 544102
rect 363306 544046 363374 544102
rect 363430 544046 363498 544102
rect 363554 544046 363622 544102
rect 363678 544046 381250 544102
rect 381306 544046 381374 544102
rect 381430 544046 381498 544102
rect 381554 544046 381622 544102
rect 381678 544046 399250 544102
rect 399306 544046 399374 544102
rect 399430 544046 399498 544102
rect 399554 544046 399622 544102
rect 399678 544046 417250 544102
rect 417306 544046 417374 544102
rect 417430 544046 417498 544102
rect 417554 544046 417622 544102
rect 417678 544046 453250 544102
rect 453306 544046 453374 544102
rect 453430 544046 453498 544102
rect 453554 544046 453622 544102
rect 453678 544046 471250 544102
rect 471306 544046 471374 544102
rect 471430 544046 471498 544102
rect 471554 544046 471622 544102
rect 471678 544046 489250 544102
rect 489306 544046 489374 544102
rect 489430 544046 489498 544102
rect 489554 544046 489622 544102
rect 489678 544046 507250 544102
rect 507306 544046 507374 544102
rect 507430 544046 507498 544102
rect 507554 544046 507622 544102
rect 507678 544046 543250 544102
rect 543306 544046 543374 544102
rect 543430 544046 543498 544102
rect 543554 544046 543622 544102
rect 543678 544046 561250 544102
rect 561306 544046 561374 544102
rect 561430 544046 561498 544102
rect 561554 544046 561622 544102
rect 561678 544046 579250 544102
rect 579306 544046 579374 544102
rect 579430 544046 579498 544102
rect 579554 544046 579622 544102
rect 579678 544046 596496 544102
rect 596552 544046 596620 544102
rect 596676 544046 596744 544102
rect 596800 544046 596868 544102
rect 596924 544046 597980 544102
rect -1916 543978 597980 544046
rect -1916 543922 -860 543978
rect -804 543922 -736 543978
rect -680 543922 -612 543978
rect -556 543922 -488 543978
rect -432 543922 3250 543978
rect 3306 543922 3374 543978
rect 3430 543922 3498 543978
rect 3554 543922 3622 543978
rect 3678 543922 21250 543978
rect 21306 543922 21374 543978
rect 21430 543922 21498 543978
rect 21554 543922 21622 543978
rect 21678 543922 39250 543978
rect 39306 543922 39374 543978
rect 39430 543922 39498 543978
rect 39554 543922 39622 543978
rect 39678 543922 57250 543978
rect 57306 543922 57374 543978
rect 57430 543922 57498 543978
rect 57554 543922 57622 543978
rect 57678 543922 93250 543978
rect 93306 543922 93374 543978
rect 93430 543922 93498 543978
rect 93554 543922 93622 543978
rect 93678 543922 111250 543978
rect 111306 543922 111374 543978
rect 111430 543922 111498 543978
rect 111554 543922 111622 543978
rect 111678 543922 129250 543978
rect 129306 543922 129374 543978
rect 129430 543922 129498 543978
rect 129554 543922 129622 543978
rect 129678 543922 147250 543978
rect 147306 543922 147374 543978
rect 147430 543922 147498 543978
rect 147554 543922 147622 543978
rect 147678 543922 183250 543978
rect 183306 543922 183374 543978
rect 183430 543922 183498 543978
rect 183554 543922 183622 543978
rect 183678 543922 201250 543978
rect 201306 543922 201374 543978
rect 201430 543922 201498 543978
rect 201554 543922 201622 543978
rect 201678 543922 219250 543978
rect 219306 543922 219374 543978
rect 219430 543922 219498 543978
rect 219554 543922 219622 543978
rect 219678 543922 237250 543978
rect 237306 543922 237374 543978
rect 237430 543922 237498 543978
rect 237554 543922 237622 543978
rect 237678 543922 273250 543978
rect 273306 543922 273374 543978
rect 273430 543922 273498 543978
rect 273554 543922 273622 543978
rect 273678 543922 291250 543978
rect 291306 543922 291374 543978
rect 291430 543922 291498 543978
rect 291554 543922 291622 543978
rect 291678 543922 309250 543978
rect 309306 543922 309374 543978
rect 309430 543922 309498 543978
rect 309554 543922 309622 543978
rect 309678 543922 327250 543978
rect 327306 543922 327374 543978
rect 327430 543922 327498 543978
rect 327554 543922 327622 543978
rect 327678 543922 363250 543978
rect 363306 543922 363374 543978
rect 363430 543922 363498 543978
rect 363554 543922 363622 543978
rect 363678 543922 381250 543978
rect 381306 543922 381374 543978
rect 381430 543922 381498 543978
rect 381554 543922 381622 543978
rect 381678 543922 399250 543978
rect 399306 543922 399374 543978
rect 399430 543922 399498 543978
rect 399554 543922 399622 543978
rect 399678 543922 417250 543978
rect 417306 543922 417374 543978
rect 417430 543922 417498 543978
rect 417554 543922 417622 543978
rect 417678 543922 453250 543978
rect 453306 543922 453374 543978
rect 453430 543922 453498 543978
rect 453554 543922 453622 543978
rect 453678 543922 471250 543978
rect 471306 543922 471374 543978
rect 471430 543922 471498 543978
rect 471554 543922 471622 543978
rect 471678 543922 489250 543978
rect 489306 543922 489374 543978
rect 489430 543922 489498 543978
rect 489554 543922 489622 543978
rect 489678 543922 507250 543978
rect 507306 543922 507374 543978
rect 507430 543922 507498 543978
rect 507554 543922 507622 543978
rect 507678 543922 543250 543978
rect 543306 543922 543374 543978
rect 543430 543922 543498 543978
rect 543554 543922 543622 543978
rect 543678 543922 561250 543978
rect 561306 543922 561374 543978
rect 561430 543922 561498 543978
rect 561554 543922 561622 543978
rect 561678 543922 579250 543978
rect 579306 543922 579374 543978
rect 579430 543922 579498 543978
rect 579554 543922 579622 543978
rect 579678 543922 596496 543978
rect 596552 543922 596620 543978
rect 596676 543922 596744 543978
rect 596800 543922 596868 543978
rect 596924 543922 597980 543978
rect -1916 543826 597980 543922
rect -1916 532350 597980 532446
rect -1916 532294 -1820 532350
rect -1764 532294 -1696 532350
rect -1640 532294 -1572 532350
rect -1516 532294 -1448 532350
rect -1392 532294 6970 532350
rect 7026 532294 7094 532350
rect 7150 532294 7218 532350
rect 7274 532294 7342 532350
rect 7398 532294 24970 532350
rect 25026 532294 25094 532350
rect 25150 532294 25218 532350
rect 25274 532294 25342 532350
rect 25398 532294 42970 532350
rect 43026 532294 43094 532350
rect 43150 532294 43218 532350
rect 43274 532294 43342 532350
rect 43398 532294 60970 532350
rect 61026 532294 61094 532350
rect 61150 532294 61218 532350
rect 61274 532294 61342 532350
rect 61398 532294 78970 532350
rect 79026 532294 79094 532350
rect 79150 532294 79218 532350
rect 79274 532294 79342 532350
rect 79398 532294 96970 532350
rect 97026 532294 97094 532350
rect 97150 532294 97218 532350
rect 97274 532294 97342 532350
rect 97398 532294 132970 532350
rect 133026 532294 133094 532350
rect 133150 532294 133218 532350
rect 133274 532294 133342 532350
rect 133398 532294 150970 532350
rect 151026 532294 151094 532350
rect 151150 532294 151218 532350
rect 151274 532294 151342 532350
rect 151398 532294 168970 532350
rect 169026 532294 169094 532350
rect 169150 532294 169218 532350
rect 169274 532294 169342 532350
rect 169398 532294 186970 532350
rect 187026 532294 187094 532350
rect 187150 532294 187218 532350
rect 187274 532294 187342 532350
rect 187398 532294 222970 532350
rect 223026 532294 223094 532350
rect 223150 532294 223218 532350
rect 223274 532294 223342 532350
rect 223398 532294 240970 532350
rect 241026 532294 241094 532350
rect 241150 532294 241218 532350
rect 241274 532294 241342 532350
rect 241398 532294 258970 532350
rect 259026 532294 259094 532350
rect 259150 532294 259218 532350
rect 259274 532294 259342 532350
rect 259398 532294 276970 532350
rect 277026 532294 277094 532350
rect 277150 532294 277218 532350
rect 277274 532294 277342 532350
rect 277398 532294 312970 532350
rect 313026 532294 313094 532350
rect 313150 532294 313218 532350
rect 313274 532294 313342 532350
rect 313398 532294 330970 532350
rect 331026 532294 331094 532350
rect 331150 532294 331218 532350
rect 331274 532294 331342 532350
rect 331398 532294 348970 532350
rect 349026 532294 349094 532350
rect 349150 532294 349218 532350
rect 349274 532294 349342 532350
rect 349398 532294 366970 532350
rect 367026 532294 367094 532350
rect 367150 532294 367218 532350
rect 367274 532294 367342 532350
rect 367398 532294 402970 532350
rect 403026 532294 403094 532350
rect 403150 532294 403218 532350
rect 403274 532294 403342 532350
rect 403398 532294 420970 532350
rect 421026 532294 421094 532350
rect 421150 532294 421218 532350
rect 421274 532294 421342 532350
rect 421398 532294 438970 532350
rect 439026 532294 439094 532350
rect 439150 532294 439218 532350
rect 439274 532294 439342 532350
rect 439398 532294 456970 532350
rect 457026 532294 457094 532350
rect 457150 532294 457218 532350
rect 457274 532294 457342 532350
rect 457398 532294 492970 532350
rect 493026 532294 493094 532350
rect 493150 532294 493218 532350
rect 493274 532294 493342 532350
rect 493398 532294 510970 532350
rect 511026 532294 511094 532350
rect 511150 532294 511218 532350
rect 511274 532294 511342 532350
rect 511398 532294 528970 532350
rect 529026 532294 529094 532350
rect 529150 532294 529218 532350
rect 529274 532294 529342 532350
rect 529398 532294 546970 532350
rect 547026 532294 547094 532350
rect 547150 532294 547218 532350
rect 547274 532294 547342 532350
rect 547398 532294 564970 532350
rect 565026 532294 565094 532350
rect 565150 532294 565218 532350
rect 565274 532294 565342 532350
rect 565398 532294 582970 532350
rect 583026 532294 583094 532350
rect 583150 532294 583218 532350
rect 583274 532294 583342 532350
rect 583398 532294 597456 532350
rect 597512 532294 597580 532350
rect 597636 532294 597704 532350
rect 597760 532294 597828 532350
rect 597884 532294 597980 532350
rect -1916 532226 597980 532294
rect -1916 532170 -1820 532226
rect -1764 532170 -1696 532226
rect -1640 532170 -1572 532226
rect -1516 532170 -1448 532226
rect -1392 532170 6970 532226
rect 7026 532170 7094 532226
rect 7150 532170 7218 532226
rect 7274 532170 7342 532226
rect 7398 532170 24970 532226
rect 25026 532170 25094 532226
rect 25150 532170 25218 532226
rect 25274 532170 25342 532226
rect 25398 532170 42970 532226
rect 43026 532170 43094 532226
rect 43150 532170 43218 532226
rect 43274 532170 43342 532226
rect 43398 532170 60970 532226
rect 61026 532170 61094 532226
rect 61150 532170 61218 532226
rect 61274 532170 61342 532226
rect 61398 532170 78970 532226
rect 79026 532170 79094 532226
rect 79150 532170 79218 532226
rect 79274 532170 79342 532226
rect 79398 532170 96970 532226
rect 97026 532170 97094 532226
rect 97150 532170 97218 532226
rect 97274 532170 97342 532226
rect 97398 532170 132970 532226
rect 133026 532170 133094 532226
rect 133150 532170 133218 532226
rect 133274 532170 133342 532226
rect 133398 532170 150970 532226
rect 151026 532170 151094 532226
rect 151150 532170 151218 532226
rect 151274 532170 151342 532226
rect 151398 532170 168970 532226
rect 169026 532170 169094 532226
rect 169150 532170 169218 532226
rect 169274 532170 169342 532226
rect 169398 532170 186970 532226
rect 187026 532170 187094 532226
rect 187150 532170 187218 532226
rect 187274 532170 187342 532226
rect 187398 532170 222970 532226
rect 223026 532170 223094 532226
rect 223150 532170 223218 532226
rect 223274 532170 223342 532226
rect 223398 532170 240970 532226
rect 241026 532170 241094 532226
rect 241150 532170 241218 532226
rect 241274 532170 241342 532226
rect 241398 532170 258970 532226
rect 259026 532170 259094 532226
rect 259150 532170 259218 532226
rect 259274 532170 259342 532226
rect 259398 532170 276970 532226
rect 277026 532170 277094 532226
rect 277150 532170 277218 532226
rect 277274 532170 277342 532226
rect 277398 532170 312970 532226
rect 313026 532170 313094 532226
rect 313150 532170 313218 532226
rect 313274 532170 313342 532226
rect 313398 532170 330970 532226
rect 331026 532170 331094 532226
rect 331150 532170 331218 532226
rect 331274 532170 331342 532226
rect 331398 532170 348970 532226
rect 349026 532170 349094 532226
rect 349150 532170 349218 532226
rect 349274 532170 349342 532226
rect 349398 532170 366970 532226
rect 367026 532170 367094 532226
rect 367150 532170 367218 532226
rect 367274 532170 367342 532226
rect 367398 532170 402970 532226
rect 403026 532170 403094 532226
rect 403150 532170 403218 532226
rect 403274 532170 403342 532226
rect 403398 532170 420970 532226
rect 421026 532170 421094 532226
rect 421150 532170 421218 532226
rect 421274 532170 421342 532226
rect 421398 532170 438970 532226
rect 439026 532170 439094 532226
rect 439150 532170 439218 532226
rect 439274 532170 439342 532226
rect 439398 532170 456970 532226
rect 457026 532170 457094 532226
rect 457150 532170 457218 532226
rect 457274 532170 457342 532226
rect 457398 532170 492970 532226
rect 493026 532170 493094 532226
rect 493150 532170 493218 532226
rect 493274 532170 493342 532226
rect 493398 532170 510970 532226
rect 511026 532170 511094 532226
rect 511150 532170 511218 532226
rect 511274 532170 511342 532226
rect 511398 532170 528970 532226
rect 529026 532170 529094 532226
rect 529150 532170 529218 532226
rect 529274 532170 529342 532226
rect 529398 532170 546970 532226
rect 547026 532170 547094 532226
rect 547150 532170 547218 532226
rect 547274 532170 547342 532226
rect 547398 532170 564970 532226
rect 565026 532170 565094 532226
rect 565150 532170 565218 532226
rect 565274 532170 565342 532226
rect 565398 532170 582970 532226
rect 583026 532170 583094 532226
rect 583150 532170 583218 532226
rect 583274 532170 583342 532226
rect 583398 532170 597456 532226
rect 597512 532170 597580 532226
rect 597636 532170 597704 532226
rect 597760 532170 597828 532226
rect 597884 532170 597980 532226
rect -1916 532102 597980 532170
rect -1916 532046 -1820 532102
rect -1764 532046 -1696 532102
rect -1640 532046 -1572 532102
rect -1516 532046 -1448 532102
rect -1392 532046 6970 532102
rect 7026 532046 7094 532102
rect 7150 532046 7218 532102
rect 7274 532046 7342 532102
rect 7398 532046 24970 532102
rect 25026 532046 25094 532102
rect 25150 532046 25218 532102
rect 25274 532046 25342 532102
rect 25398 532046 42970 532102
rect 43026 532046 43094 532102
rect 43150 532046 43218 532102
rect 43274 532046 43342 532102
rect 43398 532046 60970 532102
rect 61026 532046 61094 532102
rect 61150 532046 61218 532102
rect 61274 532046 61342 532102
rect 61398 532046 78970 532102
rect 79026 532046 79094 532102
rect 79150 532046 79218 532102
rect 79274 532046 79342 532102
rect 79398 532046 96970 532102
rect 97026 532046 97094 532102
rect 97150 532046 97218 532102
rect 97274 532046 97342 532102
rect 97398 532046 132970 532102
rect 133026 532046 133094 532102
rect 133150 532046 133218 532102
rect 133274 532046 133342 532102
rect 133398 532046 150970 532102
rect 151026 532046 151094 532102
rect 151150 532046 151218 532102
rect 151274 532046 151342 532102
rect 151398 532046 168970 532102
rect 169026 532046 169094 532102
rect 169150 532046 169218 532102
rect 169274 532046 169342 532102
rect 169398 532046 186970 532102
rect 187026 532046 187094 532102
rect 187150 532046 187218 532102
rect 187274 532046 187342 532102
rect 187398 532046 222970 532102
rect 223026 532046 223094 532102
rect 223150 532046 223218 532102
rect 223274 532046 223342 532102
rect 223398 532046 240970 532102
rect 241026 532046 241094 532102
rect 241150 532046 241218 532102
rect 241274 532046 241342 532102
rect 241398 532046 258970 532102
rect 259026 532046 259094 532102
rect 259150 532046 259218 532102
rect 259274 532046 259342 532102
rect 259398 532046 276970 532102
rect 277026 532046 277094 532102
rect 277150 532046 277218 532102
rect 277274 532046 277342 532102
rect 277398 532046 312970 532102
rect 313026 532046 313094 532102
rect 313150 532046 313218 532102
rect 313274 532046 313342 532102
rect 313398 532046 330970 532102
rect 331026 532046 331094 532102
rect 331150 532046 331218 532102
rect 331274 532046 331342 532102
rect 331398 532046 348970 532102
rect 349026 532046 349094 532102
rect 349150 532046 349218 532102
rect 349274 532046 349342 532102
rect 349398 532046 366970 532102
rect 367026 532046 367094 532102
rect 367150 532046 367218 532102
rect 367274 532046 367342 532102
rect 367398 532046 402970 532102
rect 403026 532046 403094 532102
rect 403150 532046 403218 532102
rect 403274 532046 403342 532102
rect 403398 532046 420970 532102
rect 421026 532046 421094 532102
rect 421150 532046 421218 532102
rect 421274 532046 421342 532102
rect 421398 532046 438970 532102
rect 439026 532046 439094 532102
rect 439150 532046 439218 532102
rect 439274 532046 439342 532102
rect 439398 532046 456970 532102
rect 457026 532046 457094 532102
rect 457150 532046 457218 532102
rect 457274 532046 457342 532102
rect 457398 532046 492970 532102
rect 493026 532046 493094 532102
rect 493150 532046 493218 532102
rect 493274 532046 493342 532102
rect 493398 532046 510970 532102
rect 511026 532046 511094 532102
rect 511150 532046 511218 532102
rect 511274 532046 511342 532102
rect 511398 532046 528970 532102
rect 529026 532046 529094 532102
rect 529150 532046 529218 532102
rect 529274 532046 529342 532102
rect 529398 532046 546970 532102
rect 547026 532046 547094 532102
rect 547150 532046 547218 532102
rect 547274 532046 547342 532102
rect 547398 532046 564970 532102
rect 565026 532046 565094 532102
rect 565150 532046 565218 532102
rect 565274 532046 565342 532102
rect 565398 532046 582970 532102
rect 583026 532046 583094 532102
rect 583150 532046 583218 532102
rect 583274 532046 583342 532102
rect 583398 532046 597456 532102
rect 597512 532046 597580 532102
rect 597636 532046 597704 532102
rect 597760 532046 597828 532102
rect 597884 532046 597980 532102
rect -1916 531978 597980 532046
rect -1916 531922 -1820 531978
rect -1764 531922 -1696 531978
rect -1640 531922 -1572 531978
rect -1516 531922 -1448 531978
rect -1392 531922 6970 531978
rect 7026 531922 7094 531978
rect 7150 531922 7218 531978
rect 7274 531922 7342 531978
rect 7398 531922 24970 531978
rect 25026 531922 25094 531978
rect 25150 531922 25218 531978
rect 25274 531922 25342 531978
rect 25398 531922 42970 531978
rect 43026 531922 43094 531978
rect 43150 531922 43218 531978
rect 43274 531922 43342 531978
rect 43398 531922 60970 531978
rect 61026 531922 61094 531978
rect 61150 531922 61218 531978
rect 61274 531922 61342 531978
rect 61398 531922 78970 531978
rect 79026 531922 79094 531978
rect 79150 531922 79218 531978
rect 79274 531922 79342 531978
rect 79398 531922 96970 531978
rect 97026 531922 97094 531978
rect 97150 531922 97218 531978
rect 97274 531922 97342 531978
rect 97398 531922 132970 531978
rect 133026 531922 133094 531978
rect 133150 531922 133218 531978
rect 133274 531922 133342 531978
rect 133398 531922 150970 531978
rect 151026 531922 151094 531978
rect 151150 531922 151218 531978
rect 151274 531922 151342 531978
rect 151398 531922 168970 531978
rect 169026 531922 169094 531978
rect 169150 531922 169218 531978
rect 169274 531922 169342 531978
rect 169398 531922 186970 531978
rect 187026 531922 187094 531978
rect 187150 531922 187218 531978
rect 187274 531922 187342 531978
rect 187398 531922 222970 531978
rect 223026 531922 223094 531978
rect 223150 531922 223218 531978
rect 223274 531922 223342 531978
rect 223398 531922 240970 531978
rect 241026 531922 241094 531978
rect 241150 531922 241218 531978
rect 241274 531922 241342 531978
rect 241398 531922 258970 531978
rect 259026 531922 259094 531978
rect 259150 531922 259218 531978
rect 259274 531922 259342 531978
rect 259398 531922 276970 531978
rect 277026 531922 277094 531978
rect 277150 531922 277218 531978
rect 277274 531922 277342 531978
rect 277398 531922 312970 531978
rect 313026 531922 313094 531978
rect 313150 531922 313218 531978
rect 313274 531922 313342 531978
rect 313398 531922 330970 531978
rect 331026 531922 331094 531978
rect 331150 531922 331218 531978
rect 331274 531922 331342 531978
rect 331398 531922 348970 531978
rect 349026 531922 349094 531978
rect 349150 531922 349218 531978
rect 349274 531922 349342 531978
rect 349398 531922 366970 531978
rect 367026 531922 367094 531978
rect 367150 531922 367218 531978
rect 367274 531922 367342 531978
rect 367398 531922 402970 531978
rect 403026 531922 403094 531978
rect 403150 531922 403218 531978
rect 403274 531922 403342 531978
rect 403398 531922 420970 531978
rect 421026 531922 421094 531978
rect 421150 531922 421218 531978
rect 421274 531922 421342 531978
rect 421398 531922 438970 531978
rect 439026 531922 439094 531978
rect 439150 531922 439218 531978
rect 439274 531922 439342 531978
rect 439398 531922 456970 531978
rect 457026 531922 457094 531978
rect 457150 531922 457218 531978
rect 457274 531922 457342 531978
rect 457398 531922 492970 531978
rect 493026 531922 493094 531978
rect 493150 531922 493218 531978
rect 493274 531922 493342 531978
rect 493398 531922 510970 531978
rect 511026 531922 511094 531978
rect 511150 531922 511218 531978
rect 511274 531922 511342 531978
rect 511398 531922 528970 531978
rect 529026 531922 529094 531978
rect 529150 531922 529218 531978
rect 529274 531922 529342 531978
rect 529398 531922 546970 531978
rect 547026 531922 547094 531978
rect 547150 531922 547218 531978
rect 547274 531922 547342 531978
rect 547398 531922 564970 531978
rect 565026 531922 565094 531978
rect 565150 531922 565218 531978
rect 565274 531922 565342 531978
rect 565398 531922 582970 531978
rect 583026 531922 583094 531978
rect 583150 531922 583218 531978
rect 583274 531922 583342 531978
rect 583398 531922 597456 531978
rect 597512 531922 597580 531978
rect 597636 531922 597704 531978
rect 597760 531922 597828 531978
rect 597884 531922 597980 531978
rect -1916 531826 597980 531922
rect -1916 526350 597980 526446
rect -1916 526294 -860 526350
rect -804 526294 -736 526350
rect -680 526294 -612 526350
rect -556 526294 -488 526350
rect -432 526294 3250 526350
rect 3306 526294 3374 526350
rect 3430 526294 3498 526350
rect 3554 526294 3622 526350
rect 3678 526294 21250 526350
rect 21306 526294 21374 526350
rect 21430 526294 21498 526350
rect 21554 526294 21622 526350
rect 21678 526294 39250 526350
rect 39306 526294 39374 526350
rect 39430 526294 39498 526350
rect 39554 526294 39622 526350
rect 39678 526294 57250 526350
rect 57306 526294 57374 526350
rect 57430 526294 57498 526350
rect 57554 526294 57622 526350
rect 57678 526294 93250 526350
rect 93306 526294 93374 526350
rect 93430 526294 93498 526350
rect 93554 526294 93622 526350
rect 93678 526294 111250 526350
rect 111306 526294 111374 526350
rect 111430 526294 111498 526350
rect 111554 526294 111622 526350
rect 111678 526294 129250 526350
rect 129306 526294 129374 526350
rect 129430 526294 129498 526350
rect 129554 526294 129622 526350
rect 129678 526294 147250 526350
rect 147306 526294 147374 526350
rect 147430 526294 147498 526350
rect 147554 526294 147622 526350
rect 147678 526294 183250 526350
rect 183306 526294 183374 526350
rect 183430 526294 183498 526350
rect 183554 526294 183622 526350
rect 183678 526294 201250 526350
rect 201306 526294 201374 526350
rect 201430 526294 201498 526350
rect 201554 526294 201622 526350
rect 201678 526294 219250 526350
rect 219306 526294 219374 526350
rect 219430 526294 219498 526350
rect 219554 526294 219622 526350
rect 219678 526294 237250 526350
rect 237306 526294 237374 526350
rect 237430 526294 237498 526350
rect 237554 526294 237622 526350
rect 237678 526294 273250 526350
rect 273306 526294 273374 526350
rect 273430 526294 273498 526350
rect 273554 526294 273622 526350
rect 273678 526294 291250 526350
rect 291306 526294 291374 526350
rect 291430 526294 291498 526350
rect 291554 526294 291622 526350
rect 291678 526294 309250 526350
rect 309306 526294 309374 526350
rect 309430 526294 309498 526350
rect 309554 526294 309622 526350
rect 309678 526294 327250 526350
rect 327306 526294 327374 526350
rect 327430 526294 327498 526350
rect 327554 526294 327622 526350
rect 327678 526294 363250 526350
rect 363306 526294 363374 526350
rect 363430 526294 363498 526350
rect 363554 526294 363622 526350
rect 363678 526294 381250 526350
rect 381306 526294 381374 526350
rect 381430 526294 381498 526350
rect 381554 526294 381622 526350
rect 381678 526294 399250 526350
rect 399306 526294 399374 526350
rect 399430 526294 399498 526350
rect 399554 526294 399622 526350
rect 399678 526294 417250 526350
rect 417306 526294 417374 526350
rect 417430 526294 417498 526350
rect 417554 526294 417622 526350
rect 417678 526294 453250 526350
rect 453306 526294 453374 526350
rect 453430 526294 453498 526350
rect 453554 526294 453622 526350
rect 453678 526294 471250 526350
rect 471306 526294 471374 526350
rect 471430 526294 471498 526350
rect 471554 526294 471622 526350
rect 471678 526294 489250 526350
rect 489306 526294 489374 526350
rect 489430 526294 489498 526350
rect 489554 526294 489622 526350
rect 489678 526294 507250 526350
rect 507306 526294 507374 526350
rect 507430 526294 507498 526350
rect 507554 526294 507622 526350
rect 507678 526294 543250 526350
rect 543306 526294 543374 526350
rect 543430 526294 543498 526350
rect 543554 526294 543622 526350
rect 543678 526294 561250 526350
rect 561306 526294 561374 526350
rect 561430 526294 561498 526350
rect 561554 526294 561622 526350
rect 561678 526294 579250 526350
rect 579306 526294 579374 526350
rect 579430 526294 579498 526350
rect 579554 526294 579622 526350
rect 579678 526294 596496 526350
rect 596552 526294 596620 526350
rect 596676 526294 596744 526350
rect 596800 526294 596868 526350
rect 596924 526294 597980 526350
rect -1916 526226 597980 526294
rect -1916 526170 -860 526226
rect -804 526170 -736 526226
rect -680 526170 -612 526226
rect -556 526170 -488 526226
rect -432 526170 3250 526226
rect 3306 526170 3374 526226
rect 3430 526170 3498 526226
rect 3554 526170 3622 526226
rect 3678 526170 21250 526226
rect 21306 526170 21374 526226
rect 21430 526170 21498 526226
rect 21554 526170 21622 526226
rect 21678 526170 39250 526226
rect 39306 526170 39374 526226
rect 39430 526170 39498 526226
rect 39554 526170 39622 526226
rect 39678 526170 57250 526226
rect 57306 526170 57374 526226
rect 57430 526170 57498 526226
rect 57554 526170 57622 526226
rect 57678 526170 93250 526226
rect 93306 526170 93374 526226
rect 93430 526170 93498 526226
rect 93554 526170 93622 526226
rect 93678 526170 111250 526226
rect 111306 526170 111374 526226
rect 111430 526170 111498 526226
rect 111554 526170 111622 526226
rect 111678 526170 129250 526226
rect 129306 526170 129374 526226
rect 129430 526170 129498 526226
rect 129554 526170 129622 526226
rect 129678 526170 147250 526226
rect 147306 526170 147374 526226
rect 147430 526170 147498 526226
rect 147554 526170 147622 526226
rect 147678 526170 183250 526226
rect 183306 526170 183374 526226
rect 183430 526170 183498 526226
rect 183554 526170 183622 526226
rect 183678 526170 201250 526226
rect 201306 526170 201374 526226
rect 201430 526170 201498 526226
rect 201554 526170 201622 526226
rect 201678 526170 219250 526226
rect 219306 526170 219374 526226
rect 219430 526170 219498 526226
rect 219554 526170 219622 526226
rect 219678 526170 237250 526226
rect 237306 526170 237374 526226
rect 237430 526170 237498 526226
rect 237554 526170 237622 526226
rect 237678 526170 273250 526226
rect 273306 526170 273374 526226
rect 273430 526170 273498 526226
rect 273554 526170 273622 526226
rect 273678 526170 291250 526226
rect 291306 526170 291374 526226
rect 291430 526170 291498 526226
rect 291554 526170 291622 526226
rect 291678 526170 309250 526226
rect 309306 526170 309374 526226
rect 309430 526170 309498 526226
rect 309554 526170 309622 526226
rect 309678 526170 327250 526226
rect 327306 526170 327374 526226
rect 327430 526170 327498 526226
rect 327554 526170 327622 526226
rect 327678 526170 363250 526226
rect 363306 526170 363374 526226
rect 363430 526170 363498 526226
rect 363554 526170 363622 526226
rect 363678 526170 381250 526226
rect 381306 526170 381374 526226
rect 381430 526170 381498 526226
rect 381554 526170 381622 526226
rect 381678 526170 399250 526226
rect 399306 526170 399374 526226
rect 399430 526170 399498 526226
rect 399554 526170 399622 526226
rect 399678 526170 417250 526226
rect 417306 526170 417374 526226
rect 417430 526170 417498 526226
rect 417554 526170 417622 526226
rect 417678 526170 453250 526226
rect 453306 526170 453374 526226
rect 453430 526170 453498 526226
rect 453554 526170 453622 526226
rect 453678 526170 471250 526226
rect 471306 526170 471374 526226
rect 471430 526170 471498 526226
rect 471554 526170 471622 526226
rect 471678 526170 489250 526226
rect 489306 526170 489374 526226
rect 489430 526170 489498 526226
rect 489554 526170 489622 526226
rect 489678 526170 507250 526226
rect 507306 526170 507374 526226
rect 507430 526170 507498 526226
rect 507554 526170 507622 526226
rect 507678 526170 543250 526226
rect 543306 526170 543374 526226
rect 543430 526170 543498 526226
rect 543554 526170 543622 526226
rect 543678 526170 561250 526226
rect 561306 526170 561374 526226
rect 561430 526170 561498 526226
rect 561554 526170 561622 526226
rect 561678 526170 579250 526226
rect 579306 526170 579374 526226
rect 579430 526170 579498 526226
rect 579554 526170 579622 526226
rect 579678 526170 596496 526226
rect 596552 526170 596620 526226
rect 596676 526170 596744 526226
rect 596800 526170 596868 526226
rect 596924 526170 597980 526226
rect -1916 526102 597980 526170
rect -1916 526046 -860 526102
rect -804 526046 -736 526102
rect -680 526046 -612 526102
rect -556 526046 -488 526102
rect -432 526046 3250 526102
rect 3306 526046 3374 526102
rect 3430 526046 3498 526102
rect 3554 526046 3622 526102
rect 3678 526046 21250 526102
rect 21306 526046 21374 526102
rect 21430 526046 21498 526102
rect 21554 526046 21622 526102
rect 21678 526046 39250 526102
rect 39306 526046 39374 526102
rect 39430 526046 39498 526102
rect 39554 526046 39622 526102
rect 39678 526046 57250 526102
rect 57306 526046 57374 526102
rect 57430 526046 57498 526102
rect 57554 526046 57622 526102
rect 57678 526046 93250 526102
rect 93306 526046 93374 526102
rect 93430 526046 93498 526102
rect 93554 526046 93622 526102
rect 93678 526046 111250 526102
rect 111306 526046 111374 526102
rect 111430 526046 111498 526102
rect 111554 526046 111622 526102
rect 111678 526046 129250 526102
rect 129306 526046 129374 526102
rect 129430 526046 129498 526102
rect 129554 526046 129622 526102
rect 129678 526046 147250 526102
rect 147306 526046 147374 526102
rect 147430 526046 147498 526102
rect 147554 526046 147622 526102
rect 147678 526046 183250 526102
rect 183306 526046 183374 526102
rect 183430 526046 183498 526102
rect 183554 526046 183622 526102
rect 183678 526046 201250 526102
rect 201306 526046 201374 526102
rect 201430 526046 201498 526102
rect 201554 526046 201622 526102
rect 201678 526046 219250 526102
rect 219306 526046 219374 526102
rect 219430 526046 219498 526102
rect 219554 526046 219622 526102
rect 219678 526046 237250 526102
rect 237306 526046 237374 526102
rect 237430 526046 237498 526102
rect 237554 526046 237622 526102
rect 237678 526046 273250 526102
rect 273306 526046 273374 526102
rect 273430 526046 273498 526102
rect 273554 526046 273622 526102
rect 273678 526046 291250 526102
rect 291306 526046 291374 526102
rect 291430 526046 291498 526102
rect 291554 526046 291622 526102
rect 291678 526046 309250 526102
rect 309306 526046 309374 526102
rect 309430 526046 309498 526102
rect 309554 526046 309622 526102
rect 309678 526046 327250 526102
rect 327306 526046 327374 526102
rect 327430 526046 327498 526102
rect 327554 526046 327622 526102
rect 327678 526046 363250 526102
rect 363306 526046 363374 526102
rect 363430 526046 363498 526102
rect 363554 526046 363622 526102
rect 363678 526046 381250 526102
rect 381306 526046 381374 526102
rect 381430 526046 381498 526102
rect 381554 526046 381622 526102
rect 381678 526046 399250 526102
rect 399306 526046 399374 526102
rect 399430 526046 399498 526102
rect 399554 526046 399622 526102
rect 399678 526046 417250 526102
rect 417306 526046 417374 526102
rect 417430 526046 417498 526102
rect 417554 526046 417622 526102
rect 417678 526046 453250 526102
rect 453306 526046 453374 526102
rect 453430 526046 453498 526102
rect 453554 526046 453622 526102
rect 453678 526046 471250 526102
rect 471306 526046 471374 526102
rect 471430 526046 471498 526102
rect 471554 526046 471622 526102
rect 471678 526046 489250 526102
rect 489306 526046 489374 526102
rect 489430 526046 489498 526102
rect 489554 526046 489622 526102
rect 489678 526046 507250 526102
rect 507306 526046 507374 526102
rect 507430 526046 507498 526102
rect 507554 526046 507622 526102
rect 507678 526046 543250 526102
rect 543306 526046 543374 526102
rect 543430 526046 543498 526102
rect 543554 526046 543622 526102
rect 543678 526046 561250 526102
rect 561306 526046 561374 526102
rect 561430 526046 561498 526102
rect 561554 526046 561622 526102
rect 561678 526046 579250 526102
rect 579306 526046 579374 526102
rect 579430 526046 579498 526102
rect 579554 526046 579622 526102
rect 579678 526046 596496 526102
rect 596552 526046 596620 526102
rect 596676 526046 596744 526102
rect 596800 526046 596868 526102
rect 596924 526046 597980 526102
rect -1916 525978 597980 526046
rect -1916 525922 -860 525978
rect -804 525922 -736 525978
rect -680 525922 -612 525978
rect -556 525922 -488 525978
rect -432 525922 3250 525978
rect 3306 525922 3374 525978
rect 3430 525922 3498 525978
rect 3554 525922 3622 525978
rect 3678 525922 21250 525978
rect 21306 525922 21374 525978
rect 21430 525922 21498 525978
rect 21554 525922 21622 525978
rect 21678 525922 39250 525978
rect 39306 525922 39374 525978
rect 39430 525922 39498 525978
rect 39554 525922 39622 525978
rect 39678 525922 57250 525978
rect 57306 525922 57374 525978
rect 57430 525922 57498 525978
rect 57554 525922 57622 525978
rect 57678 525922 93250 525978
rect 93306 525922 93374 525978
rect 93430 525922 93498 525978
rect 93554 525922 93622 525978
rect 93678 525922 111250 525978
rect 111306 525922 111374 525978
rect 111430 525922 111498 525978
rect 111554 525922 111622 525978
rect 111678 525922 129250 525978
rect 129306 525922 129374 525978
rect 129430 525922 129498 525978
rect 129554 525922 129622 525978
rect 129678 525922 147250 525978
rect 147306 525922 147374 525978
rect 147430 525922 147498 525978
rect 147554 525922 147622 525978
rect 147678 525922 183250 525978
rect 183306 525922 183374 525978
rect 183430 525922 183498 525978
rect 183554 525922 183622 525978
rect 183678 525922 201250 525978
rect 201306 525922 201374 525978
rect 201430 525922 201498 525978
rect 201554 525922 201622 525978
rect 201678 525922 219250 525978
rect 219306 525922 219374 525978
rect 219430 525922 219498 525978
rect 219554 525922 219622 525978
rect 219678 525922 237250 525978
rect 237306 525922 237374 525978
rect 237430 525922 237498 525978
rect 237554 525922 237622 525978
rect 237678 525922 273250 525978
rect 273306 525922 273374 525978
rect 273430 525922 273498 525978
rect 273554 525922 273622 525978
rect 273678 525922 291250 525978
rect 291306 525922 291374 525978
rect 291430 525922 291498 525978
rect 291554 525922 291622 525978
rect 291678 525922 309250 525978
rect 309306 525922 309374 525978
rect 309430 525922 309498 525978
rect 309554 525922 309622 525978
rect 309678 525922 327250 525978
rect 327306 525922 327374 525978
rect 327430 525922 327498 525978
rect 327554 525922 327622 525978
rect 327678 525922 363250 525978
rect 363306 525922 363374 525978
rect 363430 525922 363498 525978
rect 363554 525922 363622 525978
rect 363678 525922 381250 525978
rect 381306 525922 381374 525978
rect 381430 525922 381498 525978
rect 381554 525922 381622 525978
rect 381678 525922 399250 525978
rect 399306 525922 399374 525978
rect 399430 525922 399498 525978
rect 399554 525922 399622 525978
rect 399678 525922 417250 525978
rect 417306 525922 417374 525978
rect 417430 525922 417498 525978
rect 417554 525922 417622 525978
rect 417678 525922 453250 525978
rect 453306 525922 453374 525978
rect 453430 525922 453498 525978
rect 453554 525922 453622 525978
rect 453678 525922 471250 525978
rect 471306 525922 471374 525978
rect 471430 525922 471498 525978
rect 471554 525922 471622 525978
rect 471678 525922 489250 525978
rect 489306 525922 489374 525978
rect 489430 525922 489498 525978
rect 489554 525922 489622 525978
rect 489678 525922 507250 525978
rect 507306 525922 507374 525978
rect 507430 525922 507498 525978
rect 507554 525922 507622 525978
rect 507678 525922 543250 525978
rect 543306 525922 543374 525978
rect 543430 525922 543498 525978
rect 543554 525922 543622 525978
rect 543678 525922 561250 525978
rect 561306 525922 561374 525978
rect 561430 525922 561498 525978
rect 561554 525922 561622 525978
rect 561678 525922 579250 525978
rect 579306 525922 579374 525978
rect 579430 525922 579498 525978
rect 579554 525922 579622 525978
rect 579678 525922 596496 525978
rect 596552 525922 596620 525978
rect 596676 525922 596744 525978
rect 596800 525922 596868 525978
rect 596924 525922 597980 525978
rect -1916 525826 597980 525922
rect -1916 514350 597980 514446
rect -1916 514294 -1820 514350
rect -1764 514294 -1696 514350
rect -1640 514294 -1572 514350
rect -1516 514294 -1448 514350
rect -1392 514294 6970 514350
rect 7026 514294 7094 514350
rect 7150 514294 7218 514350
rect 7274 514294 7342 514350
rect 7398 514294 24970 514350
rect 25026 514294 25094 514350
rect 25150 514294 25218 514350
rect 25274 514294 25342 514350
rect 25398 514294 42970 514350
rect 43026 514294 43094 514350
rect 43150 514294 43218 514350
rect 43274 514294 43342 514350
rect 43398 514294 60970 514350
rect 61026 514294 61094 514350
rect 61150 514294 61218 514350
rect 61274 514294 61342 514350
rect 61398 514294 78970 514350
rect 79026 514294 79094 514350
rect 79150 514294 79218 514350
rect 79274 514294 79342 514350
rect 79398 514294 96970 514350
rect 97026 514294 97094 514350
rect 97150 514294 97218 514350
rect 97274 514294 97342 514350
rect 97398 514294 132970 514350
rect 133026 514294 133094 514350
rect 133150 514294 133218 514350
rect 133274 514294 133342 514350
rect 133398 514294 150970 514350
rect 151026 514294 151094 514350
rect 151150 514294 151218 514350
rect 151274 514294 151342 514350
rect 151398 514294 168970 514350
rect 169026 514294 169094 514350
rect 169150 514294 169218 514350
rect 169274 514294 169342 514350
rect 169398 514294 186970 514350
rect 187026 514294 187094 514350
rect 187150 514294 187218 514350
rect 187274 514294 187342 514350
rect 187398 514294 222970 514350
rect 223026 514294 223094 514350
rect 223150 514294 223218 514350
rect 223274 514294 223342 514350
rect 223398 514294 240970 514350
rect 241026 514294 241094 514350
rect 241150 514294 241218 514350
rect 241274 514294 241342 514350
rect 241398 514294 258970 514350
rect 259026 514294 259094 514350
rect 259150 514294 259218 514350
rect 259274 514294 259342 514350
rect 259398 514294 276970 514350
rect 277026 514294 277094 514350
rect 277150 514294 277218 514350
rect 277274 514294 277342 514350
rect 277398 514294 312970 514350
rect 313026 514294 313094 514350
rect 313150 514294 313218 514350
rect 313274 514294 313342 514350
rect 313398 514294 330970 514350
rect 331026 514294 331094 514350
rect 331150 514294 331218 514350
rect 331274 514294 331342 514350
rect 331398 514294 348970 514350
rect 349026 514294 349094 514350
rect 349150 514294 349218 514350
rect 349274 514294 349342 514350
rect 349398 514294 366970 514350
rect 367026 514294 367094 514350
rect 367150 514294 367218 514350
rect 367274 514294 367342 514350
rect 367398 514294 402970 514350
rect 403026 514294 403094 514350
rect 403150 514294 403218 514350
rect 403274 514294 403342 514350
rect 403398 514294 420970 514350
rect 421026 514294 421094 514350
rect 421150 514294 421218 514350
rect 421274 514294 421342 514350
rect 421398 514294 438970 514350
rect 439026 514294 439094 514350
rect 439150 514294 439218 514350
rect 439274 514294 439342 514350
rect 439398 514294 456970 514350
rect 457026 514294 457094 514350
rect 457150 514294 457218 514350
rect 457274 514294 457342 514350
rect 457398 514294 492970 514350
rect 493026 514294 493094 514350
rect 493150 514294 493218 514350
rect 493274 514294 493342 514350
rect 493398 514294 510970 514350
rect 511026 514294 511094 514350
rect 511150 514294 511218 514350
rect 511274 514294 511342 514350
rect 511398 514294 528970 514350
rect 529026 514294 529094 514350
rect 529150 514294 529218 514350
rect 529274 514294 529342 514350
rect 529398 514294 546970 514350
rect 547026 514294 547094 514350
rect 547150 514294 547218 514350
rect 547274 514294 547342 514350
rect 547398 514294 564970 514350
rect 565026 514294 565094 514350
rect 565150 514294 565218 514350
rect 565274 514294 565342 514350
rect 565398 514294 582970 514350
rect 583026 514294 583094 514350
rect 583150 514294 583218 514350
rect 583274 514294 583342 514350
rect 583398 514294 597456 514350
rect 597512 514294 597580 514350
rect 597636 514294 597704 514350
rect 597760 514294 597828 514350
rect 597884 514294 597980 514350
rect -1916 514226 597980 514294
rect -1916 514170 -1820 514226
rect -1764 514170 -1696 514226
rect -1640 514170 -1572 514226
rect -1516 514170 -1448 514226
rect -1392 514170 6970 514226
rect 7026 514170 7094 514226
rect 7150 514170 7218 514226
rect 7274 514170 7342 514226
rect 7398 514170 24970 514226
rect 25026 514170 25094 514226
rect 25150 514170 25218 514226
rect 25274 514170 25342 514226
rect 25398 514170 42970 514226
rect 43026 514170 43094 514226
rect 43150 514170 43218 514226
rect 43274 514170 43342 514226
rect 43398 514170 60970 514226
rect 61026 514170 61094 514226
rect 61150 514170 61218 514226
rect 61274 514170 61342 514226
rect 61398 514170 78970 514226
rect 79026 514170 79094 514226
rect 79150 514170 79218 514226
rect 79274 514170 79342 514226
rect 79398 514170 96970 514226
rect 97026 514170 97094 514226
rect 97150 514170 97218 514226
rect 97274 514170 97342 514226
rect 97398 514170 132970 514226
rect 133026 514170 133094 514226
rect 133150 514170 133218 514226
rect 133274 514170 133342 514226
rect 133398 514170 150970 514226
rect 151026 514170 151094 514226
rect 151150 514170 151218 514226
rect 151274 514170 151342 514226
rect 151398 514170 168970 514226
rect 169026 514170 169094 514226
rect 169150 514170 169218 514226
rect 169274 514170 169342 514226
rect 169398 514170 186970 514226
rect 187026 514170 187094 514226
rect 187150 514170 187218 514226
rect 187274 514170 187342 514226
rect 187398 514170 222970 514226
rect 223026 514170 223094 514226
rect 223150 514170 223218 514226
rect 223274 514170 223342 514226
rect 223398 514170 240970 514226
rect 241026 514170 241094 514226
rect 241150 514170 241218 514226
rect 241274 514170 241342 514226
rect 241398 514170 258970 514226
rect 259026 514170 259094 514226
rect 259150 514170 259218 514226
rect 259274 514170 259342 514226
rect 259398 514170 276970 514226
rect 277026 514170 277094 514226
rect 277150 514170 277218 514226
rect 277274 514170 277342 514226
rect 277398 514170 312970 514226
rect 313026 514170 313094 514226
rect 313150 514170 313218 514226
rect 313274 514170 313342 514226
rect 313398 514170 330970 514226
rect 331026 514170 331094 514226
rect 331150 514170 331218 514226
rect 331274 514170 331342 514226
rect 331398 514170 348970 514226
rect 349026 514170 349094 514226
rect 349150 514170 349218 514226
rect 349274 514170 349342 514226
rect 349398 514170 366970 514226
rect 367026 514170 367094 514226
rect 367150 514170 367218 514226
rect 367274 514170 367342 514226
rect 367398 514170 402970 514226
rect 403026 514170 403094 514226
rect 403150 514170 403218 514226
rect 403274 514170 403342 514226
rect 403398 514170 420970 514226
rect 421026 514170 421094 514226
rect 421150 514170 421218 514226
rect 421274 514170 421342 514226
rect 421398 514170 438970 514226
rect 439026 514170 439094 514226
rect 439150 514170 439218 514226
rect 439274 514170 439342 514226
rect 439398 514170 456970 514226
rect 457026 514170 457094 514226
rect 457150 514170 457218 514226
rect 457274 514170 457342 514226
rect 457398 514170 492970 514226
rect 493026 514170 493094 514226
rect 493150 514170 493218 514226
rect 493274 514170 493342 514226
rect 493398 514170 510970 514226
rect 511026 514170 511094 514226
rect 511150 514170 511218 514226
rect 511274 514170 511342 514226
rect 511398 514170 528970 514226
rect 529026 514170 529094 514226
rect 529150 514170 529218 514226
rect 529274 514170 529342 514226
rect 529398 514170 546970 514226
rect 547026 514170 547094 514226
rect 547150 514170 547218 514226
rect 547274 514170 547342 514226
rect 547398 514170 564970 514226
rect 565026 514170 565094 514226
rect 565150 514170 565218 514226
rect 565274 514170 565342 514226
rect 565398 514170 582970 514226
rect 583026 514170 583094 514226
rect 583150 514170 583218 514226
rect 583274 514170 583342 514226
rect 583398 514170 597456 514226
rect 597512 514170 597580 514226
rect 597636 514170 597704 514226
rect 597760 514170 597828 514226
rect 597884 514170 597980 514226
rect -1916 514102 597980 514170
rect -1916 514046 -1820 514102
rect -1764 514046 -1696 514102
rect -1640 514046 -1572 514102
rect -1516 514046 -1448 514102
rect -1392 514046 6970 514102
rect 7026 514046 7094 514102
rect 7150 514046 7218 514102
rect 7274 514046 7342 514102
rect 7398 514046 24970 514102
rect 25026 514046 25094 514102
rect 25150 514046 25218 514102
rect 25274 514046 25342 514102
rect 25398 514046 42970 514102
rect 43026 514046 43094 514102
rect 43150 514046 43218 514102
rect 43274 514046 43342 514102
rect 43398 514046 60970 514102
rect 61026 514046 61094 514102
rect 61150 514046 61218 514102
rect 61274 514046 61342 514102
rect 61398 514046 78970 514102
rect 79026 514046 79094 514102
rect 79150 514046 79218 514102
rect 79274 514046 79342 514102
rect 79398 514046 96970 514102
rect 97026 514046 97094 514102
rect 97150 514046 97218 514102
rect 97274 514046 97342 514102
rect 97398 514046 132970 514102
rect 133026 514046 133094 514102
rect 133150 514046 133218 514102
rect 133274 514046 133342 514102
rect 133398 514046 150970 514102
rect 151026 514046 151094 514102
rect 151150 514046 151218 514102
rect 151274 514046 151342 514102
rect 151398 514046 168970 514102
rect 169026 514046 169094 514102
rect 169150 514046 169218 514102
rect 169274 514046 169342 514102
rect 169398 514046 186970 514102
rect 187026 514046 187094 514102
rect 187150 514046 187218 514102
rect 187274 514046 187342 514102
rect 187398 514046 222970 514102
rect 223026 514046 223094 514102
rect 223150 514046 223218 514102
rect 223274 514046 223342 514102
rect 223398 514046 240970 514102
rect 241026 514046 241094 514102
rect 241150 514046 241218 514102
rect 241274 514046 241342 514102
rect 241398 514046 258970 514102
rect 259026 514046 259094 514102
rect 259150 514046 259218 514102
rect 259274 514046 259342 514102
rect 259398 514046 276970 514102
rect 277026 514046 277094 514102
rect 277150 514046 277218 514102
rect 277274 514046 277342 514102
rect 277398 514046 312970 514102
rect 313026 514046 313094 514102
rect 313150 514046 313218 514102
rect 313274 514046 313342 514102
rect 313398 514046 330970 514102
rect 331026 514046 331094 514102
rect 331150 514046 331218 514102
rect 331274 514046 331342 514102
rect 331398 514046 348970 514102
rect 349026 514046 349094 514102
rect 349150 514046 349218 514102
rect 349274 514046 349342 514102
rect 349398 514046 366970 514102
rect 367026 514046 367094 514102
rect 367150 514046 367218 514102
rect 367274 514046 367342 514102
rect 367398 514046 402970 514102
rect 403026 514046 403094 514102
rect 403150 514046 403218 514102
rect 403274 514046 403342 514102
rect 403398 514046 420970 514102
rect 421026 514046 421094 514102
rect 421150 514046 421218 514102
rect 421274 514046 421342 514102
rect 421398 514046 438970 514102
rect 439026 514046 439094 514102
rect 439150 514046 439218 514102
rect 439274 514046 439342 514102
rect 439398 514046 456970 514102
rect 457026 514046 457094 514102
rect 457150 514046 457218 514102
rect 457274 514046 457342 514102
rect 457398 514046 492970 514102
rect 493026 514046 493094 514102
rect 493150 514046 493218 514102
rect 493274 514046 493342 514102
rect 493398 514046 510970 514102
rect 511026 514046 511094 514102
rect 511150 514046 511218 514102
rect 511274 514046 511342 514102
rect 511398 514046 528970 514102
rect 529026 514046 529094 514102
rect 529150 514046 529218 514102
rect 529274 514046 529342 514102
rect 529398 514046 546970 514102
rect 547026 514046 547094 514102
rect 547150 514046 547218 514102
rect 547274 514046 547342 514102
rect 547398 514046 564970 514102
rect 565026 514046 565094 514102
rect 565150 514046 565218 514102
rect 565274 514046 565342 514102
rect 565398 514046 582970 514102
rect 583026 514046 583094 514102
rect 583150 514046 583218 514102
rect 583274 514046 583342 514102
rect 583398 514046 597456 514102
rect 597512 514046 597580 514102
rect 597636 514046 597704 514102
rect 597760 514046 597828 514102
rect 597884 514046 597980 514102
rect -1916 513978 597980 514046
rect -1916 513922 -1820 513978
rect -1764 513922 -1696 513978
rect -1640 513922 -1572 513978
rect -1516 513922 -1448 513978
rect -1392 513922 6970 513978
rect 7026 513922 7094 513978
rect 7150 513922 7218 513978
rect 7274 513922 7342 513978
rect 7398 513922 24970 513978
rect 25026 513922 25094 513978
rect 25150 513922 25218 513978
rect 25274 513922 25342 513978
rect 25398 513922 42970 513978
rect 43026 513922 43094 513978
rect 43150 513922 43218 513978
rect 43274 513922 43342 513978
rect 43398 513922 60970 513978
rect 61026 513922 61094 513978
rect 61150 513922 61218 513978
rect 61274 513922 61342 513978
rect 61398 513922 78970 513978
rect 79026 513922 79094 513978
rect 79150 513922 79218 513978
rect 79274 513922 79342 513978
rect 79398 513922 96970 513978
rect 97026 513922 97094 513978
rect 97150 513922 97218 513978
rect 97274 513922 97342 513978
rect 97398 513922 132970 513978
rect 133026 513922 133094 513978
rect 133150 513922 133218 513978
rect 133274 513922 133342 513978
rect 133398 513922 150970 513978
rect 151026 513922 151094 513978
rect 151150 513922 151218 513978
rect 151274 513922 151342 513978
rect 151398 513922 168970 513978
rect 169026 513922 169094 513978
rect 169150 513922 169218 513978
rect 169274 513922 169342 513978
rect 169398 513922 186970 513978
rect 187026 513922 187094 513978
rect 187150 513922 187218 513978
rect 187274 513922 187342 513978
rect 187398 513922 222970 513978
rect 223026 513922 223094 513978
rect 223150 513922 223218 513978
rect 223274 513922 223342 513978
rect 223398 513922 240970 513978
rect 241026 513922 241094 513978
rect 241150 513922 241218 513978
rect 241274 513922 241342 513978
rect 241398 513922 258970 513978
rect 259026 513922 259094 513978
rect 259150 513922 259218 513978
rect 259274 513922 259342 513978
rect 259398 513922 276970 513978
rect 277026 513922 277094 513978
rect 277150 513922 277218 513978
rect 277274 513922 277342 513978
rect 277398 513922 312970 513978
rect 313026 513922 313094 513978
rect 313150 513922 313218 513978
rect 313274 513922 313342 513978
rect 313398 513922 330970 513978
rect 331026 513922 331094 513978
rect 331150 513922 331218 513978
rect 331274 513922 331342 513978
rect 331398 513922 348970 513978
rect 349026 513922 349094 513978
rect 349150 513922 349218 513978
rect 349274 513922 349342 513978
rect 349398 513922 366970 513978
rect 367026 513922 367094 513978
rect 367150 513922 367218 513978
rect 367274 513922 367342 513978
rect 367398 513922 402970 513978
rect 403026 513922 403094 513978
rect 403150 513922 403218 513978
rect 403274 513922 403342 513978
rect 403398 513922 420970 513978
rect 421026 513922 421094 513978
rect 421150 513922 421218 513978
rect 421274 513922 421342 513978
rect 421398 513922 438970 513978
rect 439026 513922 439094 513978
rect 439150 513922 439218 513978
rect 439274 513922 439342 513978
rect 439398 513922 456970 513978
rect 457026 513922 457094 513978
rect 457150 513922 457218 513978
rect 457274 513922 457342 513978
rect 457398 513922 492970 513978
rect 493026 513922 493094 513978
rect 493150 513922 493218 513978
rect 493274 513922 493342 513978
rect 493398 513922 510970 513978
rect 511026 513922 511094 513978
rect 511150 513922 511218 513978
rect 511274 513922 511342 513978
rect 511398 513922 528970 513978
rect 529026 513922 529094 513978
rect 529150 513922 529218 513978
rect 529274 513922 529342 513978
rect 529398 513922 546970 513978
rect 547026 513922 547094 513978
rect 547150 513922 547218 513978
rect 547274 513922 547342 513978
rect 547398 513922 564970 513978
rect 565026 513922 565094 513978
rect 565150 513922 565218 513978
rect 565274 513922 565342 513978
rect 565398 513922 582970 513978
rect 583026 513922 583094 513978
rect 583150 513922 583218 513978
rect 583274 513922 583342 513978
rect 583398 513922 597456 513978
rect 597512 513922 597580 513978
rect 597636 513922 597704 513978
rect 597760 513922 597828 513978
rect 597884 513922 597980 513978
rect -1916 513826 597980 513922
rect -1916 508350 597980 508446
rect -1916 508294 -860 508350
rect -804 508294 -736 508350
rect -680 508294 -612 508350
rect -556 508294 -488 508350
rect -432 508294 3250 508350
rect 3306 508294 3374 508350
rect 3430 508294 3498 508350
rect 3554 508294 3622 508350
rect 3678 508294 21250 508350
rect 21306 508294 21374 508350
rect 21430 508294 21498 508350
rect 21554 508294 21622 508350
rect 21678 508294 39250 508350
rect 39306 508294 39374 508350
rect 39430 508294 39498 508350
rect 39554 508294 39622 508350
rect 39678 508294 57250 508350
rect 57306 508294 57374 508350
rect 57430 508294 57498 508350
rect 57554 508294 57622 508350
rect 57678 508294 93250 508350
rect 93306 508294 93374 508350
rect 93430 508294 93498 508350
rect 93554 508294 93622 508350
rect 93678 508294 111250 508350
rect 111306 508294 111374 508350
rect 111430 508294 111498 508350
rect 111554 508294 111622 508350
rect 111678 508294 129250 508350
rect 129306 508294 129374 508350
rect 129430 508294 129498 508350
rect 129554 508294 129622 508350
rect 129678 508294 147250 508350
rect 147306 508294 147374 508350
rect 147430 508294 147498 508350
rect 147554 508294 147622 508350
rect 147678 508294 183250 508350
rect 183306 508294 183374 508350
rect 183430 508294 183498 508350
rect 183554 508294 183622 508350
rect 183678 508294 201250 508350
rect 201306 508294 201374 508350
rect 201430 508294 201498 508350
rect 201554 508294 201622 508350
rect 201678 508294 219250 508350
rect 219306 508294 219374 508350
rect 219430 508294 219498 508350
rect 219554 508294 219622 508350
rect 219678 508294 237250 508350
rect 237306 508294 237374 508350
rect 237430 508294 237498 508350
rect 237554 508294 237622 508350
rect 237678 508294 273250 508350
rect 273306 508294 273374 508350
rect 273430 508294 273498 508350
rect 273554 508294 273622 508350
rect 273678 508294 291250 508350
rect 291306 508294 291374 508350
rect 291430 508294 291498 508350
rect 291554 508294 291622 508350
rect 291678 508294 309250 508350
rect 309306 508294 309374 508350
rect 309430 508294 309498 508350
rect 309554 508294 309622 508350
rect 309678 508294 327250 508350
rect 327306 508294 327374 508350
rect 327430 508294 327498 508350
rect 327554 508294 327622 508350
rect 327678 508294 363250 508350
rect 363306 508294 363374 508350
rect 363430 508294 363498 508350
rect 363554 508294 363622 508350
rect 363678 508294 381250 508350
rect 381306 508294 381374 508350
rect 381430 508294 381498 508350
rect 381554 508294 381622 508350
rect 381678 508294 399250 508350
rect 399306 508294 399374 508350
rect 399430 508294 399498 508350
rect 399554 508294 399622 508350
rect 399678 508294 417250 508350
rect 417306 508294 417374 508350
rect 417430 508294 417498 508350
rect 417554 508294 417622 508350
rect 417678 508294 453250 508350
rect 453306 508294 453374 508350
rect 453430 508294 453498 508350
rect 453554 508294 453622 508350
rect 453678 508294 471250 508350
rect 471306 508294 471374 508350
rect 471430 508294 471498 508350
rect 471554 508294 471622 508350
rect 471678 508294 489250 508350
rect 489306 508294 489374 508350
rect 489430 508294 489498 508350
rect 489554 508294 489622 508350
rect 489678 508294 507250 508350
rect 507306 508294 507374 508350
rect 507430 508294 507498 508350
rect 507554 508294 507622 508350
rect 507678 508294 543250 508350
rect 543306 508294 543374 508350
rect 543430 508294 543498 508350
rect 543554 508294 543622 508350
rect 543678 508294 561250 508350
rect 561306 508294 561374 508350
rect 561430 508294 561498 508350
rect 561554 508294 561622 508350
rect 561678 508294 579250 508350
rect 579306 508294 579374 508350
rect 579430 508294 579498 508350
rect 579554 508294 579622 508350
rect 579678 508294 596496 508350
rect 596552 508294 596620 508350
rect 596676 508294 596744 508350
rect 596800 508294 596868 508350
rect 596924 508294 597980 508350
rect -1916 508226 597980 508294
rect -1916 508170 -860 508226
rect -804 508170 -736 508226
rect -680 508170 -612 508226
rect -556 508170 -488 508226
rect -432 508170 3250 508226
rect 3306 508170 3374 508226
rect 3430 508170 3498 508226
rect 3554 508170 3622 508226
rect 3678 508170 21250 508226
rect 21306 508170 21374 508226
rect 21430 508170 21498 508226
rect 21554 508170 21622 508226
rect 21678 508170 39250 508226
rect 39306 508170 39374 508226
rect 39430 508170 39498 508226
rect 39554 508170 39622 508226
rect 39678 508170 57250 508226
rect 57306 508170 57374 508226
rect 57430 508170 57498 508226
rect 57554 508170 57622 508226
rect 57678 508170 93250 508226
rect 93306 508170 93374 508226
rect 93430 508170 93498 508226
rect 93554 508170 93622 508226
rect 93678 508170 111250 508226
rect 111306 508170 111374 508226
rect 111430 508170 111498 508226
rect 111554 508170 111622 508226
rect 111678 508170 129250 508226
rect 129306 508170 129374 508226
rect 129430 508170 129498 508226
rect 129554 508170 129622 508226
rect 129678 508170 147250 508226
rect 147306 508170 147374 508226
rect 147430 508170 147498 508226
rect 147554 508170 147622 508226
rect 147678 508170 183250 508226
rect 183306 508170 183374 508226
rect 183430 508170 183498 508226
rect 183554 508170 183622 508226
rect 183678 508170 201250 508226
rect 201306 508170 201374 508226
rect 201430 508170 201498 508226
rect 201554 508170 201622 508226
rect 201678 508170 219250 508226
rect 219306 508170 219374 508226
rect 219430 508170 219498 508226
rect 219554 508170 219622 508226
rect 219678 508170 237250 508226
rect 237306 508170 237374 508226
rect 237430 508170 237498 508226
rect 237554 508170 237622 508226
rect 237678 508170 273250 508226
rect 273306 508170 273374 508226
rect 273430 508170 273498 508226
rect 273554 508170 273622 508226
rect 273678 508170 291250 508226
rect 291306 508170 291374 508226
rect 291430 508170 291498 508226
rect 291554 508170 291622 508226
rect 291678 508170 309250 508226
rect 309306 508170 309374 508226
rect 309430 508170 309498 508226
rect 309554 508170 309622 508226
rect 309678 508170 327250 508226
rect 327306 508170 327374 508226
rect 327430 508170 327498 508226
rect 327554 508170 327622 508226
rect 327678 508170 363250 508226
rect 363306 508170 363374 508226
rect 363430 508170 363498 508226
rect 363554 508170 363622 508226
rect 363678 508170 381250 508226
rect 381306 508170 381374 508226
rect 381430 508170 381498 508226
rect 381554 508170 381622 508226
rect 381678 508170 399250 508226
rect 399306 508170 399374 508226
rect 399430 508170 399498 508226
rect 399554 508170 399622 508226
rect 399678 508170 417250 508226
rect 417306 508170 417374 508226
rect 417430 508170 417498 508226
rect 417554 508170 417622 508226
rect 417678 508170 453250 508226
rect 453306 508170 453374 508226
rect 453430 508170 453498 508226
rect 453554 508170 453622 508226
rect 453678 508170 471250 508226
rect 471306 508170 471374 508226
rect 471430 508170 471498 508226
rect 471554 508170 471622 508226
rect 471678 508170 489250 508226
rect 489306 508170 489374 508226
rect 489430 508170 489498 508226
rect 489554 508170 489622 508226
rect 489678 508170 507250 508226
rect 507306 508170 507374 508226
rect 507430 508170 507498 508226
rect 507554 508170 507622 508226
rect 507678 508170 543250 508226
rect 543306 508170 543374 508226
rect 543430 508170 543498 508226
rect 543554 508170 543622 508226
rect 543678 508170 561250 508226
rect 561306 508170 561374 508226
rect 561430 508170 561498 508226
rect 561554 508170 561622 508226
rect 561678 508170 579250 508226
rect 579306 508170 579374 508226
rect 579430 508170 579498 508226
rect 579554 508170 579622 508226
rect 579678 508170 596496 508226
rect 596552 508170 596620 508226
rect 596676 508170 596744 508226
rect 596800 508170 596868 508226
rect 596924 508170 597980 508226
rect -1916 508102 597980 508170
rect -1916 508046 -860 508102
rect -804 508046 -736 508102
rect -680 508046 -612 508102
rect -556 508046 -488 508102
rect -432 508046 3250 508102
rect 3306 508046 3374 508102
rect 3430 508046 3498 508102
rect 3554 508046 3622 508102
rect 3678 508046 21250 508102
rect 21306 508046 21374 508102
rect 21430 508046 21498 508102
rect 21554 508046 21622 508102
rect 21678 508046 39250 508102
rect 39306 508046 39374 508102
rect 39430 508046 39498 508102
rect 39554 508046 39622 508102
rect 39678 508046 57250 508102
rect 57306 508046 57374 508102
rect 57430 508046 57498 508102
rect 57554 508046 57622 508102
rect 57678 508046 93250 508102
rect 93306 508046 93374 508102
rect 93430 508046 93498 508102
rect 93554 508046 93622 508102
rect 93678 508046 111250 508102
rect 111306 508046 111374 508102
rect 111430 508046 111498 508102
rect 111554 508046 111622 508102
rect 111678 508046 129250 508102
rect 129306 508046 129374 508102
rect 129430 508046 129498 508102
rect 129554 508046 129622 508102
rect 129678 508046 147250 508102
rect 147306 508046 147374 508102
rect 147430 508046 147498 508102
rect 147554 508046 147622 508102
rect 147678 508046 183250 508102
rect 183306 508046 183374 508102
rect 183430 508046 183498 508102
rect 183554 508046 183622 508102
rect 183678 508046 201250 508102
rect 201306 508046 201374 508102
rect 201430 508046 201498 508102
rect 201554 508046 201622 508102
rect 201678 508046 219250 508102
rect 219306 508046 219374 508102
rect 219430 508046 219498 508102
rect 219554 508046 219622 508102
rect 219678 508046 237250 508102
rect 237306 508046 237374 508102
rect 237430 508046 237498 508102
rect 237554 508046 237622 508102
rect 237678 508046 273250 508102
rect 273306 508046 273374 508102
rect 273430 508046 273498 508102
rect 273554 508046 273622 508102
rect 273678 508046 291250 508102
rect 291306 508046 291374 508102
rect 291430 508046 291498 508102
rect 291554 508046 291622 508102
rect 291678 508046 309250 508102
rect 309306 508046 309374 508102
rect 309430 508046 309498 508102
rect 309554 508046 309622 508102
rect 309678 508046 327250 508102
rect 327306 508046 327374 508102
rect 327430 508046 327498 508102
rect 327554 508046 327622 508102
rect 327678 508046 363250 508102
rect 363306 508046 363374 508102
rect 363430 508046 363498 508102
rect 363554 508046 363622 508102
rect 363678 508046 381250 508102
rect 381306 508046 381374 508102
rect 381430 508046 381498 508102
rect 381554 508046 381622 508102
rect 381678 508046 399250 508102
rect 399306 508046 399374 508102
rect 399430 508046 399498 508102
rect 399554 508046 399622 508102
rect 399678 508046 417250 508102
rect 417306 508046 417374 508102
rect 417430 508046 417498 508102
rect 417554 508046 417622 508102
rect 417678 508046 453250 508102
rect 453306 508046 453374 508102
rect 453430 508046 453498 508102
rect 453554 508046 453622 508102
rect 453678 508046 471250 508102
rect 471306 508046 471374 508102
rect 471430 508046 471498 508102
rect 471554 508046 471622 508102
rect 471678 508046 489250 508102
rect 489306 508046 489374 508102
rect 489430 508046 489498 508102
rect 489554 508046 489622 508102
rect 489678 508046 507250 508102
rect 507306 508046 507374 508102
rect 507430 508046 507498 508102
rect 507554 508046 507622 508102
rect 507678 508046 543250 508102
rect 543306 508046 543374 508102
rect 543430 508046 543498 508102
rect 543554 508046 543622 508102
rect 543678 508046 561250 508102
rect 561306 508046 561374 508102
rect 561430 508046 561498 508102
rect 561554 508046 561622 508102
rect 561678 508046 579250 508102
rect 579306 508046 579374 508102
rect 579430 508046 579498 508102
rect 579554 508046 579622 508102
rect 579678 508046 596496 508102
rect 596552 508046 596620 508102
rect 596676 508046 596744 508102
rect 596800 508046 596868 508102
rect 596924 508046 597980 508102
rect -1916 507978 597980 508046
rect -1916 507922 -860 507978
rect -804 507922 -736 507978
rect -680 507922 -612 507978
rect -556 507922 -488 507978
rect -432 507922 3250 507978
rect 3306 507922 3374 507978
rect 3430 507922 3498 507978
rect 3554 507922 3622 507978
rect 3678 507922 21250 507978
rect 21306 507922 21374 507978
rect 21430 507922 21498 507978
rect 21554 507922 21622 507978
rect 21678 507922 39250 507978
rect 39306 507922 39374 507978
rect 39430 507922 39498 507978
rect 39554 507922 39622 507978
rect 39678 507922 57250 507978
rect 57306 507922 57374 507978
rect 57430 507922 57498 507978
rect 57554 507922 57622 507978
rect 57678 507922 93250 507978
rect 93306 507922 93374 507978
rect 93430 507922 93498 507978
rect 93554 507922 93622 507978
rect 93678 507922 111250 507978
rect 111306 507922 111374 507978
rect 111430 507922 111498 507978
rect 111554 507922 111622 507978
rect 111678 507922 129250 507978
rect 129306 507922 129374 507978
rect 129430 507922 129498 507978
rect 129554 507922 129622 507978
rect 129678 507922 147250 507978
rect 147306 507922 147374 507978
rect 147430 507922 147498 507978
rect 147554 507922 147622 507978
rect 147678 507922 183250 507978
rect 183306 507922 183374 507978
rect 183430 507922 183498 507978
rect 183554 507922 183622 507978
rect 183678 507922 201250 507978
rect 201306 507922 201374 507978
rect 201430 507922 201498 507978
rect 201554 507922 201622 507978
rect 201678 507922 219250 507978
rect 219306 507922 219374 507978
rect 219430 507922 219498 507978
rect 219554 507922 219622 507978
rect 219678 507922 237250 507978
rect 237306 507922 237374 507978
rect 237430 507922 237498 507978
rect 237554 507922 237622 507978
rect 237678 507922 273250 507978
rect 273306 507922 273374 507978
rect 273430 507922 273498 507978
rect 273554 507922 273622 507978
rect 273678 507922 291250 507978
rect 291306 507922 291374 507978
rect 291430 507922 291498 507978
rect 291554 507922 291622 507978
rect 291678 507922 309250 507978
rect 309306 507922 309374 507978
rect 309430 507922 309498 507978
rect 309554 507922 309622 507978
rect 309678 507922 327250 507978
rect 327306 507922 327374 507978
rect 327430 507922 327498 507978
rect 327554 507922 327622 507978
rect 327678 507922 363250 507978
rect 363306 507922 363374 507978
rect 363430 507922 363498 507978
rect 363554 507922 363622 507978
rect 363678 507922 381250 507978
rect 381306 507922 381374 507978
rect 381430 507922 381498 507978
rect 381554 507922 381622 507978
rect 381678 507922 399250 507978
rect 399306 507922 399374 507978
rect 399430 507922 399498 507978
rect 399554 507922 399622 507978
rect 399678 507922 417250 507978
rect 417306 507922 417374 507978
rect 417430 507922 417498 507978
rect 417554 507922 417622 507978
rect 417678 507922 453250 507978
rect 453306 507922 453374 507978
rect 453430 507922 453498 507978
rect 453554 507922 453622 507978
rect 453678 507922 471250 507978
rect 471306 507922 471374 507978
rect 471430 507922 471498 507978
rect 471554 507922 471622 507978
rect 471678 507922 489250 507978
rect 489306 507922 489374 507978
rect 489430 507922 489498 507978
rect 489554 507922 489622 507978
rect 489678 507922 507250 507978
rect 507306 507922 507374 507978
rect 507430 507922 507498 507978
rect 507554 507922 507622 507978
rect 507678 507922 543250 507978
rect 543306 507922 543374 507978
rect 543430 507922 543498 507978
rect 543554 507922 543622 507978
rect 543678 507922 561250 507978
rect 561306 507922 561374 507978
rect 561430 507922 561498 507978
rect 561554 507922 561622 507978
rect 561678 507922 579250 507978
rect 579306 507922 579374 507978
rect 579430 507922 579498 507978
rect 579554 507922 579622 507978
rect 579678 507922 596496 507978
rect 596552 507922 596620 507978
rect 596676 507922 596744 507978
rect 596800 507922 596868 507978
rect 596924 507922 597980 507978
rect -1916 507826 597980 507922
rect -1916 496350 597980 496446
rect -1916 496294 -1820 496350
rect -1764 496294 -1696 496350
rect -1640 496294 -1572 496350
rect -1516 496294 -1448 496350
rect -1392 496294 6970 496350
rect 7026 496294 7094 496350
rect 7150 496294 7218 496350
rect 7274 496294 7342 496350
rect 7398 496294 24970 496350
rect 25026 496294 25094 496350
rect 25150 496294 25218 496350
rect 25274 496294 25342 496350
rect 25398 496294 42970 496350
rect 43026 496294 43094 496350
rect 43150 496294 43218 496350
rect 43274 496294 43342 496350
rect 43398 496294 60970 496350
rect 61026 496294 61094 496350
rect 61150 496294 61218 496350
rect 61274 496294 61342 496350
rect 61398 496294 78970 496350
rect 79026 496294 79094 496350
rect 79150 496294 79218 496350
rect 79274 496294 79342 496350
rect 79398 496294 96970 496350
rect 97026 496294 97094 496350
rect 97150 496294 97218 496350
rect 97274 496294 97342 496350
rect 97398 496294 132970 496350
rect 133026 496294 133094 496350
rect 133150 496294 133218 496350
rect 133274 496294 133342 496350
rect 133398 496294 150970 496350
rect 151026 496294 151094 496350
rect 151150 496294 151218 496350
rect 151274 496294 151342 496350
rect 151398 496294 168970 496350
rect 169026 496294 169094 496350
rect 169150 496294 169218 496350
rect 169274 496294 169342 496350
rect 169398 496294 186970 496350
rect 187026 496294 187094 496350
rect 187150 496294 187218 496350
rect 187274 496294 187342 496350
rect 187398 496294 222970 496350
rect 223026 496294 223094 496350
rect 223150 496294 223218 496350
rect 223274 496294 223342 496350
rect 223398 496294 240970 496350
rect 241026 496294 241094 496350
rect 241150 496294 241218 496350
rect 241274 496294 241342 496350
rect 241398 496294 258970 496350
rect 259026 496294 259094 496350
rect 259150 496294 259218 496350
rect 259274 496294 259342 496350
rect 259398 496294 276970 496350
rect 277026 496294 277094 496350
rect 277150 496294 277218 496350
rect 277274 496294 277342 496350
rect 277398 496294 312970 496350
rect 313026 496294 313094 496350
rect 313150 496294 313218 496350
rect 313274 496294 313342 496350
rect 313398 496294 330970 496350
rect 331026 496294 331094 496350
rect 331150 496294 331218 496350
rect 331274 496294 331342 496350
rect 331398 496294 348970 496350
rect 349026 496294 349094 496350
rect 349150 496294 349218 496350
rect 349274 496294 349342 496350
rect 349398 496294 366970 496350
rect 367026 496294 367094 496350
rect 367150 496294 367218 496350
rect 367274 496294 367342 496350
rect 367398 496294 402970 496350
rect 403026 496294 403094 496350
rect 403150 496294 403218 496350
rect 403274 496294 403342 496350
rect 403398 496294 420970 496350
rect 421026 496294 421094 496350
rect 421150 496294 421218 496350
rect 421274 496294 421342 496350
rect 421398 496294 438970 496350
rect 439026 496294 439094 496350
rect 439150 496294 439218 496350
rect 439274 496294 439342 496350
rect 439398 496294 456970 496350
rect 457026 496294 457094 496350
rect 457150 496294 457218 496350
rect 457274 496294 457342 496350
rect 457398 496294 492970 496350
rect 493026 496294 493094 496350
rect 493150 496294 493218 496350
rect 493274 496294 493342 496350
rect 493398 496294 510970 496350
rect 511026 496294 511094 496350
rect 511150 496294 511218 496350
rect 511274 496294 511342 496350
rect 511398 496294 528970 496350
rect 529026 496294 529094 496350
rect 529150 496294 529218 496350
rect 529274 496294 529342 496350
rect 529398 496294 546970 496350
rect 547026 496294 547094 496350
rect 547150 496294 547218 496350
rect 547274 496294 547342 496350
rect 547398 496294 568058 496350
rect 568114 496294 568182 496350
rect 568238 496294 574862 496350
rect 574918 496294 574986 496350
rect 575042 496294 581666 496350
rect 581722 496294 581790 496350
rect 581846 496294 582970 496350
rect 583026 496294 583094 496350
rect 583150 496294 583218 496350
rect 583274 496294 583342 496350
rect 583398 496294 588470 496350
rect 588526 496294 588594 496350
rect 588650 496294 597456 496350
rect 597512 496294 597580 496350
rect 597636 496294 597704 496350
rect 597760 496294 597828 496350
rect 597884 496294 597980 496350
rect -1916 496226 597980 496294
rect -1916 496170 -1820 496226
rect -1764 496170 -1696 496226
rect -1640 496170 -1572 496226
rect -1516 496170 -1448 496226
rect -1392 496170 6970 496226
rect 7026 496170 7094 496226
rect 7150 496170 7218 496226
rect 7274 496170 7342 496226
rect 7398 496170 24970 496226
rect 25026 496170 25094 496226
rect 25150 496170 25218 496226
rect 25274 496170 25342 496226
rect 25398 496170 42970 496226
rect 43026 496170 43094 496226
rect 43150 496170 43218 496226
rect 43274 496170 43342 496226
rect 43398 496170 60970 496226
rect 61026 496170 61094 496226
rect 61150 496170 61218 496226
rect 61274 496170 61342 496226
rect 61398 496170 78970 496226
rect 79026 496170 79094 496226
rect 79150 496170 79218 496226
rect 79274 496170 79342 496226
rect 79398 496170 96970 496226
rect 97026 496170 97094 496226
rect 97150 496170 97218 496226
rect 97274 496170 97342 496226
rect 97398 496170 132970 496226
rect 133026 496170 133094 496226
rect 133150 496170 133218 496226
rect 133274 496170 133342 496226
rect 133398 496170 150970 496226
rect 151026 496170 151094 496226
rect 151150 496170 151218 496226
rect 151274 496170 151342 496226
rect 151398 496170 168970 496226
rect 169026 496170 169094 496226
rect 169150 496170 169218 496226
rect 169274 496170 169342 496226
rect 169398 496170 186970 496226
rect 187026 496170 187094 496226
rect 187150 496170 187218 496226
rect 187274 496170 187342 496226
rect 187398 496170 222970 496226
rect 223026 496170 223094 496226
rect 223150 496170 223218 496226
rect 223274 496170 223342 496226
rect 223398 496170 240970 496226
rect 241026 496170 241094 496226
rect 241150 496170 241218 496226
rect 241274 496170 241342 496226
rect 241398 496170 258970 496226
rect 259026 496170 259094 496226
rect 259150 496170 259218 496226
rect 259274 496170 259342 496226
rect 259398 496170 276970 496226
rect 277026 496170 277094 496226
rect 277150 496170 277218 496226
rect 277274 496170 277342 496226
rect 277398 496170 312970 496226
rect 313026 496170 313094 496226
rect 313150 496170 313218 496226
rect 313274 496170 313342 496226
rect 313398 496170 330970 496226
rect 331026 496170 331094 496226
rect 331150 496170 331218 496226
rect 331274 496170 331342 496226
rect 331398 496170 348970 496226
rect 349026 496170 349094 496226
rect 349150 496170 349218 496226
rect 349274 496170 349342 496226
rect 349398 496170 366970 496226
rect 367026 496170 367094 496226
rect 367150 496170 367218 496226
rect 367274 496170 367342 496226
rect 367398 496170 402970 496226
rect 403026 496170 403094 496226
rect 403150 496170 403218 496226
rect 403274 496170 403342 496226
rect 403398 496170 420970 496226
rect 421026 496170 421094 496226
rect 421150 496170 421218 496226
rect 421274 496170 421342 496226
rect 421398 496170 438970 496226
rect 439026 496170 439094 496226
rect 439150 496170 439218 496226
rect 439274 496170 439342 496226
rect 439398 496170 456970 496226
rect 457026 496170 457094 496226
rect 457150 496170 457218 496226
rect 457274 496170 457342 496226
rect 457398 496170 492970 496226
rect 493026 496170 493094 496226
rect 493150 496170 493218 496226
rect 493274 496170 493342 496226
rect 493398 496170 510970 496226
rect 511026 496170 511094 496226
rect 511150 496170 511218 496226
rect 511274 496170 511342 496226
rect 511398 496170 528970 496226
rect 529026 496170 529094 496226
rect 529150 496170 529218 496226
rect 529274 496170 529342 496226
rect 529398 496170 546970 496226
rect 547026 496170 547094 496226
rect 547150 496170 547218 496226
rect 547274 496170 547342 496226
rect 547398 496170 568058 496226
rect 568114 496170 568182 496226
rect 568238 496170 574862 496226
rect 574918 496170 574986 496226
rect 575042 496170 581666 496226
rect 581722 496170 581790 496226
rect 581846 496170 582970 496226
rect 583026 496170 583094 496226
rect 583150 496170 583218 496226
rect 583274 496170 583342 496226
rect 583398 496170 588470 496226
rect 588526 496170 588594 496226
rect 588650 496170 597456 496226
rect 597512 496170 597580 496226
rect 597636 496170 597704 496226
rect 597760 496170 597828 496226
rect 597884 496170 597980 496226
rect -1916 496102 597980 496170
rect -1916 496046 -1820 496102
rect -1764 496046 -1696 496102
rect -1640 496046 -1572 496102
rect -1516 496046 -1448 496102
rect -1392 496046 6970 496102
rect 7026 496046 7094 496102
rect 7150 496046 7218 496102
rect 7274 496046 7342 496102
rect 7398 496046 24970 496102
rect 25026 496046 25094 496102
rect 25150 496046 25218 496102
rect 25274 496046 25342 496102
rect 25398 496046 42970 496102
rect 43026 496046 43094 496102
rect 43150 496046 43218 496102
rect 43274 496046 43342 496102
rect 43398 496046 60970 496102
rect 61026 496046 61094 496102
rect 61150 496046 61218 496102
rect 61274 496046 61342 496102
rect 61398 496046 78970 496102
rect 79026 496046 79094 496102
rect 79150 496046 79218 496102
rect 79274 496046 79342 496102
rect 79398 496046 96970 496102
rect 97026 496046 97094 496102
rect 97150 496046 97218 496102
rect 97274 496046 97342 496102
rect 97398 496046 132970 496102
rect 133026 496046 133094 496102
rect 133150 496046 133218 496102
rect 133274 496046 133342 496102
rect 133398 496046 150970 496102
rect 151026 496046 151094 496102
rect 151150 496046 151218 496102
rect 151274 496046 151342 496102
rect 151398 496046 168970 496102
rect 169026 496046 169094 496102
rect 169150 496046 169218 496102
rect 169274 496046 169342 496102
rect 169398 496046 186970 496102
rect 187026 496046 187094 496102
rect 187150 496046 187218 496102
rect 187274 496046 187342 496102
rect 187398 496046 222970 496102
rect 223026 496046 223094 496102
rect 223150 496046 223218 496102
rect 223274 496046 223342 496102
rect 223398 496046 240970 496102
rect 241026 496046 241094 496102
rect 241150 496046 241218 496102
rect 241274 496046 241342 496102
rect 241398 496046 258970 496102
rect 259026 496046 259094 496102
rect 259150 496046 259218 496102
rect 259274 496046 259342 496102
rect 259398 496046 276970 496102
rect 277026 496046 277094 496102
rect 277150 496046 277218 496102
rect 277274 496046 277342 496102
rect 277398 496046 312970 496102
rect 313026 496046 313094 496102
rect 313150 496046 313218 496102
rect 313274 496046 313342 496102
rect 313398 496046 330970 496102
rect 331026 496046 331094 496102
rect 331150 496046 331218 496102
rect 331274 496046 331342 496102
rect 331398 496046 348970 496102
rect 349026 496046 349094 496102
rect 349150 496046 349218 496102
rect 349274 496046 349342 496102
rect 349398 496046 366970 496102
rect 367026 496046 367094 496102
rect 367150 496046 367218 496102
rect 367274 496046 367342 496102
rect 367398 496046 402970 496102
rect 403026 496046 403094 496102
rect 403150 496046 403218 496102
rect 403274 496046 403342 496102
rect 403398 496046 420970 496102
rect 421026 496046 421094 496102
rect 421150 496046 421218 496102
rect 421274 496046 421342 496102
rect 421398 496046 438970 496102
rect 439026 496046 439094 496102
rect 439150 496046 439218 496102
rect 439274 496046 439342 496102
rect 439398 496046 456970 496102
rect 457026 496046 457094 496102
rect 457150 496046 457218 496102
rect 457274 496046 457342 496102
rect 457398 496046 492970 496102
rect 493026 496046 493094 496102
rect 493150 496046 493218 496102
rect 493274 496046 493342 496102
rect 493398 496046 510970 496102
rect 511026 496046 511094 496102
rect 511150 496046 511218 496102
rect 511274 496046 511342 496102
rect 511398 496046 528970 496102
rect 529026 496046 529094 496102
rect 529150 496046 529218 496102
rect 529274 496046 529342 496102
rect 529398 496046 546970 496102
rect 547026 496046 547094 496102
rect 547150 496046 547218 496102
rect 547274 496046 547342 496102
rect 547398 496046 568058 496102
rect 568114 496046 568182 496102
rect 568238 496046 574862 496102
rect 574918 496046 574986 496102
rect 575042 496046 581666 496102
rect 581722 496046 581790 496102
rect 581846 496046 582970 496102
rect 583026 496046 583094 496102
rect 583150 496046 583218 496102
rect 583274 496046 583342 496102
rect 583398 496046 588470 496102
rect 588526 496046 588594 496102
rect 588650 496046 597456 496102
rect 597512 496046 597580 496102
rect 597636 496046 597704 496102
rect 597760 496046 597828 496102
rect 597884 496046 597980 496102
rect -1916 495978 597980 496046
rect -1916 495922 -1820 495978
rect -1764 495922 -1696 495978
rect -1640 495922 -1572 495978
rect -1516 495922 -1448 495978
rect -1392 495922 6970 495978
rect 7026 495922 7094 495978
rect 7150 495922 7218 495978
rect 7274 495922 7342 495978
rect 7398 495922 24970 495978
rect 25026 495922 25094 495978
rect 25150 495922 25218 495978
rect 25274 495922 25342 495978
rect 25398 495922 42970 495978
rect 43026 495922 43094 495978
rect 43150 495922 43218 495978
rect 43274 495922 43342 495978
rect 43398 495922 60970 495978
rect 61026 495922 61094 495978
rect 61150 495922 61218 495978
rect 61274 495922 61342 495978
rect 61398 495922 78970 495978
rect 79026 495922 79094 495978
rect 79150 495922 79218 495978
rect 79274 495922 79342 495978
rect 79398 495922 96970 495978
rect 97026 495922 97094 495978
rect 97150 495922 97218 495978
rect 97274 495922 97342 495978
rect 97398 495922 132970 495978
rect 133026 495922 133094 495978
rect 133150 495922 133218 495978
rect 133274 495922 133342 495978
rect 133398 495922 150970 495978
rect 151026 495922 151094 495978
rect 151150 495922 151218 495978
rect 151274 495922 151342 495978
rect 151398 495922 168970 495978
rect 169026 495922 169094 495978
rect 169150 495922 169218 495978
rect 169274 495922 169342 495978
rect 169398 495922 186970 495978
rect 187026 495922 187094 495978
rect 187150 495922 187218 495978
rect 187274 495922 187342 495978
rect 187398 495922 222970 495978
rect 223026 495922 223094 495978
rect 223150 495922 223218 495978
rect 223274 495922 223342 495978
rect 223398 495922 240970 495978
rect 241026 495922 241094 495978
rect 241150 495922 241218 495978
rect 241274 495922 241342 495978
rect 241398 495922 258970 495978
rect 259026 495922 259094 495978
rect 259150 495922 259218 495978
rect 259274 495922 259342 495978
rect 259398 495922 276970 495978
rect 277026 495922 277094 495978
rect 277150 495922 277218 495978
rect 277274 495922 277342 495978
rect 277398 495922 312970 495978
rect 313026 495922 313094 495978
rect 313150 495922 313218 495978
rect 313274 495922 313342 495978
rect 313398 495922 330970 495978
rect 331026 495922 331094 495978
rect 331150 495922 331218 495978
rect 331274 495922 331342 495978
rect 331398 495922 348970 495978
rect 349026 495922 349094 495978
rect 349150 495922 349218 495978
rect 349274 495922 349342 495978
rect 349398 495922 366970 495978
rect 367026 495922 367094 495978
rect 367150 495922 367218 495978
rect 367274 495922 367342 495978
rect 367398 495922 402970 495978
rect 403026 495922 403094 495978
rect 403150 495922 403218 495978
rect 403274 495922 403342 495978
rect 403398 495922 420970 495978
rect 421026 495922 421094 495978
rect 421150 495922 421218 495978
rect 421274 495922 421342 495978
rect 421398 495922 438970 495978
rect 439026 495922 439094 495978
rect 439150 495922 439218 495978
rect 439274 495922 439342 495978
rect 439398 495922 456970 495978
rect 457026 495922 457094 495978
rect 457150 495922 457218 495978
rect 457274 495922 457342 495978
rect 457398 495922 492970 495978
rect 493026 495922 493094 495978
rect 493150 495922 493218 495978
rect 493274 495922 493342 495978
rect 493398 495922 510970 495978
rect 511026 495922 511094 495978
rect 511150 495922 511218 495978
rect 511274 495922 511342 495978
rect 511398 495922 528970 495978
rect 529026 495922 529094 495978
rect 529150 495922 529218 495978
rect 529274 495922 529342 495978
rect 529398 495922 546970 495978
rect 547026 495922 547094 495978
rect 547150 495922 547218 495978
rect 547274 495922 547342 495978
rect 547398 495922 568058 495978
rect 568114 495922 568182 495978
rect 568238 495922 574862 495978
rect 574918 495922 574986 495978
rect 575042 495922 581666 495978
rect 581722 495922 581790 495978
rect 581846 495922 582970 495978
rect 583026 495922 583094 495978
rect 583150 495922 583218 495978
rect 583274 495922 583342 495978
rect 583398 495922 588470 495978
rect 588526 495922 588594 495978
rect 588650 495922 597456 495978
rect 597512 495922 597580 495978
rect 597636 495922 597704 495978
rect 597760 495922 597828 495978
rect 597884 495922 597980 495978
rect -1916 495826 597980 495922
rect -1916 490350 597980 490446
rect -1916 490294 -860 490350
rect -804 490294 -736 490350
rect -680 490294 -612 490350
rect -556 490294 -488 490350
rect -432 490294 3250 490350
rect 3306 490294 3374 490350
rect 3430 490294 3498 490350
rect 3554 490294 3622 490350
rect 3678 490294 21250 490350
rect 21306 490294 21374 490350
rect 21430 490294 21498 490350
rect 21554 490294 21622 490350
rect 21678 490294 39250 490350
rect 39306 490294 39374 490350
rect 39430 490294 39498 490350
rect 39554 490294 39622 490350
rect 39678 490294 57250 490350
rect 57306 490294 57374 490350
rect 57430 490294 57498 490350
rect 57554 490294 57622 490350
rect 57678 490294 93250 490350
rect 93306 490294 93374 490350
rect 93430 490294 93498 490350
rect 93554 490294 93622 490350
rect 93678 490294 111250 490350
rect 111306 490294 111374 490350
rect 111430 490294 111498 490350
rect 111554 490294 111622 490350
rect 111678 490294 129250 490350
rect 129306 490294 129374 490350
rect 129430 490294 129498 490350
rect 129554 490294 129622 490350
rect 129678 490294 147250 490350
rect 147306 490294 147374 490350
rect 147430 490294 147498 490350
rect 147554 490294 147622 490350
rect 147678 490294 183250 490350
rect 183306 490294 183374 490350
rect 183430 490294 183498 490350
rect 183554 490294 183622 490350
rect 183678 490294 201250 490350
rect 201306 490294 201374 490350
rect 201430 490294 201498 490350
rect 201554 490294 201622 490350
rect 201678 490294 219250 490350
rect 219306 490294 219374 490350
rect 219430 490294 219498 490350
rect 219554 490294 219622 490350
rect 219678 490294 237250 490350
rect 237306 490294 237374 490350
rect 237430 490294 237498 490350
rect 237554 490294 237622 490350
rect 237678 490294 273250 490350
rect 273306 490294 273374 490350
rect 273430 490294 273498 490350
rect 273554 490294 273622 490350
rect 273678 490294 291250 490350
rect 291306 490294 291374 490350
rect 291430 490294 291498 490350
rect 291554 490294 291622 490350
rect 291678 490294 309250 490350
rect 309306 490294 309374 490350
rect 309430 490294 309498 490350
rect 309554 490294 309622 490350
rect 309678 490294 327250 490350
rect 327306 490294 327374 490350
rect 327430 490294 327498 490350
rect 327554 490294 327622 490350
rect 327678 490294 363250 490350
rect 363306 490294 363374 490350
rect 363430 490294 363498 490350
rect 363554 490294 363622 490350
rect 363678 490294 381250 490350
rect 381306 490294 381374 490350
rect 381430 490294 381498 490350
rect 381554 490294 381622 490350
rect 381678 490294 399250 490350
rect 399306 490294 399374 490350
rect 399430 490294 399498 490350
rect 399554 490294 399622 490350
rect 399678 490294 417250 490350
rect 417306 490294 417374 490350
rect 417430 490294 417498 490350
rect 417554 490294 417622 490350
rect 417678 490294 453250 490350
rect 453306 490294 453374 490350
rect 453430 490294 453498 490350
rect 453554 490294 453622 490350
rect 453678 490294 471250 490350
rect 471306 490294 471374 490350
rect 471430 490294 471498 490350
rect 471554 490294 471622 490350
rect 471678 490294 489250 490350
rect 489306 490294 489374 490350
rect 489430 490294 489498 490350
rect 489554 490294 489622 490350
rect 489678 490294 507250 490350
rect 507306 490294 507374 490350
rect 507430 490294 507498 490350
rect 507554 490294 507622 490350
rect 507678 490294 543250 490350
rect 543306 490294 543374 490350
rect 543430 490294 543498 490350
rect 543554 490294 543622 490350
rect 543678 490294 561250 490350
rect 561306 490294 561374 490350
rect 561430 490294 561498 490350
rect 561554 490294 561622 490350
rect 561678 490294 564656 490350
rect 564712 490294 564780 490350
rect 564836 490294 571460 490350
rect 571516 490294 571584 490350
rect 571640 490294 578264 490350
rect 578320 490294 578388 490350
rect 578444 490294 579250 490350
rect 579306 490294 579374 490350
rect 579430 490294 579498 490350
rect 579554 490294 579622 490350
rect 579678 490294 585068 490350
rect 585124 490294 585192 490350
rect 585248 490294 596496 490350
rect 596552 490294 596620 490350
rect 596676 490294 596744 490350
rect 596800 490294 596868 490350
rect 596924 490294 597980 490350
rect -1916 490226 597980 490294
rect -1916 490170 -860 490226
rect -804 490170 -736 490226
rect -680 490170 -612 490226
rect -556 490170 -488 490226
rect -432 490170 3250 490226
rect 3306 490170 3374 490226
rect 3430 490170 3498 490226
rect 3554 490170 3622 490226
rect 3678 490170 21250 490226
rect 21306 490170 21374 490226
rect 21430 490170 21498 490226
rect 21554 490170 21622 490226
rect 21678 490170 39250 490226
rect 39306 490170 39374 490226
rect 39430 490170 39498 490226
rect 39554 490170 39622 490226
rect 39678 490170 57250 490226
rect 57306 490170 57374 490226
rect 57430 490170 57498 490226
rect 57554 490170 57622 490226
rect 57678 490170 93250 490226
rect 93306 490170 93374 490226
rect 93430 490170 93498 490226
rect 93554 490170 93622 490226
rect 93678 490170 111250 490226
rect 111306 490170 111374 490226
rect 111430 490170 111498 490226
rect 111554 490170 111622 490226
rect 111678 490170 129250 490226
rect 129306 490170 129374 490226
rect 129430 490170 129498 490226
rect 129554 490170 129622 490226
rect 129678 490170 147250 490226
rect 147306 490170 147374 490226
rect 147430 490170 147498 490226
rect 147554 490170 147622 490226
rect 147678 490170 183250 490226
rect 183306 490170 183374 490226
rect 183430 490170 183498 490226
rect 183554 490170 183622 490226
rect 183678 490170 201250 490226
rect 201306 490170 201374 490226
rect 201430 490170 201498 490226
rect 201554 490170 201622 490226
rect 201678 490170 219250 490226
rect 219306 490170 219374 490226
rect 219430 490170 219498 490226
rect 219554 490170 219622 490226
rect 219678 490170 237250 490226
rect 237306 490170 237374 490226
rect 237430 490170 237498 490226
rect 237554 490170 237622 490226
rect 237678 490170 273250 490226
rect 273306 490170 273374 490226
rect 273430 490170 273498 490226
rect 273554 490170 273622 490226
rect 273678 490170 291250 490226
rect 291306 490170 291374 490226
rect 291430 490170 291498 490226
rect 291554 490170 291622 490226
rect 291678 490170 309250 490226
rect 309306 490170 309374 490226
rect 309430 490170 309498 490226
rect 309554 490170 309622 490226
rect 309678 490170 327250 490226
rect 327306 490170 327374 490226
rect 327430 490170 327498 490226
rect 327554 490170 327622 490226
rect 327678 490170 363250 490226
rect 363306 490170 363374 490226
rect 363430 490170 363498 490226
rect 363554 490170 363622 490226
rect 363678 490170 381250 490226
rect 381306 490170 381374 490226
rect 381430 490170 381498 490226
rect 381554 490170 381622 490226
rect 381678 490170 399250 490226
rect 399306 490170 399374 490226
rect 399430 490170 399498 490226
rect 399554 490170 399622 490226
rect 399678 490170 417250 490226
rect 417306 490170 417374 490226
rect 417430 490170 417498 490226
rect 417554 490170 417622 490226
rect 417678 490170 453250 490226
rect 453306 490170 453374 490226
rect 453430 490170 453498 490226
rect 453554 490170 453622 490226
rect 453678 490170 471250 490226
rect 471306 490170 471374 490226
rect 471430 490170 471498 490226
rect 471554 490170 471622 490226
rect 471678 490170 489250 490226
rect 489306 490170 489374 490226
rect 489430 490170 489498 490226
rect 489554 490170 489622 490226
rect 489678 490170 507250 490226
rect 507306 490170 507374 490226
rect 507430 490170 507498 490226
rect 507554 490170 507622 490226
rect 507678 490170 543250 490226
rect 543306 490170 543374 490226
rect 543430 490170 543498 490226
rect 543554 490170 543622 490226
rect 543678 490170 561250 490226
rect 561306 490170 561374 490226
rect 561430 490170 561498 490226
rect 561554 490170 561622 490226
rect 561678 490170 564656 490226
rect 564712 490170 564780 490226
rect 564836 490170 571460 490226
rect 571516 490170 571584 490226
rect 571640 490170 578264 490226
rect 578320 490170 578388 490226
rect 578444 490170 579250 490226
rect 579306 490170 579374 490226
rect 579430 490170 579498 490226
rect 579554 490170 579622 490226
rect 579678 490170 585068 490226
rect 585124 490170 585192 490226
rect 585248 490170 596496 490226
rect 596552 490170 596620 490226
rect 596676 490170 596744 490226
rect 596800 490170 596868 490226
rect 596924 490170 597980 490226
rect -1916 490102 597980 490170
rect -1916 490046 -860 490102
rect -804 490046 -736 490102
rect -680 490046 -612 490102
rect -556 490046 -488 490102
rect -432 490046 3250 490102
rect 3306 490046 3374 490102
rect 3430 490046 3498 490102
rect 3554 490046 3622 490102
rect 3678 490046 21250 490102
rect 21306 490046 21374 490102
rect 21430 490046 21498 490102
rect 21554 490046 21622 490102
rect 21678 490046 39250 490102
rect 39306 490046 39374 490102
rect 39430 490046 39498 490102
rect 39554 490046 39622 490102
rect 39678 490046 57250 490102
rect 57306 490046 57374 490102
rect 57430 490046 57498 490102
rect 57554 490046 57622 490102
rect 57678 490046 93250 490102
rect 93306 490046 93374 490102
rect 93430 490046 93498 490102
rect 93554 490046 93622 490102
rect 93678 490046 111250 490102
rect 111306 490046 111374 490102
rect 111430 490046 111498 490102
rect 111554 490046 111622 490102
rect 111678 490046 129250 490102
rect 129306 490046 129374 490102
rect 129430 490046 129498 490102
rect 129554 490046 129622 490102
rect 129678 490046 147250 490102
rect 147306 490046 147374 490102
rect 147430 490046 147498 490102
rect 147554 490046 147622 490102
rect 147678 490046 183250 490102
rect 183306 490046 183374 490102
rect 183430 490046 183498 490102
rect 183554 490046 183622 490102
rect 183678 490046 201250 490102
rect 201306 490046 201374 490102
rect 201430 490046 201498 490102
rect 201554 490046 201622 490102
rect 201678 490046 219250 490102
rect 219306 490046 219374 490102
rect 219430 490046 219498 490102
rect 219554 490046 219622 490102
rect 219678 490046 237250 490102
rect 237306 490046 237374 490102
rect 237430 490046 237498 490102
rect 237554 490046 237622 490102
rect 237678 490046 273250 490102
rect 273306 490046 273374 490102
rect 273430 490046 273498 490102
rect 273554 490046 273622 490102
rect 273678 490046 291250 490102
rect 291306 490046 291374 490102
rect 291430 490046 291498 490102
rect 291554 490046 291622 490102
rect 291678 490046 309250 490102
rect 309306 490046 309374 490102
rect 309430 490046 309498 490102
rect 309554 490046 309622 490102
rect 309678 490046 327250 490102
rect 327306 490046 327374 490102
rect 327430 490046 327498 490102
rect 327554 490046 327622 490102
rect 327678 490046 363250 490102
rect 363306 490046 363374 490102
rect 363430 490046 363498 490102
rect 363554 490046 363622 490102
rect 363678 490046 381250 490102
rect 381306 490046 381374 490102
rect 381430 490046 381498 490102
rect 381554 490046 381622 490102
rect 381678 490046 399250 490102
rect 399306 490046 399374 490102
rect 399430 490046 399498 490102
rect 399554 490046 399622 490102
rect 399678 490046 417250 490102
rect 417306 490046 417374 490102
rect 417430 490046 417498 490102
rect 417554 490046 417622 490102
rect 417678 490046 453250 490102
rect 453306 490046 453374 490102
rect 453430 490046 453498 490102
rect 453554 490046 453622 490102
rect 453678 490046 471250 490102
rect 471306 490046 471374 490102
rect 471430 490046 471498 490102
rect 471554 490046 471622 490102
rect 471678 490046 489250 490102
rect 489306 490046 489374 490102
rect 489430 490046 489498 490102
rect 489554 490046 489622 490102
rect 489678 490046 507250 490102
rect 507306 490046 507374 490102
rect 507430 490046 507498 490102
rect 507554 490046 507622 490102
rect 507678 490046 543250 490102
rect 543306 490046 543374 490102
rect 543430 490046 543498 490102
rect 543554 490046 543622 490102
rect 543678 490046 561250 490102
rect 561306 490046 561374 490102
rect 561430 490046 561498 490102
rect 561554 490046 561622 490102
rect 561678 490046 564656 490102
rect 564712 490046 564780 490102
rect 564836 490046 571460 490102
rect 571516 490046 571584 490102
rect 571640 490046 578264 490102
rect 578320 490046 578388 490102
rect 578444 490046 579250 490102
rect 579306 490046 579374 490102
rect 579430 490046 579498 490102
rect 579554 490046 579622 490102
rect 579678 490046 585068 490102
rect 585124 490046 585192 490102
rect 585248 490046 596496 490102
rect 596552 490046 596620 490102
rect 596676 490046 596744 490102
rect 596800 490046 596868 490102
rect 596924 490046 597980 490102
rect -1916 489978 597980 490046
rect -1916 489922 -860 489978
rect -804 489922 -736 489978
rect -680 489922 -612 489978
rect -556 489922 -488 489978
rect -432 489922 3250 489978
rect 3306 489922 3374 489978
rect 3430 489922 3498 489978
rect 3554 489922 3622 489978
rect 3678 489922 21250 489978
rect 21306 489922 21374 489978
rect 21430 489922 21498 489978
rect 21554 489922 21622 489978
rect 21678 489922 39250 489978
rect 39306 489922 39374 489978
rect 39430 489922 39498 489978
rect 39554 489922 39622 489978
rect 39678 489922 57250 489978
rect 57306 489922 57374 489978
rect 57430 489922 57498 489978
rect 57554 489922 57622 489978
rect 57678 489922 93250 489978
rect 93306 489922 93374 489978
rect 93430 489922 93498 489978
rect 93554 489922 93622 489978
rect 93678 489922 111250 489978
rect 111306 489922 111374 489978
rect 111430 489922 111498 489978
rect 111554 489922 111622 489978
rect 111678 489922 129250 489978
rect 129306 489922 129374 489978
rect 129430 489922 129498 489978
rect 129554 489922 129622 489978
rect 129678 489922 147250 489978
rect 147306 489922 147374 489978
rect 147430 489922 147498 489978
rect 147554 489922 147622 489978
rect 147678 489922 183250 489978
rect 183306 489922 183374 489978
rect 183430 489922 183498 489978
rect 183554 489922 183622 489978
rect 183678 489922 201250 489978
rect 201306 489922 201374 489978
rect 201430 489922 201498 489978
rect 201554 489922 201622 489978
rect 201678 489922 219250 489978
rect 219306 489922 219374 489978
rect 219430 489922 219498 489978
rect 219554 489922 219622 489978
rect 219678 489922 237250 489978
rect 237306 489922 237374 489978
rect 237430 489922 237498 489978
rect 237554 489922 237622 489978
rect 237678 489922 273250 489978
rect 273306 489922 273374 489978
rect 273430 489922 273498 489978
rect 273554 489922 273622 489978
rect 273678 489922 291250 489978
rect 291306 489922 291374 489978
rect 291430 489922 291498 489978
rect 291554 489922 291622 489978
rect 291678 489922 309250 489978
rect 309306 489922 309374 489978
rect 309430 489922 309498 489978
rect 309554 489922 309622 489978
rect 309678 489922 327250 489978
rect 327306 489922 327374 489978
rect 327430 489922 327498 489978
rect 327554 489922 327622 489978
rect 327678 489922 363250 489978
rect 363306 489922 363374 489978
rect 363430 489922 363498 489978
rect 363554 489922 363622 489978
rect 363678 489922 381250 489978
rect 381306 489922 381374 489978
rect 381430 489922 381498 489978
rect 381554 489922 381622 489978
rect 381678 489922 399250 489978
rect 399306 489922 399374 489978
rect 399430 489922 399498 489978
rect 399554 489922 399622 489978
rect 399678 489922 417250 489978
rect 417306 489922 417374 489978
rect 417430 489922 417498 489978
rect 417554 489922 417622 489978
rect 417678 489922 453250 489978
rect 453306 489922 453374 489978
rect 453430 489922 453498 489978
rect 453554 489922 453622 489978
rect 453678 489922 471250 489978
rect 471306 489922 471374 489978
rect 471430 489922 471498 489978
rect 471554 489922 471622 489978
rect 471678 489922 489250 489978
rect 489306 489922 489374 489978
rect 489430 489922 489498 489978
rect 489554 489922 489622 489978
rect 489678 489922 507250 489978
rect 507306 489922 507374 489978
rect 507430 489922 507498 489978
rect 507554 489922 507622 489978
rect 507678 489922 543250 489978
rect 543306 489922 543374 489978
rect 543430 489922 543498 489978
rect 543554 489922 543622 489978
rect 543678 489922 561250 489978
rect 561306 489922 561374 489978
rect 561430 489922 561498 489978
rect 561554 489922 561622 489978
rect 561678 489922 564656 489978
rect 564712 489922 564780 489978
rect 564836 489922 571460 489978
rect 571516 489922 571584 489978
rect 571640 489922 578264 489978
rect 578320 489922 578388 489978
rect 578444 489922 579250 489978
rect 579306 489922 579374 489978
rect 579430 489922 579498 489978
rect 579554 489922 579622 489978
rect 579678 489922 585068 489978
rect 585124 489922 585192 489978
rect 585248 489922 596496 489978
rect 596552 489922 596620 489978
rect 596676 489922 596744 489978
rect 596800 489922 596868 489978
rect 596924 489922 597980 489978
rect -1916 489826 597980 489922
rect -1916 478350 597980 478446
rect -1916 478294 -1820 478350
rect -1764 478294 -1696 478350
rect -1640 478294 -1572 478350
rect -1516 478294 -1448 478350
rect -1392 478294 6970 478350
rect 7026 478294 7094 478350
rect 7150 478294 7218 478350
rect 7274 478294 7342 478350
rect 7398 478294 24970 478350
rect 25026 478294 25094 478350
rect 25150 478294 25218 478350
rect 25274 478294 25342 478350
rect 25398 478294 42970 478350
rect 43026 478294 43094 478350
rect 43150 478294 43218 478350
rect 43274 478294 43342 478350
rect 43398 478294 60970 478350
rect 61026 478294 61094 478350
rect 61150 478294 61218 478350
rect 61274 478294 61342 478350
rect 61398 478294 78970 478350
rect 79026 478294 79094 478350
rect 79150 478294 79218 478350
rect 79274 478294 79342 478350
rect 79398 478294 96970 478350
rect 97026 478294 97094 478350
rect 97150 478294 97218 478350
rect 97274 478294 97342 478350
rect 97398 478294 132970 478350
rect 133026 478294 133094 478350
rect 133150 478294 133218 478350
rect 133274 478294 133342 478350
rect 133398 478294 150970 478350
rect 151026 478294 151094 478350
rect 151150 478294 151218 478350
rect 151274 478294 151342 478350
rect 151398 478294 168970 478350
rect 169026 478294 169094 478350
rect 169150 478294 169218 478350
rect 169274 478294 169342 478350
rect 169398 478294 186970 478350
rect 187026 478294 187094 478350
rect 187150 478294 187218 478350
rect 187274 478294 187342 478350
rect 187398 478294 222970 478350
rect 223026 478294 223094 478350
rect 223150 478294 223218 478350
rect 223274 478294 223342 478350
rect 223398 478294 240970 478350
rect 241026 478294 241094 478350
rect 241150 478294 241218 478350
rect 241274 478294 241342 478350
rect 241398 478294 258970 478350
rect 259026 478294 259094 478350
rect 259150 478294 259218 478350
rect 259274 478294 259342 478350
rect 259398 478294 276970 478350
rect 277026 478294 277094 478350
rect 277150 478294 277218 478350
rect 277274 478294 277342 478350
rect 277398 478294 312970 478350
rect 313026 478294 313094 478350
rect 313150 478294 313218 478350
rect 313274 478294 313342 478350
rect 313398 478294 330970 478350
rect 331026 478294 331094 478350
rect 331150 478294 331218 478350
rect 331274 478294 331342 478350
rect 331398 478294 348970 478350
rect 349026 478294 349094 478350
rect 349150 478294 349218 478350
rect 349274 478294 349342 478350
rect 349398 478294 366970 478350
rect 367026 478294 367094 478350
rect 367150 478294 367218 478350
rect 367274 478294 367342 478350
rect 367398 478294 402970 478350
rect 403026 478294 403094 478350
rect 403150 478294 403218 478350
rect 403274 478294 403342 478350
rect 403398 478294 420970 478350
rect 421026 478294 421094 478350
rect 421150 478294 421218 478350
rect 421274 478294 421342 478350
rect 421398 478294 438970 478350
rect 439026 478294 439094 478350
rect 439150 478294 439218 478350
rect 439274 478294 439342 478350
rect 439398 478294 456970 478350
rect 457026 478294 457094 478350
rect 457150 478294 457218 478350
rect 457274 478294 457342 478350
rect 457398 478294 492970 478350
rect 493026 478294 493094 478350
rect 493150 478294 493218 478350
rect 493274 478294 493342 478350
rect 493398 478294 510970 478350
rect 511026 478294 511094 478350
rect 511150 478294 511218 478350
rect 511274 478294 511342 478350
rect 511398 478294 528970 478350
rect 529026 478294 529094 478350
rect 529150 478294 529218 478350
rect 529274 478294 529342 478350
rect 529398 478294 546970 478350
rect 547026 478294 547094 478350
rect 547150 478294 547218 478350
rect 547274 478294 547342 478350
rect 547398 478294 568058 478350
rect 568114 478294 568182 478350
rect 568238 478294 574862 478350
rect 574918 478294 574986 478350
rect 575042 478294 581666 478350
rect 581722 478294 581790 478350
rect 581846 478294 588470 478350
rect 588526 478294 588594 478350
rect 588650 478294 597456 478350
rect 597512 478294 597580 478350
rect 597636 478294 597704 478350
rect 597760 478294 597828 478350
rect 597884 478294 597980 478350
rect -1916 478226 597980 478294
rect -1916 478170 -1820 478226
rect -1764 478170 -1696 478226
rect -1640 478170 -1572 478226
rect -1516 478170 -1448 478226
rect -1392 478170 6970 478226
rect 7026 478170 7094 478226
rect 7150 478170 7218 478226
rect 7274 478170 7342 478226
rect 7398 478170 24970 478226
rect 25026 478170 25094 478226
rect 25150 478170 25218 478226
rect 25274 478170 25342 478226
rect 25398 478170 42970 478226
rect 43026 478170 43094 478226
rect 43150 478170 43218 478226
rect 43274 478170 43342 478226
rect 43398 478170 60970 478226
rect 61026 478170 61094 478226
rect 61150 478170 61218 478226
rect 61274 478170 61342 478226
rect 61398 478170 78970 478226
rect 79026 478170 79094 478226
rect 79150 478170 79218 478226
rect 79274 478170 79342 478226
rect 79398 478170 96970 478226
rect 97026 478170 97094 478226
rect 97150 478170 97218 478226
rect 97274 478170 97342 478226
rect 97398 478170 132970 478226
rect 133026 478170 133094 478226
rect 133150 478170 133218 478226
rect 133274 478170 133342 478226
rect 133398 478170 150970 478226
rect 151026 478170 151094 478226
rect 151150 478170 151218 478226
rect 151274 478170 151342 478226
rect 151398 478170 168970 478226
rect 169026 478170 169094 478226
rect 169150 478170 169218 478226
rect 169274 478170 169342 478226
rect 169398 478170 186970 478226
rect 187026 478170 187094 478226
rect 187150 478170 187218 478226
rect 187274 478170 187342 478226
rect 187398 478170 222970 478226
rect 223026 478170 223094 478226
rect 223150 478170 223218 478226
rect 223274 478170 223342 478226
rect 223398 478170 240970 478226
rect 241026 478170 241094 478226
rect 241150 478170 241218 478226
rect 241274 478170 241342 478226
rect 241398 478170 258970 478226
rect 259026 478170 259094 478226
rect 259150 478170 259218 478226
rect 259274 478170 259342 478226
rect 259398 478170 276970 478226
rect 277026 478170 277094 478226
rect 277150 478170 277218 478226
rect 277274 478170 277342 478226
rect 277398 478170 312970 478226
rect 313026 478170 313094 478226
rect 313150 478170 313218 478226
rect 313274 478170 313342 478226
rect 313398 478170 330970 478226
rect 331026 478170 331094 478226
rect 331150 478170 331218 478226
rect 331274 478170 331342 478226
rect 331398 478170 348970 478226
rect 349026 478170 349094 478226
rect 349150 478170 349218 478226
rect 349274 478170 349342 478226
rect 349398 478170 366970 478226
rect 367026 478170 367094 478226
rect 367150 478170 367218 478226
rect 367274 478170 367342 478226
rect 367398 478170 402970 478226
rect 403026 478170 403094 478226
rect 403150 478170 403218 478226
rect 403274 478170 403342 478226
rect 403398 478170 420970 478226
rect 421026 478170 421094 478226
rect 421150 478170 421218 478226
rect 421274 478170 421342 478226
rect 421398 478170 438970 478226
rect 439026 478170 439094 478226
rect 439150 478170 439218 478226
rect 439274 478170 439342 478226
rect 439398 478170 456970 478226
rect 457026 478170 457094 478226
rect 457150 478170 457218 478226
rect 457274 478170 457342 478226
rect 457398 478170 492970 478226
rect 493026 478170 493094 478226
rect 493150 478170 493218 478226
rect 493274 478170 493342 478226
rect 493398 478170 510970 478226
rect 511026 478170 511094 478226
rect 511150 478170 511218 478226
rect 511274 478170 511342 478226
rect 511398 478170 528970 478226
rect 529026 478170 529094 478226
rect 529150 478170 529218 478226
rect 529274 478170 529342 478226
rect 529398 478170 546970 478226
rect 547026 478170 547094 478226
rect 547150 478170 547218 478226
rect 547274 478170 547342 478226
rect 547398 478170 568058 478226
rect 568114 478170 568182 478226
rect 568238 478170 574862 478226
rect 574918 478170 574986 478226
rect 575042 478170 581666 478226
rect 581722 478170 581790 478226
rect 581846 478170 588470 478226
rect 588526 478170 588594 478226
rect 588650 478170 597456 478226
rect 597512 478170 597580 478226
rect 597636 478170 597704 478226
rect 597760 478170 597828 478226
rect 597884 478170 597980 478226
rect -1916 478102 597980 478170
rect -1916 478046 -1820 478102
rect -1764 478046 -1696 478102
rect -1640 478046 -1572 478102
rect -1516 478046 -1448 478102
rect -1392 478046 6970 478102
rect 7026 478046 7094 478102
rect 7150 478046 7218 478102
rect 7274 478046 7342 478102
rect 7398 478046 24970 478102
rect 25026 478046 25094 478102
rect 25150 478046 25218 478102
rect 25274 478046 25342 478102
rect 25398 478046 42970 478102
rect 43026 478046 43094 478102
rect 43150 478046 43218 478102
rect 43274 478046 43342 478102
rect 43398 478046 60970 478102
rect 61026 478046 61094 478102
rect 61150 478046 61218 478102
rect 61274 478046 61342 478102
rect 61398 478046 78970 478102
rect 79026 478046 79094 478102
rect 79150 478046 79218 478102
rect 79274 478046 79342 478102
rect 79398 478046 96970 478102
rect 97026 478046 97094 478102
rect 97150 478046 97218 478102
rect 97274 478046 97342 478102
rect 97398 478046 132970 478102
rect 133026 478046 133094 478102
rect 133150 478046 133218 478102
rect 133274 478046 133342 478102
rect 133398 478046 150970 478102
rect 151026 478046 151094 478102
rect 151150 478046 151218 478102
rect 151274 478046 151342 478102
rect 151398 478046 168970 478102
rect 169026 478046 169094 478102
rect 169150 478046 169218 478102
rect 169274 478046 169342 478102
rect 169398 478046 186970 478102
rect 187026 478046 187094 478102
rect 187150 478046 187218 478102
rect 187274 478046 187342 478102
rect 187398 478046 222970 478102
rect 223026 478046 223094 478102
rect 223150 478046 223218 478102
rect 223274 478046 223342 478102
rect 223398 478046 240970 478102
rect 241026 478046 241094 478102
rect 241150 478046 241218 478102
rect 241274 478046 241342 478102
rect 241398 478046 258970 478102
rect 259026 478046 259094 478102
rect 259150 478046 259218 478102
rect 259274 478046 259342 478102
rect 259398 478046 276970 478102
rect 277026 478046 277094 478102
rect 277150 478046 277218 478102
rect 277274 478046 277342 478102
rect 277398 478046 312970 478102
rect 313026 478046 313094 478102
rect 313150 478046 313218 478102
rect 313274 478046 313342 478102
rect 313398 478046 330970 478102
rect 331026 478046 331094 478102
rect 331150 478046 331218 478102
rect 331274 478046 331342 478102
rect 331398 478046 348970 478102
rect 349026 478046 349094 478102
rect 349150 478046 349218 478102
rect 349274 478046 349342 478102
rect 349398 478046 366970 478102
rect 367026 478046 367094 478102
rect 367150 478046 367218 478102
rect 367274 478046 367342 478102
rect 367398 478046 402970 478102
rect 403026 478046 403094 478102
rect 403150 478046 403218 478102
rect 403274 478046 403342 478102
rect 403398 478046 420970 478102
rect 421026 478046 421094 478102
rect 421150 478046 421218 478102
rect 421274 478046 421342 478102
rect 421398 478046 438970 478102
rect 439026 478046 439094 478102
rect 439150 478046 439218 478102
rect 439274 478046 439342 478102
rect 439398 478046 456970 478102
rect 457026 478046 457094 478102
rect 457150 478046 457218 478102
rect 457274 478046 457342 478102
rect 457398 478046 492970 478102
rect 493026 478046 493094 478102
rect 493150 478046 493218 478102
rect 493274 478046 493342 478102
rect 493398 478046 510970 478102
rect 511026 478046 511094 478102
rect 511150 478046 511218 478102
rect 511274 478046 511342 478102
rect 511398 478046 528970 478102
rect 529026 478046 529094 478102
rect 529150 478046 529218 478102
rect 529274 478046 529342 478102
rect 529398 478046 546970 478102
rect 547026 478046 547094 478102
rect 547150 478046 547218 478102
rect 547274 478046 547342 478102
rect 547398 478046 568058 478102
rect 568114 478046 568182 478102
rect 568238 478046 574862 478102
rect 574918 478046 574986 478102
rect 575042 478046 581666 478102
rect 581722 478046 581790 478102
rect 581846 478046 588470 478102
rect 588526 478046 588594 478102
rect 588650 478046 597456 478102
rect 597512 478046 597580 478102
rect 597636 478046 597704 478102
rect 597760 478046 597828 478102
rect 597884 478046 597980 478102
rect -1916 477978 597980 478046
rect -1916 477922 -1820 477978
rect -1764 477922 -1696 477978
rect -1640 477922 -1572 477978
rect -1516 477922 -1448 477978
rect -1392 477922 6970 477978
rect 7026 477922 7094 477978
rect 7150 477922 7218 477978
rect 7274 477922 7342 477978
rect 7398 477922 24970 477978
rect 25026 477922 25094 477978
rect 25150 477922 25218 477978
rect 25274 477922 25342 477978
rect 25398 477922 42970 477978
rect 43026 477922 43094 477978
rect 43150 477922 43218 477978
rect 43274 477922 43342 477978
rect 43398 477922 60970 477978
rect 61026 477922 61094 477978
rect 61150 477922 61218 477978
rect 61274 477922 61342 477978
rect 61398 477922 78970 477978
rect 79026 477922 79094 477978
rect 79150 477922 79218 477978
rect 79274 477922 79342 477978
rect 79398 477922 96970 477978
rect 97026 477922 97094 477978
rect 97150 477922 97218 477978
rect 97274 477922 97342 477978
rect 97398 477922 132970 477978
rect 133026 477922 133094 477978
rect 133150 477922 133218 477978
rect 133274 477922 133342 477978
rect 133398 477922 150970 477978
rect 151026 477922 151094 477978
rect 151150 477922 151218 477978
rect 151274 477922 151342 477978
rect 151398 477922 168970 477978
rect 169026 477922 169094 477978
rect 169150 477922 169218 477978
rect 169274 477922 169342 477978
rect 169398 477922 186970 477978
rect 187026 477922 187094 477978
rect 187150 477922 187218 477978
rect 187274 477922 187342 477978
rect 187398 477922 222970 477978
rect 223026 477922 223094 477978
rect 223150 477922 223218 477978
rect 223274 477922 223342 477978
rect 223398 477922 240970 477978
rect 241026 477922 241094 477978
rect 241150 477922 241218 477978
rect 241274 477922 241342 477978
rect 241398 477922 258970 477978
rect 259026 477922 259094 477978
rect 259150 477922 259218 477978
rect 259274 477922 259342 477978
rect 259398 477922 276970 477978
rect 277026 477922 277094 477978
rect 277150 477922 277218 477978
rect 277274 477922 277342 477978
rect 277398 477922 312970 477978
rect 313026 477922 313094 477978
rect 313150 477922 313218 477978
rect 313274 477922 313342 477978
rect 313398 477922 330970 477978
rect 331026 477922 331094 477978
rect 331150 477922 331218 477978
rect 331274 477922 331342 477978
rect 331398 477922 348970 477978
rect 349026 477922 349094 477978
rect 349150 477922 349218 477978
rect 349274 477922 349342 477978
rect 349398 477922 366970 477978
rect 367026 477922 367094 477978
rect 367150 477922 367218 477978
rect 367274 477922 367342 477978
rect 367398 477922 402970 477978
rect 403026 477922 403094 477978
rect 403150 477922 403218 477978
rect 403274 477922 403342 477978
rect 403398 477922 420970 477978
rect 421026 477922 421094 477978
rect 421150 477922 421218 477978
rect 421274 477922 421342 477978
rect 421398 477922 438970 477978
rect 439026 477922 439094 477978
rect 439150 477922 439218 477978
rect 439274 477922 439342 477978
rect 439398 477922 456970 477978
rect 457026 477922 457094 477978
rect 457150 477922 457218 477978
rect 457274 477922 457342 477978
rect 457398 477922 492970 477978
rect 493026 477922 493094 477978
rect 493150 477922 493218 477978
rect 493274 477922 493342 477978
rect 493398 477922 510970 477978
rect 511026 477922 511094 477978
rect 511150 477922 511218 477978
rect 511274 477922 511342 477978
rect 511398 477922 528970 477978
rect 529026 477922 529094 477978
rect 529150 477922 529218 477978
rect 529274 477922 529342 477978
rect 529398 477922 546970 477978
rect 547026 477922 547094 477978
rect 547150 477922 547218 477978
rect 547274 477922 547342 477978
rect 547398 477922 568058 477978
rect 568114 477922 568182 477978
rect 568238 477922 574862 477978
rect 574918 477922 574986 477978
rect 575042 477922 581666 477978
rect 581722 477922 581790 477978
rect 581846 477922 588470 477978
rect 588526 477922 588594 477978
rect 588650 477922 597456 477978
rect 597512 477922 597580 477978
rect 597636 477922 597704 477978
rect 597760 477922 597828 477978
rect 597884 477922 597980 477978
rect -1916 477826 597980 477922
rect -1916 472350 597980 472446
rect -1916 472294 -860 472350
rect -804 472294 -736 472350
rect -680 472294 -612 472350
rect -556 472294 -488 472350
rect -432 472294 3250 472350
rect 3306 472294 3374 472350
rect 3430 472294 3498 472350
rect 3554 472294 3622 472350
rect 3678 472294 21250 472350
rect 21306 472294 21374 472350
rect 21430 472294 21498 472350
rect 21554 472294 21622 472350
rect 21678 472294 39250 472350
rect 39306 472294 39374 472350
rect 39430 472294 39498 472350
rect 39554 472294 39622 472350
rect 39678 472294 57250 472350
rect 57306 472294 57374 472350
rect 57430 472294 57498 472350
rect 57554 472294 57622 472350
rect 57678 472294 93250 472350
rect 93306 472294 93374 472350
rect 93430 472294 93498 472350
rect 93554 472294 93622 472350
rect 93678 472294 111250 472350
rect 111306 472294 111374 472350
rect 111430 472294 111498 472350
rect 111554 472294 111622 472350
rect 111678 472294 129250 472350
rect 129306 472294 129374 472350
rect 129430 472294 129498 472350
rect 129554 472294 129622 472350
rect 129678 472294 147250 472350
rect 147306 472294 147374 472350
rect 147430 472294 147498 472350
rect 147554 472294 147622 472350
rect 147678 472294 183250 472350
rect 183306 472294 183374 472350
rect 183430 472294 183498 472350
rect 183554 472294 183622 472350
rect 183678 472294 201250 472350
rect 201306 472294 201374 472350
rect 201430 472294 201498 472350
rect 201554 472294 201622 472350
rect 201678 472294 219250 472350
rect 219306 472294 219374 472350
rect 219430 472294 219498 472350
rect 219554 472294 219622 472350
rect 219678 472294 237250 472350
rect 237306 472294 237374 472350
rect 237430 472294 237498 472350
rect 237554 472294 237622 472350
rect 237678 472294 273250 472350
rect 273306 472294 273374 472350
rect 273430 472294 273498 472350
rect 273554 472294 273622 472350
rect 273678 472294 291250 472350
rect 291306 472294 291374 472350
rect 291430 472294 291498 472350
rect 291554 472294 291622 472350
rect 291678 472294 309250 472350
rect 309306 472294 309374 472350
rect 309430 472294 309498 472350
rect 309554 472294 309622 472350
rect 309678 472294 327250 472350
rect 327306 472294 327374 472350
rect 327430 472294 327498 472350
rect 327554 472294 327622 472350
rect 327678 472294 363250 472350
rect 363306 472294 363374 472350
rect 363430 472294 363498 472350
rect 363554 472294 363622 472350
rect 363678 472294 381250 472350
rect 381306 472294 381374 472350
rect 381430 472294 381498 472350
rect 381554 472294 381622 472350
rect 381678 472294 399250 472350
rect 399306 472294 399374 472350
rect 399430 472294 399498 472350
rect 399554 472294 399622 472350
rect 399678 472294 417250 472350
rect 417306 472294 417374 472350
rect 417430 472294 417498 472350
rect 417554 472294 417622 472350
rect 417678 472294 453250 472350
rect 453306 472294 453374 472350
rect 453430 472294 453498 472350
rect 453554 472294 453622 472350
rect 453678 472294 471250 472350
rect 471306 472294 471374 472350
rect 471430 472294 471498 472350
rect 471554 472294 471622 472350
rect 471678 472294 489250 472350
rect 489306 472294 489374 472350
rect 489430 472294 489498 472350
rect 489554 472294 489622 472350
rect 489678 472294 507250 472350
rect 507306 472294 507374 472350
rect 507430 472294 507498 472350
rect 507554 472294 507622 472350
rect 507678 472294 543250 472350
rect 543306 472294 543374 472350
rect 543430 472294 543498 472350
rect 543554 472294 543622 472350
rect 543678 472294 564656 472350
rect 564712 472294 564780 472350
rect 564836 472294 571460 472350
rect 571516 472294 571584 472350
rect 571640 472294 578264 472350
rect 578320 472294 578388 472350
rect 578444 472294 585068 472350
rect 585124 472294 585192 472350
rect 585248 472294 596496 472350
rect 596552 472294 596620 472350
rect 596676 472294 596744 472350
rect 596800 472294 596868 472350
rect 596924 472294 597980 472350
rect -1916 472226 597980 472294
rect -1916 472170 -860 472226
rect -804 472170 -736 472226
rect -680 472170 -612 472226
rect -556 472170 -488 472226
rect -432 472170 3250 472226
rect 3306 472170 3374 472226
rect 3430 472170 3498 472226
rect 3554 472170 3622 472226
rect 3678 472170 21250 472226
rect 21306 472170 21374 472226
rect 21430 472170 21498 472226
rect 21554 472170 21622 472226
rect 21678 472170 39250 472226
rect 39306 472170 39374 472226
rect 39430 472170 39498 472226
rect 39554 472170 39622 472226
rect 39678 472170 57250 472226
rect 57306 472170 57374 472226
rect 57430 472170 57498 472226
rect 57554 472170 57622 472226
rect 57678 472170 93250 472226
rect 93306 472170 93374 472226
rect 93430 472170 93498 472226
rect 93554 472170 93622 472226
rect 93678 472170 111250 472226
rect 111306 472170 111374 472226
rect 111430 472170 111498 472226
rect 111554 472170 111622 472226
rect 111678 472170 129250 472226
rect 129306 472170 129374 472226
rect 129430 472170 129498 472226
rect 129554 472170 129622 472226
rect 129678 472170 147250 472226
rect 147306 472170 147374 472226
rect 147430 472170 147498 472226
rect 147554 472170 147622 472226
rect 147678 472170 183250 472226
rect 183306 472170 183374 472226
rect 183430 472170 183498 472226
rect 183554 472170 183622 472226
rect 183678 472170 201250 472226
rect 201306 472170 201374 472226
rect 201430 472170 201498 472226
rect 201554 472170 201622 472226
rect 201678 472170 219250 472226
rect 219306 472170 219374 472226
rect 219430 472170 219498 472226
rect 219554 472170 219622 472226
rect 219678 472170 237250 472226
rect 237306 472170 237374 472226
rect 237430 472170 237498 472226
rect 237554 472170 237622 472226
rect 237678 472170 273250 472226
rect 273306 472170 273374 472226
rect 273430 472170 273498 472226
rect 273554 472170 273622 472226
rect 273678 472170 291250 472226
rect 291306 472170 291374 472226
rect 291430 472170 291498 472226
rect 291554 472170 291622 472226
rect 291678 472170 309250 472226
rect 309306 472170 309374 472226
rect 309430 472170 309498 472226
rect 309554 472170 309622 472226
rect 309678 472170 327250 472226
rect 327306 472170 327374 472226
rect 327430 472170 327498 472226
rect 327554 472170 327622 472226
rect 327678 472170 363250 472226
rect 363306 472170 363374 472226
rect 363430 472170 363498 472226
rect 363554 472170 363622 472226
rect 363678 472170 381250 472226
rect 381306 472170 381374 472226
rect 381430 472170 381498 472226
rect 381554 472170 381622 472226
rect 381678 472170 399250 472226
rect 399306 472170 399374 472226
rect 399430 472170 399498 472226
rect 399554 472170 399622 472226
rect 399678 472170 417250 472226
rect 417306 472170 417374 472226
rect 417430 472170 417498 472226
rect 417554 472170 417622 472226
rect 417678 472170 453250 472226
rect 453306 472170 453374 472226
rect 453430 472170 453498 472226
rect 453554 472170 453622 472226
rect 453678 472170 471250 472226
rect 471306 472170 471374 472226
rect 471430 472170 471498 472226
rect 471554 472170 471622 472226
rect 471678 472170 489250 472226
rect 489306 472170 489374 472226
rect 489430 472170 489498 472226
rect 489554 472170 489622 472226
rect 489678 472170 507250 472226
rect 507306 472170 507374 472226
rect 507430 472170 507498 472226
rect 507554 472170 507622 472226
rect 507678 472170 543250 472226
rect 543306 472170 543374 472226
rect 543430 472170 543498 472226
rect 543554 472170 543622 472226
rect 543678 472170 564656 472226
rect 564712 472170 564780 472226
rect 564836 472170 571460 472226
rect 571516 472170 571584 472226
rect 571640 472170 578264 472226
rect 578320 472170 578388 472226
rect 578444 472170 585068 472226
rect 585124 472170 585192 472226
rect 585248 472170 596496 472226
rect 596552 472170 596620 472226
rect 596676 472170 596744 472226
rect 596800 472170 596868 472226
rect 596924 472170 597980 472226
rect -1916 472102 597980 472170
rect -1916 472046 -860 472102
rect -804 472046 -736 472102
rect -680 472046 -612 472102
rect -556 472046 -488 472102
rect -432 472046 3250 472102
rect 3306 472046 3374 472102
rect 3430 472046 3498 472102
rect 3554 472046 3622 472102
rect 3678 472046 21250 472102
rect 21306 472046 21374 472102
rect 21430 472046 21498 472102
rect 21554 472046 21622 472102
rect 21678 472046 39250 472102
rect 39306 472046 39374 472102
rect 39430 472046 39498 472102
rect 39554 472046 39622 472102
rect 39678 472046 57250 472102
rect 57306 472046 57374 472102
rect 57430 472046 57498 472102
rect 57554 472046 57622 472102
rect 57678 472046 93250 472102
rect 93306 472046 93374 472102
rect 93430 472046 93498 472102
rect 93554 472046 93622 472102
rect 93678 472046 111250 472102
rect 111306 472046 111374 472102
rect 111430 472046 111498 472102
rect 111554 472046 111622 472102
rect 111678 472046 129250 472102
rect 129306 472046 129374 472102
rect 129430 472046 129498 472102
rect 129554 472046 129622 472102
rect 129678 472046 147250 472102
rect 147306 472046 147374 472102
rect 147430 472046 147498 472102
rect 147554 472046 147622 472102
rect 147678 472046 183250 472102
rect 183306 472046 183374 472102
rect 183430 472046 183498 472102
rect 183554 472046 183622 472102
rect 183678 472046 201250 472102
rect 201306 472046 201374 472102
rect 201430 472046 201498 472102
rect 201554 472046 201622 472102
rect 201678 472046 219250 472102
rect 219306 472046 219374 472102
rect 219430 472046 219498 472102
rect 219554 472046 219622 472102
rect 219678 472046 237250 472102
rect 237306 472046 237374 472102
rect 237430 472046 237498 472102
rect 237554 472046 237622 472102
rect 237678 472046 273250 472102
rect 273306 472046 273374 472102
rect 273430 472046 273498 472102
rect 273554 472046 273622 472102
rect 273678 472046 291250 472102
rect 291306 472046 291374 472102
rect 291430 472046 291498 472102
rect 291554 472046 291622 472102
rect 291678 472046 309250 472102
rect 309306 472046 309374 472102
rect 309430 472046 309498 472102
rect 309554 472046 309622 472102
rect 309678 472046 327250 472102
rect 327306 472046 327374 472102
rect 327430 472046 327498 472102
rect 327554 472046 327622 472102
rect 327678 472046 363250 472102
rect 363306 472046 363374 472102
rect 363430 472046 363498 472102
rect 363554 472046 363622 472102
rect 363678 472046 381250 472102
rect 381306 472046 381374 472102
rect 381430 472046 381498 472102
rect 381554 472046 381622 472102
rect 381678 472046 399250 472102
rect 399306 472046 399374 472102
rect 399430 472046 399498 472102
rect 399554 472046 399622 472102
rect 399678 472046 417250 472102
rect 417306 472046 417374 472102
rect 417430 472046 417498 472102
rect 417554 472046 417622 472102
rect 417678 472046 453250 472102
rect 453306 472046 453374 472102
rect 453430 472046 453498 472102
rect 453554 472046 453622 472102
rect 453678 472046 471250 472102
rect 471306 472046 471374 472102
rect 471430 472046 471498 472102
rect 471554 472046 471622 472102
rect 471678 472046 489250 472102
rect 489306 472046 489374 472102
rect 489430 472046 489498 472102
rect 489554 472046 489622 472102
rect 489678 472046 507250 472102
rect 507306 472046 507374 472102
rect 507430 472046 507498 472102
rect 507554 472046 507622 472102
rect 507678 472046 543250 472102
rect 543306 472046 543374 472102
rect 543430 472046 543498 472102
rect 543554 472046 543622 472102
rect 543678 472046 564656 472102
rect 564712 472046 564780 472102
rect 564836 472046 571460 472102
rect 571516 472046 571584 472102
rect 571640 472046 578264 472102
rect 578320 472046 578388 472102
rect 578444 472046 585068 472102
rect 585124 472046 585192 472102
rect 585248 472046 596496 472102
rect 596552 472046 596620 472102
rect 596676 472046 596744 472102
rect 596800 472046 596868 472102
rect 596924 472046 597980 472102
rect -1916 471978 597980 472046
rect -1916 471922 -860 471978
rect -804 471922 -736 471978
rect -680 471922 -612 471978
rect -556 471922 -488 471978
rect -432 471922 3250 471978
rect 3306 471922 3374 471978
rect 3430 471922 3498 471978
rect 3554 471922 3622 471978
rect 3678 471922 21250 471978
rect 21306 471922 21374 471978
rect 21430 471922 21498 471978
rect 21554 471922 21622 471978
rect 21678 471922 39250 471978
rect 39306 471922 39374 471978
rect 39430 471922 39498 471978
rect 39554 471922 39622 471978
rect 39678 471922 57250 471978
rect 57306 471922 57374 471978
rect 57430 471922 57498 471978
rect 57554 471922 57622 471978
rect 57678 471922 93250 471978
rect 93306 471922 93374 471978
rect 93430 471922 93498 471978
rect 93554 471922 93622 471978
rect 93678 471922 111250 471978
rect 111306 471922 111374 471978
rect 111430 471922 111498 471978
rect 111554 471922 111622 471978
rect 111678 471922 129250 471978
rect 129306 471922 129374 471978
rect 129430 471922 129498 471978
rect 129554 471922 129622 471978
rect 129678 471922 147250 471978
rect 147306 471922 147374 471978
rect 147430 471922 147498 471978
rect 147554 471922 147622 471978
rect 147678 471922 183250 471978
rect 183306 471922 183374 471978
rect 183430 471922 183498 471978
rect 183554 471922 183622 471978
rect 183678 471922 201250 471978
rect 201306 471922 201374 471978
rect 201430 471922 201498 471978
rect 201554 471922 201622 471978
rect 201678 471922 219250 471978
rect 219306 471922 219374 471978
rect 219430 471922 219498 471978
rect 219554 471922 219622 471978
rect 219678 471922 237250 471978
rect 237306 471922 237374 471978
rect 237430 471922 237498 471978
rect 237554 471922 237622 471978
rect 237678 471922 273250 471978
rect 273306 471922 273374 471978
rect 273430 471922 273498 471978
rect 273554 471922 273622 471978
rect 273678 471922 291250 471978
rect 291306 471922 291374 471978
rect 291430 471922 291498 471978
rect 291554 471922 291622 471978
rect 291678 471922 309250 471978
rect 309306 471922 309374 471978
rect 309430 471922 309498 471978
rect 309554 471922 309622 471978
rect 309678 471922 327250 471978
rect 327306 471922 327374 471978
rect 327430 471922 327498 471978
rect 327554 471922 327622 471978
rect 327678 471922 363250 471978
rect 363306 471922 363374 471978
rect 363430 471922 363498 471978
rect 363554 471922 363622 471978
rect 363678 471922 381250 471978
rect 381306 471922 381374 471978
rect 381430 471922 381498 471978
rect 381554 471922 381622 471978
rect 381678 471922 399250 471978
rect 399306 471922 399374 471978
rect 399430 471922 399498 471978
rect 399554 471922 399622 471978
rect 399678 471922 417250 471978
rect 417306 471922 417374 471978
rect 417430 471922 417498 471978
rect 417554 471922 417622 471978
rect 417678 471922 453250 471978
rect 453306 471922 453374 471978
rect 453430 471922 453498 471978
rect 453554 471922 453622 471978
rect 453678 471922 471250 471978
rect 471306 471922 471374 471978
rect 471430 471922 471498 471978
rect 471554 471922 471622 471978
rect 471678 471922 489250 471978
rect 489306 471922 489374 471978
rect 489430 471922 489498 471978
rect 489554 471922 489622 471978
rect 489678 471922 507250 471978
rect 507306 471922 507374 471978
rect 507430 471922 507498 471978
rect 507554 471922 507622 471978
rect 507678 471922 543250 471978
rect 543306 471922 543374 471978
rect 543430 471922 543498 471978
rect 543554 471922 543622 471978
rect 543678 471922 564656 471978
rect 564712 471922 564780 471978
rect 564836 471922 571460 471978
rect 571516 471922 571584 471978
rect 571640 471922 578264 471978
rect 578320 471922 578388 471978
rect 578444 471922 585068 471978
rect 585124 471922 585192 471978
rect 585248 471922 596496 471978
rect 596552 471922 596620 471978
rect 596676 471922 596744 471978
rect 596800 471922 596868 471978
rect 596924 471922 597980 471978
rect -1916 471826 597980 471922
rect -1916 460350 597980 460446
rect -1916 460294 -1820 460350
rect -1764 460294 -1696 460350
rect -1640 460294 -1572 460350
rect -1516 460294 -1448 460350
rect -1392 460294 6970 460350
rect 7026 460294 7094 460350
rect 7150 460294 7218 460350
rect 7274 460294 7342 460350
rect 7398 460294 24970 460350
rect 25026 460294 25094 460350
rect 25150 460294 25218 460350
rect 25274 460294 25342 460350
rect 25398 460294 42970 460350
rect 43026 460294 43094 460350
rect 43150 460294 43218 460350
rect 43274 460294 43342 460350
rect 43398 460294 60970 460350
rect 61026 460294 61094 460350
rect 61150 460294 61218 460350
rect 61274 460294 61342 460350
rect 61398 460294 78970 460350
rect 79026 460294 79094 460350
rect 79150 460294 79218 460350
rect 79274 460294 79342 460350
rect 79398 460294 96970 460350
rect 97026 460294 97094 460350
rect 97150 460294 97218 460350
rect 97274 460294 97342 460350
rect 97398 460294 132970 460350
rect 133026 460294 133094 460350
rect 133150 460294 133218 460350
rect 133274 460294 133342 460350
rect 133398 460294 150970 460350
rect 151026 460294 151094 460350
rect 151150 460294 151218 460350
rect 151274 460294 151342 460350
rect 151398 460294 168970 460350
rect 169026 460294 169094 460350
rect 169150 460294 169218 460350
rect 169274 460294 169342 460350
rect 169398 460294 186970 460350
rect 187026 460294 187094 460350
rect 187150 460294 187218 460350
rect 187274 460294 187342 460350
rect 187398 460294 222970 460350
rect 223026 460294 223094 460350
rect 223150 460294 223218 460350
rect 223274 460294 223342 460350
rect 223398 460294 240970 460350
rect 241026 460294 241094 460350
rect 241150 460294 241218 460350
rect 241274 460294 241342 460350
rect 241398 460294 258970 460350
rect 259026 460294 259094 460350
rect 259150 460294 259218 460350
rect 259274 460294 259342 460350
rect 259398 460294 276970 460350
rect 277026 460294 277094 460350
rect 277150 460294 277218 460350
rect 277274 460294 277342 460350
rect 277398 460294 312970 460350
rect 313026 460294 313094 460350
rect 313150 460294 313218 460350
rect 313274 460294 313342 460350
rect 313398 460294 330970 460350
rect 331026 460294 331094 460350
rect 331150 460294 331218 460350
rect 331274 460294 331342 460350
rect 331398 460294 348970 460350
rect 349026 460294 349094 460350
rect 349150 460294 349218 460350
rect 349274 460294 349342 460350
rect 349398 460294 366970 460350
rect 367026 460294 367094 460350
rect 367150 460294 367218 460350
rect 367274 460294 367342 460350
rect 367398 460294 402970 460350
rect 403026 460294 403094 460350
rect 403150 460294 403218 460350
rect 403274 460294 403342 460350
rect 403398 460294 420970 460350
rect 421026 460294 421094 460350
rect 421150 460294 421218 460350
rect 421274 460294 421342 460350
rect 421398 460294 438970 460350
rect 439026 460294 439094 460350
rect 439150 460294 439218 460350
rect 439274 460294 439342 460350
rect 439398 460294 456970 460350
rect 457026 460294 457094 460350
rect 457150 460294 457218 460350
rect 457274 460294 457342 460350
rect 457398 460294 492970 460350
rect 493026 460294 493094 460350
rect 493150 460294 493218 460350
rect 493274 460294 493342 460350
rect 493398 460294 510970 460350
rect 511026 460294 511094 460350
rect 511150 460294 511218 460350
rect 511274 460294 511342 460350
rect 511398 460294 528970 460350
rect 529026 460294 529094 460350
rect 529150 460294 529218 460350
rect 529274 460294 529342 460350
rect 529398 460294 546970 460350
rect 547026 460294 547094 460350
rect 547150 460294 547218 460350
rect 547274 460294 547342 460350
rect 547398 460294 568058 460350
rect 568114 460294 568182 460350
rect 568238 460294 574862 460350
rect 574918 460294 574986 460350
rect 575042 460294 581666 460350
rect 581722 460294 581790 460350
rect 581846 460294 588470 460350
rect 588526 460294 588594 460350
rect 588650 460294 597456 460350
rect 597512 460294 597580 460350
rect 597636 460294 597704 460350
rect 597760 460294 597828 460350
rect 597884 460294 597980 460350
rect -1916 460226 597980 460294
rect -1916 460170 -1820 460226
rect -1764 460170 -1696 460226
rect -1640 460170 -1572 460226
rect -1516 460170 -1448 460226
rect -1392 460170 6970 460226
rect 7026 460170 7094 460226
rect 7150 460170 7218 460226
rect 7274 460170 7342 460226
rect 7398 460170 24970 460226
rect 25026 460170 25094 460226
rect 25150 460170 25218 460226
rect 25274 460170 25342 460226
rect 25398 460170 42970 460226
rect 43026 460170 43094 460226
rect 43150 460170 43218 460226
rect 43274 460170 43342 460226
rect 43398 460170 60970 460226
rect 61026 460170 61094 460226
rect 61150 460170 61218 460226
rect 61274 460170 61342 460226
rect 61398 460170 78970 460226
rect 79026 460170 79094 460226
rect 79150 460170 79218 460226
rect 79274 460170 79342 460226
rect 79398 460170 96970 460226
rect 97026 460170 97094 460226
rect 97150 460170 97218 460226
rect 97274 460170 97342 460226
rect 97398 460170 132970 460226
rect 133026 460170 133094 460226
rect 133150 460170 133218 460226
rect 133274 460170 133342 460226
rect 133398 460170 150970 460226
rect 151026 460170 151094 460226
rect 151150 460170 151218 460226
rect 151274 460170 151342 460226
rect 151398 460170 168970 460226
rect 169026 460170 169094 460226
rect 169150 460170 169218 460226
rect 169274 460170 169342 460226
rect 169398 460170 186970 460226
rect 187026 460170 187094 460226
rect 187150 460170 187218 460226
rect 187274 460170 187342 460226
rect 187398 460170 222970 460226
rect 223026 460170 223094 460226
rect 223150 460170 223218 460226
rect 223274 460170 223342 460226
rect 223398 460170 240970 460226
rect 241026 460170 241094 460226
rect 241150 460170 241218 460226
rect 241274 460170 241342 460226
rect 241398 460170 258970 460226
rect 259026 460170 259094 460226
rect 259150 460170 259218 460226
rect 259274 460170 259342 460226
rect 259398 460170 276970 460226
rect 277026 460170 277094 460226
rect 277150 460170 277218 460226
rect 277274 460170 277342 460226
rect 277398 460170 312970 460226
rect 313026 460170 313094 460226
rect 313150 460170 313218 460226
rect 313274 460170 313342 460226
rect 313398 460170 330970 460226
rect 331026 460170 331094 460226
rect 331150 460170 331218 460226
rect 331274 460170 331342 460226
rect 331398 460170 348970 460226
rect 349026 460170 349094 460226
rect 349150 460170 349218 460226
rect 349274 460170 349342 460226
rect 349398 460170 366970 460226
rect 367026 460170 367094 460226
rect 367150 460170 367218 460226
rect 367274 460170 367342 460226
rect 367398 460170 402970 460226
rect 403026 460170 403094 460226
rect 403150 460170 403218 460226
rect 403274 460170 403342 460226
rect 403398 460170 420970 460226
rect 421026 460170 421094 460226
rect 421150 460170 421218 460226
rect 421274 460170 421342 460226
rect 421398 460170 438970 460226
rect 439026 460170 439094 460226
rect 439150 460170 439218 460226
rect 439274 460170 439342 460226
rect 439398 460170 456970 460226
rect 457026 460170 457094 460226
rect 457150 460170 457218 460226
rect 457274 460170 457342 460226
rect 457398 460170 492970 460226
rect 493026 460170 493094 460226
rect 493150 460170 493218 460226
rect 493274 460170 493342 460226
rect 493398 460170 510970 460226
rect 511026 460170 511094 460226
rect 511150 460170 511218 460226
rect 511274 460170 511342 460226
rect 511398 460170 528970 460226
rect 529026 460170 529094 460226
rect 529150 460170 529218 460226
rect 529274 460170 529342 460226
rect 529398 460170 546970 460226
rect 547026 460170 547094 460226
rect 547150 460170 547218 460226
rect 547274 460170 547342 460226
rect 547398 460170 568058 460226
rect 568114 460170 568182 460226
rect 568238 460170 574862 460226
rect 574918 460170 574986 460226
rect 575042 460170 581666 460226
rect 581722 460170 581790 460226
rect 581846 460170 588470 460226
rect 588526 460170 588594 460226
rect 588650 460170 597456 460226
rect 597512 460170 597580 460226
rect 597636 460170 597704 460226
rect 597760 460170 597828 460226
rect 597884 460170 597980 460226
rect -1916 460102 597980 460170
rect -1916 460046 -1820 460102
rect -1764 460046 -1696 460102
rect -1640 460046 -1572 460102
rect -1516 460046 -1448 460102
rect -1392 460046 6970 460102
rect 7026 460046 7094 460102
rect 7150 460046 7218 460102
rect 7274 460046 7342 460102
rect 7398 460046 24970 460102
rect 25026 460046 25094 460102
rect 25150 460046 25218 460102
rect 25274 460046 25342 460102
rect 25398 460046 42970 460102
rect 43026 460046 43094 460102
rect 43150 460046 43218 460102
rect 43274 460046 43342 460102
rect 43398 460046 60970 460102
rect 61026 460046 61094 460102
rect 61150 460046 61218 460102
rect 61274 460046 61342 460102
rect 61398 460046 78970 460102
rect 79026 460046 79094 460102
rect 79150 460046 79218 460102
rect 79274 460046 79342 460102
rect 79398 460046 96970 460102
rect 97026 460046 97094 460102
rect 97150 460046 97218 460102
rect 97274 460046 97342 460102
rect 97398 460046 132970 460102
rect 133026 460046 133094 460102
rect 133150 460046 133218 460102
rect 133274 460046 133342 460102
rect 133398 460046 150970 460102
rect 151026 460046 151094 460102
rect 151150 460046 151218 460102
rect 151274 460046 151342 460102
rect 151398 460046 168970 460102
rect 169026 460046 169094 460102
rect 169150 460046 169218 460102
rect 169274 460046 169342 460102
rect 169398 460046 186970 460102
rect 187026 460046 187094 460102
rect 187150 460046 187218 460102
rect 187274 460046 187342 460102
rect 187398 460046 222970 460102
rect 223026 460046 223094 460102
rect 223150 460046 223218 460102
rect 223274 460046 223342 460102
rect 223398 460046 240970 460102
rect 241026 460046 241094 460102
rect 241150 460046 241218 460102
rect 241274 460046 241342 460102
rect 241398 460046 258970 460102
rect 259026 460046 259094 460102
rect 259150 460046 259218 460102
rect 259274 460046 259342 460102
rect 259398 460046 276970 460102
rect 277026 460046 277094 460102
rect 277150 460046 277218 460102
rect 277274 460046 277342 460102
rect 277398 460046 312970 460102
rect 313026 460046 313094 460102
rect 313150 460046 313218 460102
rect 313274 460046 313342 460102
rect 313398 460046 330970 460102
rect 331026 460046 331094 460102
rect 331150 460046 331218 460102
rect 331274 460046 331342 460102
rect 331398 460046 348970 460102
rect 349026 460046 349094 460102
rect 349150 460046 349218 460102
rect 349274 460046 349342 460102
rect 349398 460046 366970 460102
rect 367026 460046 367094 460102
rect 367150 460046 367218 460102
rect 367274 460046 367342 460102
rect 367398 460046 402970 460102
rect 403026 460046 403094 460102
rect 403150 460046 403218 460102
rect 403274 460046 403342 460102
rect 403398 460046 420970 460102
rect 421026 460046 421094 460102
rect 421150 460046 421218 460102
rect 421274 460046 421342 460102
rect 421398 460046 438970 460102
rect 439026 460046 439094 460102
rect 439150 460046 439218 460102
rect 439274 460046 439342 460102
rect 439398 460046 456970 460102
rect 457026 460046 457094 460102
rect 457150 460046 457218 460102
rect 457274 460046 457342 460102
rect 457398 460046 492970 460102
rect 493026 460046 493094 460102
rect 493150 460046 493218 460102
rect 493274 460046 493342 460102
rect 493398 460046 510970 460102
rect 511026 460046 511094 460102
rect 511150 460046 511218 460102
rect 511274 460046 511342 460102
rect 511398 460046 528970 460102
rect 529026 460046 529094 460102
rect 529150 460046 529218 460102
rect 529274 460046 529342 460102
rect 529398 460046 546970 460102
rect 547026 460046 547094 460102
rect 547150 460046 547218 460102
rect 547274 460046 547342 460102
rect 547398 460046 568058 460102
rect 568114 460046 568182 460102
rect 568238 460046 574862 460102
rect 574918 460046 574986 460102
rect 575042 460046 581666 460102
rect 581722 460046 581790 460102
rect 581846 460046 588470 460102
rect 588526 460046 588594 460102
rect 588650 460046 597456 460102
rect 597512 460046 597580 460102
rect 597636 460046 597704 460102
rect 597760 460046 597828 460102
rect 597884 460046 597980 460102
rect -1916 459978 597980 460046
rect -1916 459922 -1820 459978
rect -1764 459922 -1696 459978
rect -1640 459922 -1572 459978
rect -1516 459922 -1448 459978
rect -1392 459922 6970 459978
rect 7026 459922 7094 459978
rect 7150 459922 7218 459978
rect 7274 459922 7342 459978
rect 7398 459922 24970 459978
rect 25026 459922 25094 459978
rect 25150 459922 25218 459978
rect 25274 459922 25342 459978
rect 25398 459922 42970 459978
rect 43026 459922 43094 459978
rect 43150 459922 43218 459978
rect 43274 459922 43342 459978
rect 43398 459922 60970 459978
rect 61026 459922 61094 459978
rect 61150 459922 61218 459978
rect 61274 459922 61342 459978
rect 61398 459922 78970 459978
rect 79026 459922 79094 459978
rect 79150 459922 79218 459978
rect 79274 459922 79342 459978
rect 79398 459922 96970 459978
rect 97026 459922 97094 459978
rect 97150 459922 97218 459978
rect 97274 459922 97342 459978
rect 97398 459922 132970 459978
rect 133026 459922 133094 459978
rect 133150 459922 133218 459978
rect 133274 459922 133342 459978
rect 133398 459922 150970 459978
rect 151026 459922 151094 459978
rect 151150 459922 151218 459978
rect 151274 459922 151342 459978
rect 151398 459922 168970 459978
rect 169026 459922 169094 459978
rect 169150 459922 169218 459978
rect 169274 459922 169342 459978
rect 169398 459922 186970 459978
rect 187026 459922 187094 459978
rect 187150 459922 187218 459978
rect 187274 459922 187342 459978
rect 187398 459922 222970 459978
rect 223026 459922 223094 459978
rect 223150 459922 223218 459978
rect 223274 459922 223342 459978
rect 223398 459922 240970 459978
rect 241026 459922 241094 459978
rect 241150 459922 241218 459978
rect 241274 459922 241342 459978
rect 241398 459922 258970 459978
rect 259026 459922 259094 459978
rect 259150 459922 259218 459978
rect 259274 459922 259342 459978
rect 259398 459922 276970 459978
rect 277026 459922 277094 459978
rect 277150 459922 277218 459978
rect 277274 459922 277342 459978
rect 277398 459922 312970 459978
rect 313026 459922 313094 459978
rect 313150 459922 313218 459978
rect 313274 459922 313342 459978
rect 313398 459922 330970 459978
rect 331026 459922 331094 459978
rect 331150 459922 331218 459978
rect 331274 459922 331342 459978
rect 331398 459922 348970 459978
rect 349026 459922 349094 459978
rect 349150 459922 349218 459978
rect 349274 459922 349342 459978
rect 349398 459922 366970 459978
rect 367026 459922 367094 459978
rect 367150 459922 367218 459978
rect 367274 459922 367342 459978
rect 367398 459922 402970 459978
rect 403026 459922 403094 459978
rect 403150 459922 403218 459978
rect 403274 459922 403342 459978
rect 403398 459922 420970 459978
rect 421026 459922 421094 459978
rect 421150 459922 421218 459978
rect 421274 459922 421342 459978
rect 421398 459922 438970 459978
rect 439026 459922 439094 459978
rect 439150 459922 439218 459978
rect 439274 459922 439342 459978
rect 439398 459922 456970 459978
rect 457026 459922 457094 459978
rect 457150 459922 457218 459978
rect 457274 459922 457342 459978
rect 457398 459922 492970 459978
rect 493026 459922 493094 459978
rect 493150 459922 493218 459978
rect 493274 459922 493342 459978
rect 493398 459922 510970 459978
rect 511026 459922 511094 459978
rect 511150 459922 511218 459978
rect 511274 459922 511342 459978
rect 511398 459922 528970 459978
rect 529026 459922 529094 459978
rect 529150 459922 529218 459978
rect 529274 459922 529342 459978
rect 529398 459922 546970 459978
rect 547026 459922 547094 459978
rect 547150 459922 547218 459978
rect 547274 459922 547342 459978
rect 547398 459922 568058 459978
rect 568114 459922 568182 459978
rect 568238 459922 574862 459978
rect 574918 459922 574986 459978
rect 575042 459922 581666 459978
rect 581722 459922 581790 459978
rect 581846 459922 588470 459978
rect 588526 459922 588594 459978
rect 588650 459922 597456 459978
rect 597512 459922 597580 459978
rect 597636 459922 597704 459978
rect 597760 459922 597828 459978
rect 597884 459922 597980 459978
rect -1916 459826 597980 459922
rect -1916 454350 597980 454446
rect -1916 454294 -860 454350
rect -804 454294 -736 454350
rect -680 454294 -612 454350
rect -556 454294 -488 454350
rect -432 454294 3250 454350
rect 3306 454294 3374 454350
rect 3430 454294 3498 454350
rect 3554 454294 3622 454350
rect 3678 454294 21250 454350
rect 21306 454294 21374 454350
rect 21430 454294 21498 454350
rect 21554 454294 21622 454350
rect 21678 454294 39250 454350
rect 39306 454294 39374 454350
rect 39430 454294 39498 454350
rect 39554 454294 39622 454350
rect 39678 454294 57250 454350
rect 57306 454294 57374 454350
rect 57430 454294 57498 454350
rect 57554 454294 57622 454350
rect 57678 454294 93250 454350
rect 93306 454294 93374 454350
rect 93430 454294 93498 454350
rect 93554 454294 93622 454350
rect 93678 454294 111250 454350
rect 111306 454294 111374 454350
rect 111430 454294 111498 454350
rect 111554 454294 111622 454350
rect 111678 454294 129250 454350
rect 129306 454294 129374 454350
rect 129430 454294 129498 454350
rect 129554 454294 129622 454350
rect 129678 454294 147250 454350
rect 147306 454294 147374 454350
rect 147430 454294 147498 454350
rect 147554 454294 147622 454350
rect 147678 454294 183250 454350
rect 183306 454294 183374 454350
rect 183430 454294 183498 454350
rect 183554 454294 183622 454350
rect 183678 454294 201250 454350
rect 201306 454294 201374 454350
rect 201430 454294 201498 454350
rect 201554 454294 201622 454350
rect 201678 454294 219250 454350
rect 219306 454294 219374 454350
rect 219430 454294 219498 454350
rect 219554 454294 219622 454350
rect 219678 454294 237250 454350
rect 237306 454294 237374 454350
rect 237430 454294 237498 454350
rect 237554 454294 237622 454350
rect 237678 454294 273250 454350
rect 273306 454294 273374 454350
rect 273430 454294 273498 454350
rect 273554 454294 273622 454350
rect 273678 454294 291250 454350
rect 291306 454294 291374 454350
rect 291430 454294 291498 454350
rect 291554 454294 291622 454350
rect 291678 454294 309250 454350
rect 309306 454294 309374 454350
rect 309430 454294 309498 454350
rect 309554 454294 309622 454350
rect 309678 454294 327250 454350
rect 327306 454294 327374 454350
rect 327430 454294 327498 454350
rect 327554 454294 327622 454350
rect 327678 454294 363250 454350
rect 363306 454294 363374 454350
rect 363430 454294 363498 454350
rect 363554 454294 363622 454350
rect 363678 454294 381250 454350
rect 381306 454294 381374 454350
rect 381430 454294 381498 454350
rect 381554 454294 381622 454350
rect 381678 454294 399250 454350
rect 399306 454294 399374 454350
rect 399430 454294 399498 454350
rect 399554 454294 399622 454350
rect 399678 454294 417250 454350
rect 417306 454294 417374 454350
rect 417430 454294 417498 454350
rect 417554 454294 417622 454350
rect 417678 454294 453250 454350
rect 453306 454294 453374 454350
rect 453430 454294 453498 454350
rect 453554 454294 453622 454350
rect 453678 454294 471250 454350
rect 471306 454294 471374 454350
rect 471430 454294 471498 454350
rect 471554 454294 471622 454350
rect 471678 454294 489250 454350
rect 489306 454294 489374 454350
rect 489430 454294 489498 454350
rect 489554 454294 489622 454350
rect 489678 454294 507250 454350
rect 507306 454294 507374 454350
rect 507430 454294 507498 454350
rect 507554 454294 507622 454350
rect 507678 454294 543250 454350
rect 543306 454294 543374 454350
rect 543430 454294 543498 454350
rect 543554 454294 543622 454350
rect 543678 454294 564656 454350
rect 564712 454294 564780 454350
rect 564836 454294 571460 454350
rect 571516 454294 571584 454350
rect 571640 454294 578264 454350
rect 578320 454294 578388 454350
rect 578444 454294 585068 454350
rect 585124 454294 585192 454350
rect 585248 454294 596496 454350
rect 596552 454294 596620 454350
rect 596676 454294 596744 454350
rect 596800 454294 596868 454350
rect 596924 454294 597980 454350
rect -1916 454226 597980 454294
rect -1916 454170 -860 454226
rect -804 454170 -736 454226
rect -680 454170 -612 454226
rect -556 454170 -488 454226
rect -432 454170 3250 454226
rect 3306 454170 3374 454226
rect 3430 454170 3498 454226
rect 3554 454170 3622 454226
rect 3678 454170 21250 454226
rect 21306 454170 21374 454226
rect 21430 454170 21498 454226
rect 21554 454170 21622 454226
rect 21678 454170 39250 454226
rect 39306 454170 39374 454226
rect 39430 454170 39498 454226
rect 39554 454170 39622 454226
rect 39678 454170 57250 454226
rect 57306 454170 57374 454226
rect 57430 454170 57498 454226
rect 57554 454170 57622 454226
rect 57678 454170 93250 454226
rect 93306 454170 93374 454226
rect 93430 454170 93498 454226
rect 93554 454170 93622 454226
rect 93678 454170 111250 454226
rect 111306 454170 111374 454226
rect 111430 454170 111498 454226
rect 111554 454170 111622 454226
rect 111678 454170 129250 454226
rect 129306 454170 129374 454226
rect 129430 454170 129498 454226
rect 129554 454170 129622 454226
rect 129678 454170 147250 454226
rect 147306 454170 147374 454226
rect 147430 454170 147498 454226
rect 147554 454170 147622 454226
rect 147678 454170 183250 454226
rect 183306 454170 183374 454226
rect 183430 454170 183498 454226
rect 183554 454170 183622 454226
rect 183678 454170 201250 454226
rect 201306 454170 201374 454226
rect 201430 454170 201498 454226
rect 201554 454170 201622 454226
rect 201678 454170 219250 454226
rect 219306 454170 219374 454226
rect 219430 454170 219498 454226
rect 219554 454170 219622 454226
rect 219678 454170 237250 454226
rect 237306 454170 237374 454226
rect 237430 454170 237498 454226
rect 237554 454170 237622 454226
rect 237678 454170 273250 454226
rect 273306 454170 273374 454226
rect 273430 454170 273498 454226
rect 273554 454170 273622 454226
rect 273678 454170 291250 454226
rect 291306 454170 291374 454226
rect 291430 454170 291498 454226
rect 291554 454170 291622 454226
rect 291678 454170 309250 454226
rect 309306 454170 309374 454226
rect 309430 454170 309498 454226
rect 309554 454170 309622 454226
rect 309678 454170 327250 454226
rect 327306 454170 327374 454226
rect 327430 454170 327498 454226
rect 327554 454170 327622 454226
rect 327678 454170 363250 454226
rect 363306 454170 363374 454226
rect 363430 454170 363498 454226
rect 363554 454170 363622 454226
rect 363678 454170 381250 454226
rect 381306 454170 381374 454226
rect 381430 454170 381498 454226
rect 381554 454170 381622 454226
rect 381678 454170 399250 454226
rect 399306 454170 399374 454226
rect 399430 454170 399498 454226
rect 399554 454170 399622 454226
rect 399678 454170 417250 454226
rect 417306 454170 417374 454226
rect 417430 454170 417498 454226
rect 417554 454170 417622 454226
rect 417678 454170 453250 454226
rect 453306 454170 453374 454226
rect 453430 454170 453498 454226
rect 453554 454170 453622 454226
rect 453678 454170 471250 454226
rect 471306 454170 471374 454226
rect 471430 454170 471498 454226
rect 471554 454170 471622 454226
rect 471678 454170 489250 454226
rect 489306 454170 489374 454226
rect 489430 454170 489498 454226
rect 489554 454170 489622 454226
rect 489678 454170 507250 454226
rect 507306 454170 507374 454226
rect 507430 454170 507498 454226
rect 507554 454170 507622 454226
rect 507678 454170 543250 454226
rect 543306 454170 543374 454226
rect 543430 454170 543498 454226
rect 543554 454170 543622 454226
rect 543678 454170 564656 454226
rect 564712 454170 564780 454226
rect 564836 454170 571460 454226
rect 571516 454170 571584 454226
rect 571640 454170 578264 454226
rect 578320 454170 578388 454226
rect 578444 454170 585068 454226
rect 585124 454170 585192 454226
rect 585248 454170 596496 454226
rect 596552 454170 596620 454226
rect 596676 454170 596744 454226
rect 596800 454170 596868 454226
rect 596924 454170 597980 454226
rect -1916 454102 597980 454170
rect -1916 454046 -860 454102
rect -804 454046 -736 454102
rect -680 454046 -612 454102
rect -556 454046 -488 454102
rect -432 454046 3250 454102
rect 3306 454046 3374 454102
rect 3430 454046 3498 454102
rect 3554 454046 3622 454102
rect 3678 454046 21250 454102
rect 21306 454046 21374 454102
rect 21430 454046 21498 454102
rect 21554 454046 21622 454102
rect 21678 454046 39250 454102
rect 39306 454046 39374 454102
rect 39430 454046 39498 454102
rect 39554 454046 39622 454102
rect 39678 454046 57250 454102
rect 57306 454046 57374 454102
rect 57430 454046 57498 454102
rect 57554 454046 57622 454102
rect 57678 454046 93250 454102
rect 93306 454046 93374 454102
rect 93430 454046 93498 454102
rect 93554 454046 93622 454102
rect 93678 454046 111250 454102
rect 111306 454046 111374 454102
rect 111430 454046 111498 454102
rect 111554 454046 111622 454102
rect 111678 454046 129250 454102
rect 129306 454046 129374 454102
rect 129430 454046 129498 454102
rect 129554 454046 129622 454102
rect 129678 454046 147250 454102
rect 147306 454046 147374 454102
rect 147430 454046 147498 454102
rect 147554 454046 147622 454102
rect 147678 454046 183250 454102
rect 183306 454046 183374 454102
rect 183430 454046 183498 454102
rect 183554 454046 183622 454102
rect 183678 454046 201250 454102
rect 201306 454046 201374 454102
rect 201430 454046 201498 454102
rect 201554 454046 201622 454102
rect 201678 454046 219250 454102
rect 219306 454046 219374 454102
rect 219430 454046 219498 454102
rect 219554 454046 219622 454102
rect 219678 454046 237250 454102
rect 237306 454046 237374 454102
rect 237430 454046 237498 454102
rect 237554 454046 237622 454102
rect 237678 454046 273250 454102
rect 273306 454046 273374 454102
rect 273430 454046 273498 454102
rect 273554 454046 273622 454102
rect 273678 454046 291250 454102
rect 291306 454046 291374 454102
rect 291430 454046 291498 454102
rect 291554 454046 291622 454102
rect 291678 454046 309250 454102
rect 309306 454046 309374 454102
rect 309430 454046 309498 454102
rect 309554 454046 309622 454102
rect 309678 454046 327250 454102
rect 327306 454046 327374 454102
rect 327430 454046 327498 454102
rect 327554 454046 327622 454102
rect 327678 454046 363250 454102
rect 363306 454046 363374 454102
rect 363430 454046 363498 454102
rect 363554 454046 363622 454102
rect 363678 454046 381250 454102
rect 381306 454046 381374 454102
rect 381430 454046 381498 454102
rect 381554 454046 381622 454102
rect 381678 454046 399250 454102
rect 399306 454046 399374 454102
rect 399430 454046 399498 454102
rect 399554 454046 399622 454102
rect 399678 454046 417250 454102
rect 417306 454046 417374 454102
rect 417430 454046 417498 454102
rect 417554 454046 417622 454102
rect 417678 454046 453250 454102
rect 453306 454046 453374 454102
rect 453430 454046 453498 454102
rect 453554 454046 453622 454102
rect 453678 454046 471250 454102
rect 471306 454046 471374 454102
rect 471430 454046 471498 454102
rect 471554 454046 471622 454102
rect 471678 454046 489250 454102
rect 489306 454046 489374 454102
rect 489430 454046 489498 454102
rect 489554 454046 489622 454102
rect 489678 454046 507250 454102
rect 507306 454046 507374 454102
rect 507430 454046 507498 454102
rect 507554 454046 507622 454102
rect 507678 454046 543250 454102
rect 543306 454046 543374 454102
rect 543430 454046 543498 454102
rect 543554 454046 543622 454102
rect 543678 454046 564656 454102
rect 564712 454046 564780 454102
rect 564836 454046 571460 454102
rect 571516 454046 571584 454102
rect 571640 454046 578264 454102
rect 578320 454046 578388 454102
rect 578444 454046 585068 454102
rect 585124 454046 585192 454102
rect 585248 454046 596496 454102
rect 596552 454046 596620 454102
rect 596676 454046 596744 454102
rect 596800 454046 596868 454102
rect 596924 454046 597980 454102
rect -1916 453978 597980 454046
rect -1916 453922 -860 453978
rect -804 453922 -736 453978
rect -680 453922 -612 453978
rect -556 453922 -488 453978
rect -432 453922 3250 453978
rect 3306 453922 3374 453978
rect 3430 453922 3498 453978
rect 3554 453922 3622 453978
rect 3678 453922 21250 453978
rect 21306 453922 21374 453978
rect 21430 453922 21498 453978
rect 21554 453922 21622 453978
rect 21678 453922 39250 453978
rect 39306 453922 39374 453978
rect 39430 453922 39498 453978
rect 39554 453922 39622 453978
rect 39678 453922 57250 453978
rect 57306 453922 57374 453978
rect 57430 453922 57498 453978
rect 57554 453922 57622 453978
rect 57678 453922 93250 453978
rect 93306 453922 93374 453978
rect 93430 453922 93498 453978
rect 93554 453922 93622 453978
rect 93678 453922 111250 453978
rect 111306 453922 111374 453978
rect 111430 453922 111498 453978
rect 111554 453922 111622 453978
rect 111678 453922 129250 453978
rect 129306 453922 129374 453978
rect 129430 453922 129498 453978
rect 129554 453922 129622 453978
rect 129678 453922 147250 453978
rect 147306 453922 147374 453978
rect 147430 453922 147498 453978
rect 147554 453922 147622 453978
rect 147678 453922 183250 453978
rect 183306 453922 183374 453978
rect 183430 453922 183498 453978
rect 183554 453922 183622 453978
rect 183678 453922 201250 453978
rect 201306 453922 201374 453978
rect 201430 453922 201498 453978
rect 201554 453922 201622 453978
rect 201678 453922 219250 453978
rect 219306 453922 219374 453978
rect 219430 453922 219498 453978
rect 219554 453922 219622 453978
rect 219678 453922 237250 453978
rect 237306 453922 237374 453978
rect 237430 453922 237498 453978
rect 237554 453922 237622 453978
rect 237678 453922 273250 453978
rect 273306 453922 273374 453978
rect 273430 453922 273498 453978
rect 273554 453922 273622 453978
rect 273678 453922 291250 453978
rect 291306 453922 291374 453978
rect 291430 453922 291498 453978
rect 291554 453922 291622 453978
rect 291678 453922 309250 453978
rect 309306 453922 309374 453978
rect 309430 453922 309498 453978
rect 309554 453922 309622 453978
rect 309678 453922 327250 453978
rect 327306 453922 327374 453978
rect 327430 453922 327498 453978
rect 327554 453922 327622 453978
rect 327678 453922 363250 453978
rect 363306 453922 363374 453978
rect 363430 453922 363498 453978
rect 363554 453922 363622 453978
rect 363678 453922 381250 453978
rect 381306 453922 381374 453978
rect 381430 453922 381498 453978
rect 381554 453922 381622 453978
rect 381678 453922 399250 453978
rect 399306 453922 399374 453978
rect 399430 453922 399498 453978
rect 399554 453922 399622 453978
rect 399678 453922 417250 453978
rect 417306 453922 417374 453978
rect 417430 453922 417498 453978
rect 417554 453922 417622 453978
rect 417678 453922 453250 453978
rect 453306 453922 453374 453978
rect 453430 453922 453498 453978
rect 453554 453922 453622 453978
rect 453678 453922 471250 453978
rect 471306 453922 471374 453978
rect 471430 453922 471498 453978
rect 471554 453922 471622 453978
rect 471678 453922 489250 453978
rect 489306 453922 489374 453978
rect 489430 453922 489498 453978
rect 489554 453922 489622 453978
rect 489678 453922 507250 453978
rect 507306 453922 507374 453978
rect 507430 453922 507498 453978
rect 507554 453922 507622 453978
rect 507678 453922 543250 453978
rect 543306 453922 543374 453978
rect 543430 453922 543498 453978
rect 543554 453922 543622 453978
rect 543678 453922 564656 453978
rect 564712 453922 564780 453978
rect 564836 453922 571460 453978
rect 571516 453922 571584 453978
rect 571640 453922 578264 453978
rect 578320 453922 578388 453978
rect 578444 453922 585068 453978
rect 585124 453922 585192 453978
rect 585248 453922 596496 453978
rect 596552 453922 596620 453978
rect 596676 453922 596744 453978
rect 596800 453922 596868 453978
rect 596924 453922 597980 453978
rect -1916 453826 597980 453922
rect -1916 442350 597980 442446
rect -1916 442294 -1820 442350
rect -1764 442294 -1696 442350
rect -1640 442294 -1572 442350
rect -1516 442294 -1448 442350
rect -1392 442294 6970 442350
rect 7026 442294 7094 442350
rect 7150 442294 7218 442350
rect 7274 442294 7342 442350
rect 7398 442294 24970 442350
rect 25026 442294 25094 442350
rect 25150 442294 25218 442350
rect 25274 442294 25342 442350
rect 25398 442294 42970 442350
rect 43026 442294 43094 442350
rect 43150 442294 43218 442350
rect 43274 442294 43342 442350
rect 43398 442294 60970 442350
rect 61026 442294 61094 442350
rect 61150 442294 61218 442350
rect 61274 442294 61342 442350
rect 61398 442294 78970 442350
rect 79026 442294 79094 442350
rect 79150 442294 79218 442350
rect 79274 442294 79342 442350
rect 79398 442294 96970 442350
rect 97026 442294 97094 442350
rect 97150 442294 97218 442350
rect 97274 442294 97342 442350
rect 97398 442294 132970 442350
rect 133026 442294 133094 442350
rect 133150 442294 133218 442350
rect 133274 442294 133342 442350
rect 133398 442294 150970 442350
rect 151026 442294 151094 442350
rect 151150 442294 151218 442350
rect 151274 442294 151342 442350
rect 151398 442294 168970 442350
rect 169026 442294 169094 442350
rect 169150 442294 169218 442350
rect 169274 442294 169342 442350
rect 169398 442294 186970 442350
rect 187026 442294 187094 442350
rect 187150 442294 187218 442350
rect 187274 442294 187342 442350
rect 187398 442294 222970 442350
rect 223026 442294 223094 442350
rect 223150 442294 223218 442350
rect 223274 442294 223342 442350
rect 223398 442294 240970 442350
rect 241026 442294 241094 442350
rect 241150 442294 241218 442350
rect 241274 442294 241342 442350
rect 241398 442294 258970 442350
rect 259026 442294 259094 442350
rect 259150 442294 259218 442350
rect 259274 442294 259342 442350
rect 259398 442294 276970 442350
rect 277026 442294 277094 442350
rect 277150 442294 277218 442350
rect 277274 442294 277342 442350
rect 277398 442294 312970 442350
rect 313026 442294 313094 442350
rect 313150 442294 313218 442350
rect 313274 442294 313342 442350
rect 313398 442294 330970 442350
rect 331026 442294 331094 442350
rect 331150 442294 331218 442350
rect 331274 442294 331342 442350
rect 331398 442294 348970 442350
rect 349026 442294 349094 442350
rect 349150 442294 349218 442350
rect 349274 442294 349342 442350
rect 349398 442294 366970 442350
rect 367026 442294 367094 442350
rect 367150 442294 367218 442350
rect 367274 442294 367342 442350
rect 367398 442294 402970 442350
rect 403026 442294 403094 442350
rect 403150 442294 403218 442350
rect 403274 442294 403342 442350
rect 403398 442294 420970 442350
rect 421026 442294 421094 442350
rect 421150 442294 421218 442350
rect 421274 442294 421342 442350
rect 421398 442294 438970 442350
rect 439026 442294 439094 442350
rect 439150 442294 439218 442350
rect 439274 442294 439342 442350
rect 439398 442294 456970 442350
rect 457026 442294 457094 442350
rect 457150 442294 457218 442350
rect 457274 442294 457342 442350
rect 457398 442294 492970 442350
rect 493026 442294 493094 442350
rect 493150 442294 493218 442350
rect 493274 442294 493342 442350
rect 493398 442294 510970 442350
rect 511026 442294 511094 442350
rect 511150 442294 511218 442350
rect 511274 442294 511342 442350
rect 511398 442294 528970 442350
rect 529026 442294 529094 442350
rect 529150 442294 529218 442350
rect 529274 442294 529342 442350
rect 529398 442294 546970 442350
rect 547026 442294 547094 442350
rect 547150 442294 547218 442350
rect 547274 442294 547342 442350
rect 547398 442294 568058 442350
rect 568114 442294 568182 442350
rect 568238 442294 574862 442350
rect 574918 442294 574986 442350
rect 575042 442294 581666 442350
rect 581722 442294 581790 442350
rect 581846 442294 588470 442350
rect 588526 442294 588594 442350
rect 588650 442294 597456 442350
rect 597512 442294 597580 442350
rect 597636 442294 597704 442350
rect 597760 442294 597828 442350
rect 597884 442294 597980 442350
rect -1916 442226 597980 442294
rect -1916 442170 -1820 442226
rect -1764 442170 -1696 442226
rect -1640 442170 -1572 442226
rect -1516 442170 -1448 442226
rect -1392 442170 6970 442226
rect 7026 442170 7094 442226
rect 7150 442170 7218 442226
rect 7274 442170 7342 442226
rect 7398 442170 24970 442226
rect 25026 442170 25094 442226
rect 25150 442170 25218 442226
rect 25274 442170 25342 442226
rect 25398 442170 42970 442226
rect 43026 442170 43094 442226
rect 43150 442170 43218 442226
rect 43274 442170 43342 442226
rect 43398 442170 60970 442226
rect 61026 442170 61094 442226
rect 61150 442170 61218 442226
rect 61274 442170 61342 442226
rect 61398 442170 78970 442226
rect 79026 442170 79094 442226
rect 79150 442170 79218 442226
rect 79274 442170 79342 442226
rect 79398 442170 96970 442226
rect 97026 442170 97094 442226
rect 97150 442170 97218 442226
rect 97274 442170 97342 442226
rect 97398 442170 132970 442226
rect 133026 442170 133094 442226
rect 133150 442170 133218 442226
rect 133274 442170 133342 442226
rect 133398 442170 150970 442226
rect 151026 442170 151094 442226
rect 151150 442170 151218 442226
rect 151274 442170 151342 442226
rect 151398 442170 168970 442226
rect 169026 442170 169094 442226
rect 169150 442170 169218 442226
rect 169274 442170 169342 442226
rect 169398 442170 186970 442226
rect 187026 442170 187094 442226
rect 187150 442170 187218 442226
rect 187274 442170 187342 442226
rect 187398 442170 222970 442226
rect 223026 442170 223094 442226
rect 223150 442170 223218 442226
rect 223274 442170 223342 442226
rect 223398 442170 240970 442226
rect 241026 442170 241094 442226
rect 241150 442170 241218 442226
rect 241274 442170 241342 442226
rect 241398 442170 258970 442226
rect 259026 442170 259094 442226
rect 259150 442170 259218 442226
rect 259274 442170 259342 442226
rect 259398 442170 276970 442226
rect 277026 442170 277094 442226
rect 277150 442170 277218 442226
rect 277274 442170 277342 442226
rect 277398 442170 312970 442226
rect 313026 442170 313094 442226
rect 313150 442170 313218 442226
rect 313274 442170 313342 442226
rect 313398 442170 330970 442226
rect 331026 442170 331094 442226
rect 331150 442170 331218 442226
rect 331274 442170 331342 442226
rect 331398 442170 348970 442226
rect 349026 442170 349094 442226
rect 349150 442170 349218 442226
rect 349274 442170 349342 442226
rect 349398 442170 366970 442226
rect 367026 442170 367094 442226
rect 367150 442170 367218 442226
rect 367274 442170 367342 442226
rect 367398 442170 402970 442226
rect 403026 442170 403094 442226
rect 403150 442170 403218 442226
rect 403274 442170 403342 442226
rect 403398 442170 420970 442226
rect 421026 442170 421094 442226
rect 421150 442170 421218 442226
rect 421274 442170 421342 442226
rect 421398 442170 438970 442226
rect 439026 442170 439094 442226
rect 439150 442170 439218 442226
rect 439274 442170 439342 442226
rect 439398 442170 456970 442226
rect 457026 442170 457094 442226
rect 457150 442170 457218 442226
rect 457274 442170 457342 442226
rect 457398 442170 492970 442226
rect 493026 442170 493094 442226
rect 493150 442170 493218 442226
rect 493274 442170 493342 442226
rect 493398 442170 510970 442226
rect 511026 442170 511094 442226
rect 511150 442170 511218 442226
rect 511274 442170 511342 442226
rect 511398 442170 528970 442226
rect 529026 442170 529094 442226
rect 529150 442170 529218 442226
rect 529274 442170 529342 442226
rect 529398 442170 546970 442226
rect 547026 442170 547094 442226
rect 547150 442170 547218 442226
rect 547274 442170 547342 442226
rect 547398 442170 568058 442226
rect 568114 442170 568182 442226
rect 568238 442170 574862 442226
rect 574918 442170 574986 442226
rect 575042 442170 581666 442226
rect 581722 442170 581790 442226
rect 581846 442170 588470 442226
rect 588526 442170 588594 442226
rect 588650 442170 597456 442226
rect 597512 442170 597580 442226
rect 597636 442170 597704 442226
rect 597760 442170 597828 442226
rect 597884 442170 597980 442226
rect -1916 442102 597980 442170
rect -1916 442046 -1820 442102
rect -1764 442046 -1696 442102
rect -1640 442046 -1572 442102
rect -1516 442046 -1448 442102
rect -1392 442046 6970 442102
rect 7026 442046 7094 442102
rect 7150 442046 7218 442102
rect 7274 442046 7342 442102
rect 7398 442046 24970 442102
rect 25026 442046 25094 442102
rect 25150 442046 25218 442102
rect 25274 442046 25342 442102
rect 25398 442046 42970 442102
rect 43026 442046 43094 442102
rect 43150 442046 43218 442102
rect 43274 442046 43342 442102
rect 43398 442046 60970 442102
rect 61026 442046 61094 442102
rect 61150 442046 61218 442102
rect 61274 442046 61342 442102
rect 61398 442046 78970 442102
rect 79026 442046 79094 442102
rect 79150 442046 79218 442102
rect 79274 442046 79342 442102
rect 79398 442046 96970 442102
rect 97026 442046 97094 442102
rect 97150 442046 97218 442102
rect 97274 442046 97342 442102
rect 97398 442046 132970 442102
rect 133026 442046 133094 442102
rect 133150 442046 133218 442102
rect 133274 442046 133342 442102
rect 133398 442046 150970 442102
rect 151026 442046 151094 442102
rect 151150 442046 151218 442102
rect 151274 442046 151342 442102
rect 151398 442046 168970 442102
rect 169026 442046 169094 442102
rect 169150 442046 169218 442102
rect 169274 442046 169342 442102
rect 169398 442046 186970 442102
rect 187026 442046 187094 442102
rect 187150 442046 187218 442102
rect 187274 442046 187342 442102
rect 187398 442046 222970 442102
rect 223026 442046 223094 442102
rect 223150 442046 223218 442102
rect 223274 442046 223342 442102
rect 223398 442046 240970 442102
rect 241026 442046 241094 442102
rect 241150 442046 241218 442102
rect 241274 442046 241342 442102
rect 241398 442046 258970 442102
rect 259026 442046 259094 442102
rect 259150 442046 259218 442102
rect 259274 442046 259342 442102
rect 259398 442046 276970 442102
rect 277026 442046 277094 442102
rect 277150 442046 277218 442102
rect 277274 442046 277342 442102
rect 277398 442046 312970 442102
rect 313026 442046 313094 442102
rect 313150 442046 313218 442102
rect 313274 442046 313342 442102
rect 313398 442046 330970 442102
rect 331026 442046 331094 442102
rect 331150 442046 331218 442102
rect 331274 442046 331342 442102
rect 331398 442046 348970 442102
rect 349026 442046 349094 442102
rect 349150 442046 349218 442102
rect 349274 442046 349342 442102
rect 349398 442046 366970 442102
rect 367026 442046 367094 442102
rect 367150 442046 367218 442102
rect 367274 442046 367342 442102
rect 367398 442046 402970 442102
rect 403026 442046 403094 442102
rect 403150 442046 403218 442102
rect 403274 442046 403342 442102
rect 403398 442046 420970 442102
rect 421026 442046 421094 442102
rect 421150 442046 421218 442102
rect 421274 442046 421342 442102
rect 421398 442046 438970 442102
rect 439026 442046 439094 442102
rect 439150 442046 439218 442102
rect 439274 442046 439342 442102
rect 439398 442046 456970 442102
rect 457026 442046 457094 442102
rect 457150 442046 457218 442102
rect 457274 442046 457342 442102
rect 457398 442046 492970 442102
rect 493026 442046 493094 442102
rect 493150 442046 493218 442102
rect 493274 442046 493342 442102
rect 493398 442046 510970 442102
rect 511026 442046 511094 442102
rect 511150 442046 511218 442102
rect 511274 442046 511342 442102
rect 511398 442046 528970 442102
rect 529026 442046 529094 442102
rect 529150 442046 529218 442102
rect 529274 442046 529342 442102
rect 529398 442046 546970 442102
rect 547026 442046 547094 442102
rect 547150 442046 547218 442102
rect 547274 442046 547342 442102
rect 547398 442046 568058 442102
rect 568114 442046 568182 442102
rect 568238 442046 574862 442102
rect 574918 442046 574986 442102
rect 575042 442046 581666 442102
rect 581722 442046 581790 442102
rect 581846 442046 588470 442102
rect 588526 442046 588594 442102
rect 588650 442046 597456 442102
rect 597512 442046 597580 442102
rect 597636 442046 597704 442102
rect 597760 442046 597828 442102
rect 597884 442046 597980 442102
rect -1916 441978 597980 442046
rect -1916 441922 -1820 441978
rect -1764 441922 -1696 441978
rect -1640 441922 -1572 441978
rect -1516 441922 -1448 441978
rect -1392 441922 6970 441978
rect 7026 441922 7094 441978
rect 7150 441922 7218 441978
rect 7274 441922 7342 441978
rect 7398 441922 24970 441978
rect 25026 441922 25094 441978
rect 25150 441922 25218 441978
rect 25274 441922 25342 441978
rect 25398 441922 42970 441978
rect 43026 441922 43094 441978
rect 43150 441922 43218 441978
rect 43274 441922 43342 441978
rect 43398 441922 60970 441978
rect 61026 441922 61094 441978
rect 61150 441922 61218 441978
rect 61274 441922 61342 441978
rect 61398 441922 78970 441978
rect 79026 441922 79094 441978
rect 79150 441922 79218 441978
rect 79274 441922 79342 441978
rect 79398 441922 96970 441978
rect 97026 441922 97094 441978
rect 97150 441922 97218 441978
rect 97274 441922 97342 441978
rect 97398 441922 132970 441978
rect 133026 441922 133094 441978
rect 133150 441922 133218 441978
rect 133274 441922 133342 441978
rect 133398 441922 150970 441978
rect 151026 441922 151094 441978
rect 151150 441922 151218 441978
rect 151274 441922 151342 441978
rect 151398 441922 168970 441978
rect 169026 441922 169094 441978
rect 169150 441922 169218 441978
rect 169274 441922 169342 441978
rect 169398 441922 186970 441978
rect 187026 441922 187094 441978
rect 187150 441922 187218 441978
rect 187274 441922 187342 441978
rect 187398 441922 222970 441978
rect 223026 441922 223094 441978
rect 223150 441922 223218 441978
rect 223274 441922 223342 441978
rect 223398 441922 240970 441978
rect 241026 441922 241094 441978
rect 241150 441922 241218 441978
rect 241274 441922 241342 441978
rect 241398 441922 258970 441978
rect 259026 441922 259094 441978
rect 259150 441922 259218 441978
rect 259274 441922 259342 441978
rect 259398 441922 276970 441978
rect 277026 441922 277094 441978
rect 277150 441922 277218 441978
rect 277274 441922 277342 441978
rect 277398 441922 312970 441978
rect 313026 441922 313094 441978
rect 313150 441922 313218 441978
rect 313274 441922 313342 441978
rect 313398 441922 330970 441978
rect 331026 441922 331094 441978
rect 331150 441922 331218 441978
rect 331274 441922 331342 441978
rect 331398 441922 348970 441978
rect 349026 441922 349094 441978
rect 349150 441922 349218 441978
rect 349274 441922 349342 441978
rect 349398 441922 366970 441978
rect 367026 441922 367094 441978
rect 367150 441922 367218 441978
rect 367274 441922 367342 441978
rect 367398 441922 402970 441978
rect 403026 441922 403094 441978
rect 403150 441922 403218 441978
rect 403274 441922 403342 441978
rect 403398 441922 420970 441978
rect 421026 441922 421094 441978
rect 421150 441922 421218 441978
rect 421274 441922 421342 441978
rect 421398 441922 438970 441978
rect 439026 441922 439094 441978
rect 439150 441922 439218 441978
rect 439274 441922 439342 441978
rect 439398 441922 456970 441978
rect 457026 441922 457094 441978
rect 457150 441922 457218 441978
rect 457274 441922 457342 441978
rect 457398 441922 492970 441978
rect 493026 441922 493094 441978
rect 493150 441922 493218 441978
rect 493274 441922 493342 441978
rect 493398 441922 510970 441978
rect 511026 441922 511094 441978
rect 511150 441922 511218 441978
rect 511274 441922 511342 441978
rect 511398 441922 528970 441978
rect 529026 441922 529094 441978
rect 529150 441922 529218 441978
rect 529274 441922 529342 441978
rect 529398 441922 546970 441978
rect 547026 441922 547094 441978
rect 547150 441922 547218 441978
rect 547274 441922 547342 441978
rect 547398 441922 568058 441978
rect 568114 441922 568182 441978
rect 568238 441922 574862 441978
rect 574918 441922 574986 441978
rect 575042 441922 581666 441978
rect 581722 441922 581790 441978
rect 581846 441922 588470 441978
rect 588526 441922 588594 441978
rect 588650 441922 597456 441978
rect 597512 441922 597580 441978
rect 597636 441922 597704 441978
rect 597760 441922 597828 441978
rect 597884 441922 597980 441978
rect -1916 441826 597980 441922
rect -1916 436350 597980 436446
rect -1916 436294 -860 436350
rect -804 436294 -736 436350
rect -680 436294 -612 436350
rect -556 436294 -488 436350
rect -432 436294 3250 436350
rect 3306 436294 3374 436350
rect 3430 436294 3498 436350
rect 3554 436294 3622 436350
rect 3678 436294 21250 436350
rect 21306 436294 21374 436350
rect 21430 436294 21498 436350
rect 21554 436294 21622 436350
rect 21678 436294 39250 436350
rect 39306 436294 39374 436350
rect 39430 436294 39498 436350
rect 39554 436294 39622 436350
rect 39678 436294 57250 436350
rect 57306 436294 57374 436350
rect 57430 436294 57498 436350
rect 57554 436294 57622 436350
rect 57678 436294 93250 436350
rect 93306 436294 93374 436350
rect 93430 436294 93498 436350
rect 93554 436294 93622 436350
rect 93678 436294 111250 436350
rect 111306 436294 111374 436350
rect 111430 436294 111498 436350
rect 111554 436294 111622 436350
rect 111678 436294 129250 436350
rect 129306 436294 129374 436350
rect 129430 436294 129498 436350
rect 129554 436294 129622 436350
rect 129678 436294 147250 436350
rect 147306 436294 147374 436350
rect 147430 436294 147498 436350
rect 147554 436294 147622 436350
rect 147678 436294 183250 436350
rect 183306 436294 183374 436350
rect 183430 436294 183498 436350
rect 183554 436294 183622 436350
rect 183678 436294 201250 436350
rect 201306 436294 201374 436350
rect 201430 436294 201498 436350
rect 201554 436294 201622 436350
rect 201678 436294 219250 436350
rect 219306 436294 219374 436350
rect 219430 436294 219498 436350
rect 219554 436294 219622 436350
rect 219678 436294 237250 436350
rect 237306 436294 237374 436350
rect 237430 436294 237498 436350
rect 237554 436294 237622 436350
rect 237678 436294 273250 436350
rect 273306 436294 273374 436350
rect 273430 436294 273498 436350
rect 273554 436294 273622 436350
rect 273678 436294 291250 436350
rect 291306 436294 291374 436350
rect 291430 436294 291498 436350
rect 291554 436294 291622 436350
rect 291678 436294 309250 436350
rect 309306 436294 309374 436350
rect 309430 436294 309498 436350
rect 309554 436294 309622 436350
rect 309678 436294 327250 436350
rect 327306 436294 327374 436350
rect 327430 436294 327498 436350
rect 327554 436294 327622 436350
rect 327678 436294 363250 436350
rect 363306 436294 363374 436350
rect 363430 436294 363498 436350
rect 363554 436294 363622 436350
rect 363678 436294 381250 436350
rect 381306 436294 381374 436350
rect 381430 436294 381498 436350
rect 381554 436294 381622 436350
rect 381678 436294 399250 436350
rect 399306 436294 399374 436350
rect 399430 436294 399498 436350
rect 399554 436294 399622 436350
rect 399678 436294 417250 436350
rect 417306 436294 417374 436350
rect 417430 436294 417498 436350
rect 417554 436294 417622 436350
rect 417678 436294 453250 436350
rect 453306 436294 453374 436350
rect 453430 436294 453498 436350
rect 453554 436294 453622 436350
rect 453678 436294 471250 436350
rect 471306 436294 471374 436350
rect 471430 436294 471498 436350
rect 471554 436294 471622 436350
rect 471678 436294 489250 436350
rect 489306 436294 489374 436350
rect 489430 436294 489498 436350
rect 489554 436294 489622 436350
rect 489678 436294 507250 436350
rect 507306 436294 507374 436350
rect 507430 436294 507498 436350
rect 507554 436294 507622 436350
rect 507678 436294 543250 436350
rect 543306 436294 543374 436350
rect 543430 436294 543498 436350
rect 543554 436294 543622 436350
rect 543678 436294 564656 436350
rect 564712 436294 564780 436350
rect 564836 436294 571460 436350
rect 571516 436294 571584 436350
rect 571640 436294 578264 436350
rect 578320 436294 578388 436350
rect 578444 436294 585068 436350
rect 585124 436294 585192 436350
rect 585248 436294 596496 436350
rect 596552 436294 596620 436350
rect 596676 436294 596744 436350
rect 596800 436294 596868 436350
rect 596924 436294 597980 436350
rect -1916 436226 597980 436294
rect -1916 436170 -860 436226
rect -804 436170 -736 436226
rect -680 436170 -612 436226
rect -556 436170 -488 436226
rect -432 436170 3250 436226
rect 3306 436170 3374 436226
rect 3430 436170 3498 436226
rect 3554 436170 3622 436226
rect 3678 436170 21250 436226
rect 21306 436170 21374 436226
rect 21430 436170 21498 436226
rect 21554 436170 21622 436226
rect 21678 436170 39250 436226
rect 39306 436170 39374 436226
rect 39430 436170 39498 436226
rect 39554 436170 39622 436226
rect 39678 436170 57250 436226
rect 57306 436170 57374 436226
rect 57430 436170 57498 436226
rect 57554 436170 57622 436226
rect 57678 436170 93250 436226
rect 93306 436170 93374 436226
rect 93430 436170 93498 436226
rect 93554 436170 93622 436226
rect 93678 436170 111250 436226
rect 111306 436170 111374 436226
rect 111430 436170 111498 436226
rect 111554 436170 111622 436226
rect 111678 436170 129250 436226
rect 129306 436170 129374 436226
rect 129430 436170 129498 436226
rect 129554 436170 129622 436226
rect 129678 436170 147250 436226
rect 147306 436170 147374 436226
rect 147430 436170 147498 436226
rect 147554 436170 147622 436226
rect 147678 436170 183250 436226
rect 183306 436170 183374 436226
rect 183430 436170 183498 436226
rect 183554 436170 183622 436226
rect 183678 436170 201250 436226
rect 201306 436170 201374 436226
rect 201430 436170 201498 436226
rect 201554 436170 201622 436226
rect 201678 436170 219250 436226
rect 219306 436170 219374 436226
rect 219430 436170 219498 436226
rect 219554 436170 219622 436226
rect 219678 436170 237250 436226
rect 237306 436170 237374 436226
rect 237430 436170 237498 436226
rect 237554 436170 237622 436226
rect 237678 436170 273250 436226
rect 273306 436170 273374 436226
rect 273430 436170 273498 436226
rect 273554 436170 273622 436226
rect 273678 436170 291250 436226
rect 291306 436170 291374 436226
rect 291430 436170 291498 436226
rect 291554 436170 291622 436226
rect 291678 436170 309250 436226
rect 309306 436170 309374 436226
rect 309430 436170 309498 436226
rect 309554 436170 309622 436226
rect 309678 436170 327250 436226
rect 327306 436170 327374 436226
rect 327430 436170 327498 436226
rect 327554 436170 327622 436226
rect 327678 436170 363250 436226
rect 363306 436170 363374 436226
rect 363430 436170 363498 436226
rect 363554 436170 363622 436226
rect 363678 436170 381250 436226
rect 381306 436170 381374 436226
rect 381430 436170 381498 436226
rect 381554 436170 381622 436226
rect 381678 436170 399250 436226
rect 399306 436170 399374 436226
rect 399430 436170 399498 436226
rect 399554 436170 399622 436226
rect 399678 436170 417250 436226
rect 417306 436170 417374 436226
rect 417430 436170 417498 436226
rect 417554 436170 417622 436226
rect 417678 436170 453250 436226
rect 453306 436170 453374 436226
rect 453430 436170 453498 436226
rect 453554 436170 453622 436226
rect 453678 436170 471250 436226
rect 471306 436170 471374 436226
rect 471430 436170 471498 436226
rect 471554 436170 471622 436226
rect 471678 436170 489250 436226
rect 489306 436170 489374 436226
rect 489430 436170 489498 436226
rect 489554 436170 489622 436226
rect 489678 436170 507250 436226
rect 507306 436170 507374 436226
rect 507430 436170 507498 436226
rect 507554 436170 507622 436226
rect 507678 436170 543250 436226
rect 543306 436170 543374 436226
rect 543430 436170 543498 436226
rect 543554 436170 543622 436226
rect 543678 436170 564656 436226
rect 564712 436170 564780 436226
rect 564836 436170 571460 436226
rect 571516 436170 571584 436226
rect 571640 436170 578264 436226
rect 578320 436170 578388 436226
rect 578444 436170 585068 436226
rect 585124 436170 585192 436226
rect 585248 436170 596496 436226
rect 596552 436170 596620 436226
rect 596676 436170 596744 436226
rect 596800 436170 596868 436226
rect 596924 436170 597980 436226
rect -1916 436102 597980 436170
rect -1916 436046 -860 436102
rect -804 436046 -736 436102
rect -680 436046 -612 436102
rect -556 436046 -488 436102
rect -432 436046 3250 436102
rect 3306 436046 3374 436102
rect 3430 436046 3498 436102
rect 3554 436046 3622 436102
rect 3678 436046 21250 436102
rect 21306 436046 21374 436102
rect 21430 436046 21498 436102
rect 21554 436046 21622 436102
rect 21678 436046 39250 436102
rect 39306 436046 39374 436102
rect 39430 436046 39498 436102
rect 39554 436046 39622 436102
rect 39678 436046 57250 436102
rect 57306 436046 57374 436102
rect 57430 436046 57498 436102
rect 57554 436046 57622 436102
rect 57678 436046 93250 436102
rect 93306 436046 93374 436102
rect 93430 436046 93498 436102
rect 93554 436046 93622 436102
rect 93678 436046 111250 436102
rect 111306 436046 111374 436102
rect 111430 436046 111498 436102
rect 111554 436046 111622 436102
rect 111678 436046 129250 436102
rect 129306 436046 129374 436102
rect 129430 436046 129498 436102
rect 129554 436046 129622 436102
rect 129678 436046 147250 436102
rect 147306 436046 147374 436102
rect 147430 436046 147498 436102
rect 147554 436046 147622 436102
rect 147678 436046 183250 436102
rect 183306 436046 183374 436102
rect 183430 436046 183498 436102
rect 183554 436046 183622 436102
rect 183678 436046 201250 436102
rect 201306 436046 201374 436102
rect 201430 436046 201498 436102
rect 201554 436046 201622 436102
rect 201678 436046 219250 436102
rect 219306 436046 219374 436102
rect 219430 436046 219498 436102
rect 219554 436046 219622 436102
rect 219678 436046 237250 436102
rect 237306 436046 237374 436102
rect 237430 436046 237498 436102
rect 237554 436046 237622 436102
rect 237678 436046 273250 436102
rect 273306 436046 273374 436102
rect 273430 436046 273498 436102
rect 273554 436046 273622 436102
rect 273678 436046 291250 436102
rect 291306 436046 291374 436102
rect 291430 436046 291498 436102
rect 291554 436046 291622 436102
rect 291678 436046 309250 436102
rect 309306 436046 309374 436102
rect 309430 436046 309498 436102
rect 309554 436046 309622 436102
rect 309678 436046 327250 436102
rect 327306 436046 327374 436102
rect 327430 436046 327498 436102
rect 327554 436046 327622 436102
rect 327678 436046 363250 436102
rect 363306 436046 363374 436102
rect 363430 436046 363498 436102
rect 363554 436046 363622 436102
rect 363678 436046 381250 436102
rect 381306 436046 381374 436102
rect 381430 436046 381498 436102
rect 381554 436046 381622 436102
rect 381678 436046 399250 436102
rect 399306 436046 399374 436102
rect 399430 436046 399498 436102
rect 399554 436046 399622 436102
rect 399678 436046 417250 436102
rect 417306 436046 417374 436102
rect 417430 436046 417498 436102
rect 417554 436046 417622 436102
rect 417678 436046 453250 436102
rect 453306 436046 453374 436102
rect 453430 436046 453498 436102
rect 453554 436046 453622 436102
rect 453678 436046 471250 436102
rect 471306 436046 471374 436102
rect 471430 436046 471498 436102
rect 471554 436046 471622 436102
rect 471678 436046 489250 436102
rect 489306 436046 489374 436102
rect 489430 436046 489498 436102
rect 489554 436046 489622 436102
rect 489678 436046 507250 436102
rect 507306 436046 507374 436102
rect 507430 436046 507498 436102
rect 507554 436046 507622 436102
rect 507678 436046 543250 436102
rect 543306 436046 543374 436102
rect 543430 436046 543498 436102
rect 543554 436046 543622 436102
rect 543678 436046 564656 436102
rect 564712 436046 564780 436102
rect 564836 436046 571460 436102
rect 571516 436046 571584 436102
rect 571640 436046 578264 436102
rect 578320 436046 578388 436102
rect 578444 436046 585068 436102
rect 585124 436046 585192 436102
rect 585248 436046 596496 436102
rect 596552 436046 596620 436102
rect 596676 436046 596744 436102
rect 596800 436046 596868 436102
rect 596924 436046 597980 436102
rect -1916 435978 597980 436046
rect -1916 435922 -860 435978
rect -804 435922 -736 435978
rect -680 435922 -612 435978
rect -556 435922 -488 435978
rect -432 435922 3250 435978
rect 3306 435922 3374 435978
rect 3430 435922 3498 435978
rect 3554 435922 3622 435978
rect 3678 435922 21250 435978
rect 21306 435922 21374 435978
rect 21430 435922 21498 435978
rect 21554 435922 21622 435978
rect 21678 435922 39250 435978
rect 39306 435922 39374 435978
rect 39430 435922 39498 435978
rect 39554 435922 39622 435978
rect 39678 435922 57250 435978
rect 57306 435922 57374 435978
rect 57430 435922 57498 435978
rect 57554 435922 57622 435978
rect 57678 435922 93250 435978
rect 93306 435922 93374 435978
rect 93430 435922 93498 435978
rect 93554 435922 93622 435978
rect 93678 435922 111250 435978
rect 111306 435922 111374 435978
rect 111430 435922 111498 435978
rect 111554 435922 111622 435978
rect 111678 435922 129250 435978
rect 129306 435922 129374 435978
rect 129430 435922 129498 435978
rect 129554 435922 129622 435978
rect 129678 435922 147250 435978
rect 147306 435922 147374 435978
rect 147430 435922 147498 435978
rect 147554 435922 147622 435978
rect 147678 435922 183250 435978
rect 183306 435922 183374 435978
rect 183430 435922 183498 435978
rect 183554 435922 183622 435978
rect 183678 435922 201250 435978
rect 201306 435922 201374 435978
rect 201430 435922 201498 435978
rect 201554 435922 201622 435978
rect 201678 435922 219250 435978
rect 219306 435922 219374 435978
rect 219430 435922 219498 435978
rect 219554 435922 219622 435978
rect 219678 435922 237250 435978
rect 237306 435922 237374 435978
rect 237430 435922 237498 435978
rect 237554 435922 237622 435978
rect 237678 435922 273250 435978
rect 273306 435922 273374 435978
rect 273430 435922 273498 435978
rect 273554 435922 273622 435978
rect 273678 435922 291250 435978
rect 291306 435922 291374 435978
rect 291430 435922 291498 435978
rect 291554 435922 291622 435978
rect 291678 435922 309250 435978
rect 309306 435922 309374 435978
rect 309430 435922 309498 435978
rect 309554 435922 309622 435978
rect 309678 435922 327250 435978
rect 327306 435922 327374 435978
rect 327430 435922 327498 435978
rect 327554 435922 327622 435978
rect 327678 435922 363250 435978
rect 363306 435922 363374 435978
rect 363430 435922 363498 435978
rect 363554 435922 363622 435978
rect 363678 435922 381250 435978
rect 381306 435922 381374 435978
rect 381430 435922 381498 435978
rect 381554 435922 381622 435978
rect 381678 435922 399250 435978
rect 399306 435922 399374 435978
rect 399430 435922 399498 435978
rect 399554 435922 399622 435978
rect 399678 435922 417250 435978
rect 417306 435922 417374 435978
rect 417430 435922 417498 435978
rect 417554 435922 417622 435978
rect 417678 435922 453250 435978
rect 453306 435922 453374 435978
rect 453430 435922 453498 435978
rect 453554 435922 453622 435978
rect 453678 435922 471250 435978
rect 471306 435922 471374 435978
rect 471430 435922 471498 435978
rect 471554 435922 471622 435978
rect 471678 435922 489250 435978
rect 489306 435922 489374 435978
rect 489430 435922 489498 435978
rect 489554 435922 489622 435978
rect 489678 435922 507250 435978
rect 507306 435922 507374 435978
rect 507430 435922 507498 435978
rect 507554 435922 507622 435978
rect 507678 435922 543250 435978
rect 543306 435922 543374 435978
rect 543430 435922 543498 435978
rect 543554 435922 543622 435978
rect 543678 435922 564656 435978
rect 564712 435922 564780 435978
rect 564836 435922 571460 435978
rect 571516 435922 571584 435978
rect 571640 435922 578264 435978
rect 578320 435922 578388 435978
rect 578444 435922 585068 435978
rect 585124 435922 585192 435978
rect 585248 435922 596496 435978
rect 596552 435922 596620 435978
rect 596676 435922 596744 435978
rect 596800 435922 596868 435978
rect 596924 435922 597980 435978
rect -1916 435826 597980 435922
rect -1916 424350 597980 424446
rect -1916 424294 -1820 424350
rect -1764 424294 -1696 424350
rect -1640 424294 -1572 424350
rect -1516 424294 -1448 424350
rect -1392 424294 6970 424350
rect 7026 424294 7094 424350
rect 7150 424294 7218 424350
rect 7274 424294 7342 424350
rect 7398 424294 24970 424350
rect 25026 424294 25094 424350
rect 25150 424294 25218 424350
rect 25274 424294 25342 424350
rect 25398 424294 42970 424350
rect 43026 424294 43094 424350
rect 43150 424294 43218 424350
rect 43274 424294 43342 424350
rect 43398 424294 60970 424350
rect 61026 424294 61094 424350
rect 61150 424294 61218 424350
rect 61274 424294 61342 424350
rect 61398 424294 78970 424350
rect 79026 424294 79094 424350
rect 79150 424294 79218 424350
rect 79274 424294 79342 424350
rect 79398 424294 96970 424350
rect 97026 424294 97094 424350
rect 97150 424294 97218 424350
rect 97274 424294 97342 424350
rect 97398 424294 132970 424350
rect 133026 424294 133094 424350
rect 133150 424294 133218 424350
rect 133274 424294 133342 424350
rect 133398 424294 150970 424350
rect 151026 424294 151094 424350
rect 151150 424294 151218 424350
rect 151274 424294 151342 424350
rect 151398 424294 168970 424350
rect 169026 424294 169094 424350
rect 169150 424294 169218 424350
rect 169274 424294 169342 424350
rect 169398 424294 186970 424350
rect 187026 424294 187094 424350
rect 187150 424294 187218 424350
rect 187274 424294 187342 424350
rect 187398 424294 222970 424350
rect 223026 424294 223094 424350
rect 223150 424294 223218 424350
rect 223274 424294 223342 424350
rect 223398 424294 240970 424350
rect 241026 424294 241094 424350
rect 241150 424294 241218 424350
rect 241274 424294 241342 424350
rect 241398 424294 258970 424350
rect 259026 424294 259094 424350
rect 259150 424294 259218 424350
rect 259274 424294 259342 424350
rect 259398 424294 276970 424350
rect 277026 424294 277094 424350
rect 277150 424294 277218 424350
rect 277274 424294 277342 424350
rect 277398 424294 312970 424350
rect 313026 424294 313094 424350
rect 313150 424294 313218 424350
rect 313274 424294 313342 424350
rect 313398 424294 330970 424350
rect 331026 424294 331094 424350
rect 331150 424294 331218 424350
rect 331274 424294 331342 424350
rect 331398 424294 348970 424350
rect 349026 424294 349094 424350
rect 349150 424294 349218 424350
rect 349274 424294 349342 424350
rect 349398 424294 366970 424350
rect 367026 424294 367094 424350
rect 367150 424294 367218 424350
rect 367274 424294 367342 424350
rect 367398 424294 402970 424350
rect 403026 424294 403094 424350
rect 403150 424294 403218 424350
rect 403274 424294 403342 424350
rect 403398 424294 420970 424350
rect 421026 424294 421094 424350
rect 421150 424294 421218 424350
rect 421274 424294 421342 424350
rect 421398 424294 438970 424350
rect 439026 424294 439094 424350
rect 439150 424294 439218 424350
rect 439274 424294 439342 424350
rect 439398 424294 456970 424350
rect 457026 424294 457094 424350
rect 457150 424294 457218 424350
rect 457274 424294 457342 424350
rect 457398 424294 492970 424350
rect 493026 424294 493094 424350
rect 493150 424294 493218 424350
rect 493274 424294 493342 424350
rect 493398 424294 510970 424350
rect 511026 424294 511094 424350
rect 511150 424294 511218 424350
rect 511274 424294 511342 424350
rect 511398 424294 528970 424350
rect 529026 424294 529094 424350
rect 529150 424294 529218 424350
rect 529274 424294 529342 424350
rect 529398 424294 546970 424350
rect 547026 424294 547094 424350
rect 547150 424294 547218 424350
rect 547274 424294 547342 424350
rect 547398 424294 568058 424350
rect 568114 424294 568182 424350
rect 568238 424294 574862 424350
rect 574918 424294 574986 424350
rect 575042 424294 581666 424350
rect 581722 424294 581790 424350
rect 581846 424294 588470 424350
rect 588526 424294 588594 424350
rect 588650 424294 597456 424350
rect 597512 424294 597580 424350
rect 597636 424294 597704 424350
rect 597760 424294 597828 424350
rect 597884 424294 597980 424350
rect -1916 424226 597980 424294
rect -1916 424170 -1820 424226
rect -1764 424170 -1696 424226
rect -1640 424170 -1572 424226
rect -1516 424170 -1448 424226
rect -1392 424170 6970 424226
rect 7026 424170 7094 424226
rect 7150 424170 7218 424226
rect 7274 424170 7342 424226
rect 7398 424170 24970 424226
rect 25026 424170 25094 424226
rect 25150 424170 25218 424226
rect 25274 424170 25342 424226
rect 25398 424170 42970 424226
rect 43026 424170 43094 424226
rect 43150 424170 43218 424226
rect 43274 424170 43342 424226
rect 43398 424170 60970 424226
rect 61026 424170 61094 424226
rect 61150 424170 61218 424226
rect 61274 424170 61342 424226
rect 61398 424170 78970 424226
rect 79026 424170 79094 424226
rect 79150 424170 79218 424226
rect 79274 424170 79342 424226
rect 79398 424170 96970 424226
rect 97026 424170 97094 424226
rect 97150 424170 97218 424226
rect 97274 424170 97342 424226
rect 97398 424170 132970 424226
rect 133026 424170 133094 424226
rect 133150 424170 133218 424226
rect 133274 424170 133342 424226
rect 133398 424170 150970 424226
rect 151026 424170 151094 424226
rect 151150 424170 151218 424226
rect 151274 424170 151342 424226
rect 151398 424170 168970 424226
rect 169026 424170 169094 424226
rect 169150 424170 169218 424226
rect 169274 424170 169342 424226
rect 169398 424170 186970 424226
rect 187026 424170 187094 424226
rect 187150 424170 187218 424226
rect 187274 424170 187342 424226
rect 187398 424170 222970 424226
rect 223026 424170 223094 424226
rect 223150 424170 223218 424226
rect 223274 424170 223342 424226
rect 223398 424170 240970 424226
rect 241026 424170 241094 424226
rect 241150 424170 241218 424226
rect 241274 424170 241342 424226
rect 241398 424170 258970 424226
rect 259026 424170 259094 424226
rect 259150 424170 259218 424226
rect 259274 424170 259342 424226
rect 259398 424170 276970 424226
rect 277026 424170 277094 424226
rect 277150 424170 277218 424226
rect 277274 424170 277342 424226
rect 277398 424170 312970 424226
rect 313026 424170 313094 424226
rect 313150 424170 313218 424226
rect 313274 424170 313342 424226
rect 313398 424170 330970 424226
rect 331026 424170 331094 424226
rect 331150 424170 331218 424226
rect 331274 424170 331342 424226
rect 331398 424170 348970 424226
rect 349026 424170 349094 424226
rect 349150 424170 349218 424226
rect 349274 424170 349342 424226
rect 349398 424170 366970 424226
rect 367026 424170 367094 424226
rect 367150 424170 367218 424226
rect 367274 424170 367342 424226
rect 367398 424170 402970 424226
rect 403026 424170 403094 424226
rect 403150 424170 403218 424226
rect 403274 424170 403342 424226
rect 403398 424170 420970 424226
rect 421026 424170 421094 424226
rect 421150 424170 421218 424226
rect 421274 424170 421342 424226
rect 421398 424170 438970 424226
rect 439026 424170 439094 424226
rect 439150 424170 439218 424226
rect 439274 424170 439342 424226
rect 439398 424170 456970 424226
rect 457026 424170 457094 424226
rect 457150 424170 457218 424226
rect 457274 424170 457342 424226
rect 457398 424170 492970 424226
rect 493026 424170 493094 424226
rect 493150 424170 493218 424226
rect 493274 424170 493342 424226
rect 493398 424170 510970 424226
rect 511026 424170 511094 424226
rect 511150 424170 511218 424226
rect 511274 424170 511342 424226
rect 511398 424170 528970 424226
rect 529026 424170 529094 424226
rect 529150 424170 529218 424226
rect 529274 424170 529342 424226
rect 529398 424170 546970 424226
rect 547026 424170 547094 424226
rect 547150 424170 547218 424226
rect 547274 424170 547342 424226
rect 547398 424170 568058 424226
rect 568114 424170 568182 424226
rect 568238 424170 574862 424226
rect 574918 424170 574986 424226
rect 575042 424170 581666 424226
rect 581722 424170 581790 424226
rect 581846 424170 588470 424226
rect 588526 424170 588594 424226
rect 588650 424170 597456 424226
rect 597512 424170 597580 424226
rect 597636 424170 597704 424226
rect 597760 424170 597828 424226
rect 597884 424170 597980 424226
rect -1916 424102 597980 424170
rect -1916 424046 -1820 424102
rect -1764 424046 -1696 424102
rect -1640 424046 -1572 424102
rect -1516 424046 -1448 424102
rect -1392 424046 6970 424102
rect 7026 424046 7094 424102
rect 7150 424046 7218 424102
rect 7274 424046 7342 424102
rect 7398 424046 24970 424102
rect 25026 424046 25094 424102
rect 25150 424046 25218 424102
rect 25274 424046 25342 424102
rect 25398 424046 42970 424102
rect 43026 424046 43094 424102
rect 43150 424046 43218 424102
rect 43274 424046 43342 424102
rect 43398 424046 60970 424102
rect 61026 424046 61094 424102
rect 61150 424046 61218 424102
rect 61274 424046 61342 424102
rect 61398 424046 78970 424102
rect 79026 424046 79094 424102
rect 79150 424046 79218 424102
rect 79274 424046 79342 424102
rect 79398 424046 96970 424102
rect 97026 424046 97094 424102
rect 97150 424046 97218 424102
rect 97274 424046 97342 424102
rect 97398 424046 132970 424102
rect 133026 424046 133094 424102
rect 133150 424046 133218 424102
rect 133274 424046 133342 424102
rect 133398 424046 150970 424102
rect 151026 424046 151094 424102
rect 151150 424046 151218 424102
rect 151274 424046 151342 424102
rect 151398 424046 168970 424102
rect 169026 424046 169094 424102
rect 169150 424046 169218 424102
rect 169274 424046 169342 424102
rect 169398 424046 186970 424102
rect 187026 424046 187094 424102
rect 187150 424046 187218 424102
rect 187274 424046 187342 424102
rect 187398 424046 222970 424102
rect 223026 424046 223094 424102
rect 223150 424046 223218 424102
rect 223274 424046 223342 424102
rect 223398 424046 240970 424102
rect 241026 424046 241094 424102
rect 241150 424046 241218 424102
rect 241274 424046 241342 424102
rect 241398 424046 258970 424102
rect 259026 424046 259094 424102
rect 259150 424046 259218 424102
rect 259274 424046 259342 424102
rect 259398 424046 276970 424102
rect 277026 424046 277094 424102
rect 277150 424046 277218 424102
rect 277274 424046 277342 424102
rect 277398 424046 312970 424102
rect 313026 424046 313094 424102
rect 313150 424046 313218 424102
rect 313274 424046 313342 424102
rect 313398 424046 330970 424102
rect 331026 424046 331094 424102
rect 331150 424046 331218 424102
rect 331274 424046 331342 424102
rect 331398 424046 348970 424102
rect 349026 424046 349094 424102
rect 349150 424046 349218 424102
rect 349274 424046 349342 424102
rect 349398 424046 366970 424102
rect 367026 424046 367094 424102
rect 367150 424046 367218 424102
rect 367274 424046 367342 424102
rect 367398 424046 402970 424102
rect 403026 424046 403094 424102
rect 403150 424046 403218 424102
rect 403274 424046 403342 424102
rect 403398 424046 420970 424102
rect 421026 424046 421094 424102
rect 421150 424046 421218 424102
rect 421274 424046 421342 424102
rect 421398 424046 438970 424102
rect 439026 424046 439094 424102
rect 439150 424046 439218 424102
rect 439274 424046 439342 424102
rect 439398 424046 456970 424102
rect 457026 424046 457094 424102
rect 457150 424046 457218 424102
rect 457274 424046 457342 424102
rect 457398 424046 492970 424102
rect 493026 424046 493094 424102
rect 493150 424046 493218 424102
rect 493274 424046 493342 424102
rect 493398 424046 510970 424102
rect 511026 424046 511094 424102
rect 511150 424046 511218 424102
rect 511274 424046 511342 424102
rect 511398 424046 528970 424102
rect 529026 424046 529094 424102
rect 529150 424046 529218 424102
rect 529274 424046 529342 424102
rect 529398 424046 546970 424102
rect 547026 424046 547094 424102
rect 547150 424046 547218 424102
rect 547274 424046 547342 424102
rect 547398 424046 568058 424102
rect 568114 424046 568182 424102
rect 568238 424046 574862 424102
rect 574918 424046 574986 424102
rect 575042 424046 581666 424102
rect 581722 424046 581790 424102
rect 581846 424046 588470 424102
rect 588526 424046 588594 424102
rect 588650 424046 597456 424102
rect 597512 424046 597580 424102
rect 597636 424046 597704 424102
rect 597760 424046 597828 424102
rect 597884 424046 597980 424102
rect -1916 423978 597980 424046
rect -1916 423922 -1820 423978
rect -1764 423922 -1696 423978
rect -1640 423922 -1572 423978
rect -1516 423922 -1448 423978
rect -1392 423922 6970 423978
rect 7026 423922 7094 423978
rect 7150 423922 7218 423978
rect 7274 423922 7342 423978
rect 7398 423922 24970 423978
rect 25026 423922 25094 423978
rect 25150 423922 25218 423978
rect 25274 423922 25342 423978
rect 25398 423922 42970 423978
rect 43026 423922 43094 423978
rect 43150 423922 43218 423978
rect 43274 423922 43342 423978
rect 43398 423922 60970 423978
rect 61026 423922 61094 423978
rect 61150 423922 61218 423978
rect 61274 423922 61342 423978
rect 61398 423922 78970 423978
rect 79026 423922 79094 423978
rect 79150 423922 79218 423978
rect 79274 423922 79342 423978
rect 79398 423922 96970 423978
rect 97026 423922 97094 423978
rect 97150 423922 97218 423978
rect 97274 423922 97342 423978
rect 97398 423922 132970 423978
rect 133026 423922 133094 423978
rect 133150 423922 133218 423978
rect 133274 423922 133342 423978
rect 133398 423922 150970 423978
rect 151026 423922 151094 423978
rect 151150 423922 151218 423978
rect 151274 423922 151342 423978
rect 151398 423922 168970 423978
rect 169026 423922 169094 423978
rect 169150 423922 169218 423978
rect 169274 423922 169342 423978
rect 169398 423922 186970 423978
rect 187026 423922 187094 423978
rect 187150 423922 187218 423978
rect 187274 423922 187342 423978
rect 187398 423922 222970 423978
rect 223026 423922 223094 423978
rect 223150 423922 223218 423978
rect 223274 423922 223342 423978
rect 223398 423922 240970 423978
rect 241026 423922 241094 423978
rect 241150 423922 241218 423978
rect 241274 423922 241342 423978
rect 241398 423922 258970 423978
rect 259026 423922 259094 423978
rect 259150 423922 259218 423978
rect 259274 423922 259342 423978
rect 259398 423922 276970 423978
rect 277026 423922 277094 423978
rect 277150 423922 277218 423978
rect 277274 423922 277342 423978
rect 277398 423922 312970 423978
rect 313026 423922 313094 423978
rect 313150 423922 313218 423978
rect 313274 423922 313342 423978
rect 313398 423922 330970 423978
rect 331026 423922 331094 423978
rect 331150 423922 331218 423978
rect 331274 423922 331342 423978
rect 331398 423922 348970 423978
rect 349026 423922 349094 423978
rect 349150 423922 349218 423978
rect 349274 423922 349342 423978
rect 349398 423922 366970 423978
rect 367026 423922 367094 423978
rect 367150 423922 367218 423978
rect 367274 423922 367342 423978
rect 367398 423922 402970 423978
rect 403026 423922 403094 423978
rect 403150 423922 403218 423978
rect 403274 423922 403342 423978
rect 403398 423922 420970 423978
rect 421026 423922 421094 423978
rect 421150 423922 421218 423978
rect 421274 423922 421342 423978
rect 421398 423922 438970 423978
rect 439026 423922 439094 423978
rect 439150 423922 439218 423978
rect 439274 423922 439342 423978
rect 439398 423922 456970 423978
rect 457026 423922 457094 423978
rect 457150 423922 457218 423978
rect 457274 423922 457342 423978
rect 457398 423922 492970 423978
rect 493026 423922 493094 423978
rect 493150 423922 493218 423978
rect 493274 423922 493342 423978
rect 493398 423922 510970 423978
rect 511026 423922 511094 423978
rect 511150 423922 511218 423978
rect 511274 423922 511342 423978
rect 511398 423922 528970 423978
rect 529026 423922 529094 423978
rect 529150 423922 529218 423978
rect 529274 423922 529342 423978
rect 529398 423922 546970 423978
rect 547026 423922 547094 423978
rect 547150 423922 547218 423978
rect 547274 423922 547342 423978
rect 547398 423922 568058 423978
rect 568114 423922 568182 423978
rect 568238 423922 574862 423978
rect 574918 423922 574986 423978
rect 575042 423922 581666 423978
rect 581722 423922 581790 423978
rect 581846 423922 588470 423978
rect 588526 423922 588594 423978
rect 588650 423922 597456 423978
rect 597512 423922 597580 423978
rect 597636 423922 597704 423978
rect 597760 423922 597828 423978
rect 597884 423922 597980 423978
rect -1916 423826 597980 423922
rect -1916 418350 597980 418446
rect -1916 418294 -860 418350
rect -804 418294 -736 418350
rect -680 418294 -612 418350
rect -556 418294 -488 418350
rect -432 418294 3250 418350
rect 3306 418294 3374 418350
rect 3430 418294 3498 418350
rect 3554 418294 3622 418350
rect 3678 418294 21250 418350
rect 21306 418294 21374 418350
rect 21430 418294 21498 418350
rect 21554 418294 21622 418350
rect 21678 418294 39250 418350
rect 39306 418294 39374 418350
rect 39430 418294 39498 418350
rect 39554 418294 39622 418350
rect 39678 418294 57250 418350
rect 57306 418294 57374 418350
rect 57430 418294 57498 418350
rect 57554 418294 57622 418350
rect 57678 418294 93250 418350
rect 93306 418294 93374 418350
rect 93430 418294 93498 418350
rect 93554 418294 93622 418350
rect 93678 418294 111250 418350
rect 111306 418294 111374 418350
rect 111430 418294 111498 418350
rect 111554 418294 111622 418350
rect 111678 418294 129250 418350
rect 129306 418294 129374 418350
rect 129430 418294 129498 418350
rect 129554 418294 129622 418350
rect 129678 418294 147250 418350
rect 147306 418294 147374 418350
rect 147430 418294 147498 418350
rect 147554 418294 147622 418350
rect 147678 418294 183250 418350
rect 183306 418294 183374 418350
rect 183430 418294 183498 418350
rect 183554 418294 183622 418350
rect 183678 418294 201250 418350
rect 201306 418294 201374 418350
rect 201430 418294 201498 418350
rect 201554 418294 201622 418350
rect 201678 418294 219250 418350
rect 219306 418294 219374 418350
rect 219430 418294 219498 418350
rect 219554 418294 219622 418350
rect 219678 418294 237250 418350
rect 237306 418294 237374 418350
rect 237430 418294 237498 418350
rect 237554 418294 237622 418350
rect 237678 418294 273250 418350
rect 273306 418294 273374 418350
rect 273430 418294 273498 418350
rect 273554 418294 273622 418350
rect 273678 418294 291250 418350
rect 291306 418294 291374 418350
rect 291430 418294 291498 418350
rect 291554 418294 291622 418350
rect 291678 418294 309250 418350
rect 309306 418294 309374 418350
rect 309430 418294 309498 418350
rect 309554 418294 309622 418350
rect 309678 418294 327250 418350
rect 327306 418294 327374 418350
rect 327430 418294 327498 418350
rect 327554 418294 327622 418350
rect 327678 418294 363250 418350
rect 363306 418294 363374 418350
rect 363430 418294 363498 418350
rect 363554 418294 363622 418350
rect 363678 418294 381250 418350
rect 381306 418294 381374 418350
rect 381430 418294 381498 418350
rect 381554 418294 381622 418350
rect 381678 418294 399250 418350
rect 399306 418294 399374 418350
rect 399430 418294 399498 418350
rect 399554 418294 399622 418350
rect 399678 418294 417250 418350
rect 417306 418294 417374 418350
rect 417430 418294 417498 418350
rect 417554 418294 417622 418350
rect 417678 418294 453250 418350
rect 453306 418294 453374 418350
rect 453430 418294 453498 418350
rect 453554 418294 453622 418350
rect 453678 418294 471250 418350
rect 471306 418294 471374 418350
rect 471430 418294 471498 418350
rect 471554 418294 471622 418350
rect 471678 418294 489250 418350
rect 489306 418294 489374 418350
rect 489430 418294 489498 418350
rect 489554 418294 489622 418350
rect 489678 418294 507250 418350
rect 507306 418294 507374 418350
rect 507430 418294 507498 418350
rect 507554 418294 507622 418350
rect 507678 418294 543250 418350
rect 543306 418294 543374 418350
rect 543430 418294 543498 418350
rect 543554 418294 543622 418350
rect 543678 418294 564656 418350
rect 564712 418294 564780 418350
rect 564836 418294 571460 418350
rect 571516 418294 571584 418350
rect 571640 418294 578264 418350
rect 578320 418294 578388 418350
rect 578444 418294 585068 418350
rect 585124 418294 585192 418350
rect 585248 418294 596496 418350
rect 596552 418294 596620 418350
rect 596676 418294 596744 418350
rect 596800 418294 596868 418350
rect 596924 418294 597980 418350
rect -1916 418226 597980 418294
rect -1916 418170 -860 418226
rect -804 418170 -736 418226
rect -680 418170 -612 418226
rect -556 418170 -488 418226
rect -432 418170 3250 418226
rect 3306 418170 3374 418226
rect 3430 418170 3498 418226
rect 3554 418170 3622 418226
rect 3678 418170 21250 418226
rect 21306 418170 21374 418226
rect 21430 418170 21498 418226
rect 21554 418170 21622 418226
rect 21678 418170 39250 418226
rect 39306 418170 39374 418226
rect 39430 418170 39498 418226
rect 39554 418170 39622 418226
rect 39678 418170 57250 418226
rect 57306 418170 57374 418226
rect 57430 418170 57498 418226
rect 57554 418170 57622 418226
rect 57678 418170 93250 418226
rect 93306 418170 93374 418226
rect 93430 418170 93498 418226
rect 93554 418170 93622 418226
rect 93678 418170 111250 418226
rect 111306 418170 111374 418226
rect 111430 418170 111498 418226
rect 111554 418170 111622 418226
rect 111678 418170 129250 418226
rect 129306 418170 129374 418226
rect 129430 418170 129498 418226
rect 129554 418170 129622 418226
rect 129678 418170 147250 418226
rect 147306 418170 147374 418226
rect 147430 418170 147498 418226
rect 147554 418170 147622 418226
rect 147678 418170 183250 418226
rect 183306 418170 183374 418226
rect 183430 418170 183498 418226
rect 183554 418170 183622 418226
rect 183678 418170 201250 418226
rect 201306 418170 201374 418226
rect 201430 418170 201498 418226
rect 201554 418170 201622 418226
rect 201678 418170 219250 418226
rect 219306 418170 219374 418226
rect 219430 418170 219498 418226
rect 219554 418170 219622 418226
rect 219678 418170 237250 418226
rect 237306 418170 237374 418226
rect 237430 418170 237498 418226
rect 237554 418170 237622 418226
rect 237678 418170 273250 418226
rect 273306 418170 273374 418226
rect 273430 418170 273498 418226
rect 273554 418170 273622 418226
rect 273678 418170 291250 418226
rect 291306 418170 291374 418226
rect 291430 418170 291498 418226
rect 291554 418170 291622 418226
rect 291678 418170 309250 418226
rect 309306 418170 309374 418226
rect 309430 418170 309498 418226
rect 309554 418170 309622 418226
rect 309678 418170 327250 418226
rect 327306 418170 327374 418226
rect 327430 418170 327498 418226
rect 327554 418170 327622 418226
rect 327678 418170 363250 418226
rect 363306 418170 363374 418226
rect 363430 418170 363498 418226
rect 363554 418170 363622 418226
rect 363678 418170 381250 418226
rect 381306 418170 381374 418226
rect 381430 418170 381498 418226
rect 381554 418170 381622 418226
rect 381678 418170 399250 418226
rect 399306 418170 399374 418226
rect 399430 418170 399498 418226
rect 399554 418170 399622 418226
rect 399678 418170 417250 418226
rect 417306 418170 417374 418226
rect 417430 418170 417498 418226
rect 417554 418170 417622 418226
rect 417678 418170 453250 418226
rect 453306 418170 453374 418226
rect 453430 418170 453498 418226
rect 453554 418170 453622 418226
rect 453678 418170 471250 418226
rect 471306 418170 471374 418226
rect 471430 418170 471498 418226
rect 471554 418170 471622 418226
rect 471678 418170 489250 418226
rect 489306 418170 489374 418226
rect 489430 418170 489498 418226
rect 489554 418170 489622 418226
rect 489678 418170 507250 418226
rect 507306 418170 507374 418226
rect 507430 418170 507498 418226
rect 507554 418170 507622 418226
rect 507678 418170 543250 418226
rect 543306 418170 543374 418226
rect 543430 418170 543498 418226
rect 543554 418170 543622 418226
rect 543678 418170 564656 418226
rect 564712 418170 564780 418226
rect 564836 418170 571460 418226
rect 571516 418170 571584 418226
rect 571640 418170 578264 418226
rect 578320 418170 578388 418226
rect 578444 418170 585068 418226
rect 585124 418170 585192 418226
rect 585248 418170 596496 418226
rect 596552 418170 596620 418226
rect 596676 418170 596744 418226
rect 596800 418170 596868 418226
rect 596924 418170 597980 418226
rect -1916 418102 597980 418170
rect -1916 418046 -860 418102
rect -804 418046 -736 418102
rect -680 418046 -612 418102
rect -556 418046 -488 418102
rect -432 418046 3250 418102
rect 3306 418046 3374 418102
rect 3430 418046 3498 418102
rect 3554 418046 3622 418102
rect 3678 418046 21250 418102
rect 21306 418046 21374 418102
rect 21430 418046 21498 418102
rect 21554 418046 21622 418102
rect 21678 418046 39250 418102
rect 39306 418046 39374 418102
rect 39430 418046 39498 418102
rect 39554 418046 39622 418102
rect 39678 418046 57250 418102
rect 57306 418046 57374 418102
rect 57430 418046 57498 418102
rect 57554 418046 57622 418102
rect 57678 418046 93250 418102
rect 93306 418046 93374 418102
rect 93430 418046 93498 418102
rect 93554 418046 93622 418102
rect 93678 418046 111250 418102
rect 111306 418046 111374 418102
rect 111430 418046 111498 418102
rect 111554 418046 111622 418102
rect 111678 418046 129250 418102
rect 129306 418046 129374 418102
rect 129430 418046 129498 418102
rect 129554 418046 129622 418102
rect 129678 418046 147250 418102
rect 147306 418046 147374 418102
rect 147430 418046 147498 418102
rect 147554 418046 147622 418102
rect 147678 418046 183250 418102
rect 183306 418046 183374 418102
rect 183430 418046 183498 418102
rect 183554 418046 183622 418102
rect 183678 418046 201250 418102
rect 201306 418046 201374 418102
rect 201430 418046 201498 418102
rect 201554 418046 201622 418102
rect 201678 418046 219250 418102
rect 219306 418046 219374 418102
rect 219430 418046 219498 418102
rect 219554 418046 219622 418102
rect 219678 418046 237250 418102
rect 237306 418046 237374 418102
rect 237430 418046 237498 418102
rect 237554 418046 237622 418102
rect 237678 418046 273250 418102
rect 273306 418046 273374 418102
rect 273430 418046 273498 418102
rect 273554 418046 273622 418102
rect 273678 418046 291250 418102
rect 291306 418046 291374 418102
rect 291430 418046 291498 418102
rect 291554 418046 291622 418102
rect 291678 418046 309250 418102
rect 309306 418046 309374 418102
rect 309430 418046 309498 418102
rect 309554 418046 309622 418102
rect 309678 418046 327250 418102
rect 327306 418046 327374 418102
rect 327430 418046 327498 418102
rect 327554 418046 327622 418102
rect 327678 418046 363250 418102
rect 363306 418046 363374 418102
rect 363430 418046 363498 418102
rect 363554 418046 363622 418102
rect 363678 418046 381250 418102
rect 381306 418046 381374 418102
rect 381430 418046 381498 418102
rect 381554 418046 381622 418102
rect 381678 418046 399250 418102
rect 399306 418046 399374 418102
rect 399430 418046 399498 418102
rect 399554 418046 399622 418102
rect 399678 418046 417250 418102
rect 417306 418046 417374 418102
rect 417430 418046 417498 418102
rect 417554 418046 417622 418102
rect 417678 418046 453250 418102
rect 453306 418046 453374 418102
rect 453430 418046 453498 418102
rect 453554 418046 453622 418102
rect 453678 418046 471250 418102
rect 471306 418046 471374 418102
rect 471430 418046 471498 418102
rect 471554 418046 471622 418102
rect 471678 418046 489250 418102
rect 489306 418046 489374 418102
rect 489430 418046 489498 418102
rect 489554 418046 489622 418102
rect 489678 418046 507250 418102
rect 507306 418046 507374 418102
rect 507430 418046 507498 418102
rect 507554 418046 507622 418102
rect 507678 418046 543250 418102
rect 543306 418046 543374 418102
rect 543430 418046 543498 418102
rect 543554 418046 543622 418102
rect 543678 418046 564656 418102
rect 564712 418046 564780 418102
rect 564836 418046 571460 418102
rect 571516 418046 571584 418102
rect 571640 418046 578264 418102
rect 578320 418046 578388 418102
rect 578444 418046 585068 418102
rect 585124 418046 585192 418102
rect 585248 418046 596496 418102
rect 596552 418046 596620 418102
rect 596676 418046 596744 418102
rect 596800 418046 596868 418102
rect 596924 418046 597980 418102
rect -1916 417978 597980 418046
rect -1916 417922 -860 417978
rect -804 417922 -736 417978
rect -680 417922 -612 417978
rect -556 417922 -488 417978
rect -432 417922 3250 417978
rect 3306 417922 3374 417978
rect 3430 417922 3498 417978
rect 3554 417922 3622 417978
rect 3678 417922 21250 417978
rect 21306 417922 21374 417978
rect 21430 417922 21498 417978
rect 21554 417922 21622 417978
rect 21678 417922 39250 417978
rect 39306 417922 39374 417978
rect 39430 417922 39498 417978
rect 39554 417922 39622 417978
rect 39678 417922 57250 417978
rect 57306 417922 57374 417978
rect 57430 417922 57498 417978
rect 57554 417922 57622 417978
rect 57678 417922 93250 417978
rect 93306 417922 93374 417978
rect 93430 417922 93498 417978
rect 93554 417922 93622 417978
rect 93678 417922 111250 417978
rect 111306 417922 111374 417978
rect 111430 417922 111498 417978
rect 111554 417922 111622 417978
rect 111678 417922 129250 417978
rect 129306 417922 129374 417978
rect 129430 417922 129498 417978
rect 129554 417922 129622 417978
rect 129678 417922 147250 417978
rect 147306 417922 147374 417978
rect 147430 417922 147498 417978
rect 147554 417922 147622 417978
rect 147678 417922 183250 417978
rect 183306 417922 183374 417978
rect 183430 417922 183498 417978
rect 183554 417922 183622 417978
rect 183678 417922 201250 417978
rect 201306 417922 201374 417978
rect 201430 417922 201498 417978
rect 201554 417922 201622 417978
rect 201678 417922 219250 417978
rect 219306 417922 219374 417978
rect 219430 417922 219498 417978
rect 219554 417922 219622 417978
rect 219678 417922 237250 417978
rect 237306 417922 237374 417978
rect 237430 417922 237498 417978
rect 237554 417922 237622 417978
rect 237678 417922 273250 417978
rect 273306 417922 273374 417978
rect 273430 417922 273498 417978
rect 273554 417922 273622 417978
rect 273678 417922 291250 417978
rect 291306 417922 291374 417978
rect 291430 417922 291498 417978
rect 291554 417922 291622 417978
rect 291678 417922 309250 417978
rect 309306 417922 309374 417978
rect 309430 417922 309498 417978
rect 309554 417922 309622 417978
rect 309678 417922 327250 417978
rect 327306 417922 327374 417978
rect 327430 417922 327498 417978
rect 327554 417922 327622 417978
rect 327678 417922 363250 417978
rect 363306 417922 363374 417978
rect 363430 417922 363498 417978
rect 363554 417922 363622 417978
rect 363678 417922 381250 417978
rect 381306 417922 381374 417978
rect 381430 417922 381498 417978
rect 381554 417922 381622 417978
rect 381678 417922 399250 417978
rect 399306 417922 399374 417978
rect 399430 417922 399498 417978
rect 399554 417922 399622 417978
rect 399678 417922 417250 417978
rect 417306 417922 417374 417978
rect 417430 417922 417498 417978
rect 417554 417922 417622 417978
rect 417678 417922 453250 417978
rect 453306 417922 453374 417978
rect 453430 417922 453498 417978
rect 453554 417922 453622 417978
rect 453678 417922 471250 417978
rect 471306 417922 471374 417978
rect 471430 417922 471498 417978
rect 471554 417922 471622 417978
rect 471678 417922 489250 417978
rect 489306 417922 489374 417978
rect 489430 417922 489498 417978
rect 489554 417922 489622 417978
rect 489678 417922 507250 417978
rect 507306 417922 507374 417978
rect 507430 417922 507498 417978
rect 507554 417922 507622 417978
rect 507678 417922 543250 417978
rect 543306 417922 543374 417978
rect 543430 417922 543498 417978
rect 543554 417922 543622 417978
rect 543678 417922 564656 417978
rect 564712 417922 564780 417978
rect 564836 417922 571460 417978
rect 571516 417922 571584 417978
rect 571640 417922 578264 417978
rect 578320 417922 578388 417978
rect 578444 417922 585068 417978
rect 585124 417922 585192 417978
rect 585248 417922 596496 417978
rect 596552 417922 596620 417978
rect 596676 417922 596744 417978
rect 596800 417922 596868 417978
rect 596924 417922 597980 417978
rect -1916 417826 597980 417922
rect -1916 406350 597980 406446
rect -1916 406294 -1820 406350
rect -1764 406294 -1696 406350
rect -1640 406294 -1572 406350
rect -1516 406294 -1448 406350
rect -1392 406294 6970 406350
rect 7026 406294 7094 406350
rect 7150 406294 7218 406350
rect 7274 406294 7342 406350
rect 7398 406294 24970 406350
rect 25026 406294 25094 406350
rect 25150 406294 25218 406350
rect 25274 406294 25342 406350
rect 25398 406294 42970 406350
rect 43026 406294 43094 406350
rect 43150 406294 43218 406350
rect 43274 406294 43342 406350
rect 43398 406294 60970 406350
rect 61026 406294 61094 406350
rect 61150 406294 61218 406350
rect 61274 406294 61342 406350
rect 61398 406294 78970 406350
rect 79026 406294 79094 406350
rect 79150 406294 79218 406350
rect 79274 406294 79342 406350
rect 79398 406294 96970 406350
rect 97026 406294 97094 406350
rect 97150 406294 97218 406350
rect 97274 406294 97342 406350
rect 97398 406294 132970 406350
rect 133026 406294 133094 406350
rect 133150 406294 133218 406350
rect 133274 406294 133342 406350
rect 133398 406294 150970 406350
rect 151026 406294 151094 406350
rect 151150 406294 151218 406350
rect 151274 406294 151342 406350
rect 151398 406294 168970 406350
rect 169026 406294 169094 406350
rect 169150 406294 169218 406350
rect 169274 406294 169342 406350
rect 169398 406294 186970 406350
rect 187026 406294 187094 406350
rect 187150 406294 187218 406350
rect 187274 406294 187342 406350
rect 187398 406294 222970 406350
rect 223026 406294 223094 406350
rect 223150 406294 223218 406350
rect 223274 406294 223342 406350
rect 223398 406294 240970 406350
rect 241026 406294 241094 406350
rect 241150 406294 241218 406350
rect 241274 406294 241342 406350
rect 241398 406294 258970 406350
rect 259026 406294 259094 406350
rect 259150 406294 259218 406350
rect 259274 406294 259342 406350
rect 259398 406294 276970 406350
rect 277026 406294 277094 406350
rect 277150 406294 277218 406350
rect 277274 406294 277342 406350
rect 277398 406294 312970 406350
rect 313026 406294 313094 406350
rect 313150 406294 313218 406350
rect 313274 406294 313342 406350
rect 313398 406294 330970 406350
rect 331026 406294 331094 406350
rect 331150 406294 331218 406350
rect 331274 406294 331342 406350
rect 331398 406294 348970 406350
rect 349026 406294 349094 406350
rect 349150 406294 349218 406350
rect 349274 406294 349342 406350
rect 349398 406294 366970 406350
rect 367026 406294 367094 406350
rect 367150 406294 367218 406350
rect 367274 406294 367342 406350
rect 367398 406294 402970 406350
rect 403026 406294 403094 406350
rect 403150 406294 403218 406350
rect 403274 406294 403342 406350
rect 403398 406294 420970 406350
rect 421026 406294 421094 406350
rect 421150 406294 421218 406350
rect 421274 406294 421342 406350
rect 421398 406294 438970 406350
rect 439026 406294 439094 406350
rect 439150 406294 439218 406350
rect 439274 406294 439342 406350
rect 439398 406294 456970 406350
rect 457026 406294 457094 406350
rect 457150 406294 457218 406350
rect 457274 406294 457342 406350
rect 457398 406294 492970 406350
rect 493026 406294 493094 406350
rect 493150 406294 493218 406350
rect 493274 406294 493342 406350
rect 493398 406294 510970 406350
rect 511026 406294 511094 406350
rect 511150 406294 511218 406350
rect 511274 406294 511342 406350
rect 511398 406294 528970 406350
rect 529026 406294 529094 406350
rect 529150 406294 529218 406350
rect 529274 406294 529342 406350
rect 529398 406294 546970 406350
rect 547026 406294 547094 406350
rect 547150 406294 547218 406350
rect 547274 406294 547342 406350
rect 547398 406294 568058 406350
rect 568114 406294 568182 406350
rect 568238 406294 574862 406350
rect 574918 406294 574986 406350
rect 575042 406294 581666 406350
rect 581722 406294 581790 406350
rect 581846 406294 588470 406350
rect 588526 406294 588594 406350
rect 588650 406294 597456 406350
rect 597512 406294 597580 406350
rect 597636 406294 597704 406350
rect 597760 406294 597828 406350
rect 597884 406294 597980 406350
rect -1916 406226 597980 406294
rect -1916 406170 -1820 406226
rect -1764 406170 -1696 406226
rect -1640 406170 -1572 406226
rect -1516 406170 -1448 406226
rect -1392 406170 6970 406226
rect 7026 406170 7094 406226
rect 7150 406170 7218 406226
rect 7274 406170 7342 406226
rect 7398 406170 24970 406226
rect 25026 406170 25094 406226
rect 25150 406170 25218 406226
rect 25274 406170 25342 406226
rect 25398 406170 42970 406226
rect 43026 406170 43094 406226
rect 43150 406170 43218 406226
rect 43274 406170 43342 406226
rect 43398 406170 60970 406226
rect 61026 406170 61094 406226
rect 61150 406170 61218 406226
rect 61274 406170 61342 406226
rect 61398 406170 78970 406226
rect 79026 406170 79094 406226
rect 79150 406170 79218 406226
rect 79274 406170 79342 406226
rect 79398 406170 96970 406226
rect 97026 406170 97094 406226
rect 97150 406170 97218 406226
rect 97274 406170 97342 406226
rect 97398 406170 132970 406226
rect 133026 406170 133094 406226
rect 133150 406170 133218 406226
rect 133274 406170 133342 406226
rect 133398 406170 150970 406226
rect 151026 406170 151094 406226
rect 151150 406170 151218 406226
rect 151274 406170 151342 406226
rect 151398 406170 168970 406226
rect 169026 406170 169094 406226
rect 169150 406170 169218 406226
rect 169274 406170 169342 406226
rect 169398 406170 186970 406226
rect 187026 406170 187094 406226
rect 187150 406170 187218 406226
rect 187274 406170 187342 406226
rect 187398 406170 222970 406226
rect 223026 406170 223094 406226
rect 223150 406170 223218 406226
rect 223274 406170 223342 406226
rect 223398 406170 240970 406226
rect 241026 406170 241094 406226
rect 241150 406170 241218 406226
rect 241274 406170 241342 406226
rect 241398 406170 258970 406226
rect 259026 406170 259094 406226
rect 259150 406170 259218 406226
rect 259274 406170 259342 406226
rect 259398 406170 276970 406226
rect 277026 406170 277094 406226
rect 277150 406170 277218 406226
rect 277274 406170 277342 406226
rect 277398 406170 312970 406226
rect 313026 406170 313094 406226
rect 313150 406170 313218 406226
rect 313274 406170 313342 406226
rect 313398 406170 330970 406226
rect 331026 406170 331094 406226
rect 331150 406170 331218 406226
rect 331274 406170 331342 406226
rect 331398 406170 348970 406226
rect 349026 406170 349094 406226
rect 349150 406170 349218 406226
rect 349274 406170 349342 406226
rect 349398 406170 366970 406226
rect 367026 406170 367094 406226
rect 367150 406170 367218 406226
rect 367274 406170 367342 406226
rect 367398 406170 402970 406226
rect 403026 406170 403094 406226
rect 403150 406170 403218 406226
rect 403274 406170 403342 406226
rect 403398 406170 420970 406226
rect 421026 406170 421094 406226
rect 421150 406170 421218 406226
rect 421274 406170 421342 406226
rect 421398 406170 438970 406226
rect 439026 406170 439094 406226
rect 439150 406170 439218 406226
rect 439274 406170 439342 406226
rect 439398 406170 456970 406226
rect 457026 406170 457094 406226
rect 457150 406170 457218 406226
rect 457274 406170 457342 406226
rect 457398 406170 492970 406226
rect 493026 406170 493094 406226
rect 493150 406170 493218 406226
rect 493274 406170 493342 406226
rect 493398 406170 510970 406226
rect 511026 406170 511094 406226
rect 511150 406170 511218 406226
rect 511274 406170 511342 406226
rect 511398 406170 528970 406226
rect 529026 406170 529094 406226
rect 529150 406170 529218 406226
rect 529274 406170 529342 406226
rect 529398 406170 546970 406226
rect 547026 406170 547094 406226
rect 547150 406170 547218 406226
rect 547274 406170 547342 406226
rect 547398 406170 568058 406226
rect 568114 406170 568182 406226
rect 568238 406170 574862 406226
rect 574918 406170 574986 406226
rect 575042 406170 581666 406226
rect 581722 406170 581790 406226
rect 581846 406170 588470 406226
rect 588526 406170 588594 406226
rect 588650 406170 597456 406226
rect 597512 406170 597580 406226
rect 597636 406170 597704 406226
rect 597760 406170 597828 406226
rect 597884 406170 597980 406226
rect -1916 406102 597980 406170
rect -1916 406046 -1820 406102
rect -1764 406046 -1696 406102
rect -1640 406046 -1572 406102
rect -1516 406046 -1448 406102
rect -1392 406046 6970 406102
rect 7026 406046 7094 406102
rect 7150 406046 7218 406102
rect 7274 406046 7342 406102
rect 7398 406046 24970 406102
rect 25026 406046 25094 406102
rect 25150 406046 25218 406102
rect 25274 406046 25342 406102
rect 25398 406046 42970 406102
rect 43026 406046 43094 406102
rect 43150 406046 43218 406102
rect 43274 406046 43342 406102
rect 43398 406046 60970 406102
rect 61026 406046 61094 406102
rect 61150 406046 61218 406102
rect 61274 406046 61342 406102
rect 61398 406046 78970 406102
rect 79026 406046 79094 406102
rect 79150 406046 79218 406102
rect 79274 406046 79342 406102
rect 79398 406046 96970 406102
rect 97026 406046 97094 406102
rect 97150 406046 97218 406102
rect 97274 406046 97342 406102
rect 97398 406046 132970 406102
rect 133026 406046 133094 406102
rect 133150 406046 133218 406102
rect 133274 406046 133342 406102
rect 133398 406046 150970 406102
rect 151026 406046 151094 406102
rect 151150 406046 151218 406102
rect 151274 406046 151342 406102
rect 151398 406046 168970 406102
rect 169026 406046 169094 406102
rect 169150 406046 169218 406102
rect 169274 406046 169342 406102
rect 169398 406046 186970 406102
rect 187026 406046 187094 406102
rect 187150 406046 187218 406102
rect 187274 406046 187342 406102
rect 187398 406046 222970 406102
rect 223026 406046 223094 406102
rect 223150 406046 223218 406102
rect 223274 406046 223342 406102
rect 223398 406046 240970 406102
rect 241026 406046 241094 406102
rect 241150 406046 241218 406102
rect 241274 406046 241342 406102
rect 241398 406046 258970 406102
rect 259026 406046 259094 406102
rect 259150 406046 259218 406102
rect 259274 406046 259342 406102
rect 259398 406046 276970 406102
rect 277026 406046 277094 406102
rect 277150 406046 277218 406102
rect 277274 406046 277342 406102
rect 277398 406046 312970 406102
rect 313026 406046 313094 406102
rect 313150 406046 313218 406102
rect 313274 406046 313342 406102
rect 313398 406046 330970 406102
rect 331026 406046 331094 406102
rect 331150 406046 331218 406102
rect 331274 406046 331342 406102
rect 331398 406046 348970 406102
rect 349026 406046 349094 406102
rect 349150 406046 349218 406102
rect 349274 406046 349342 406102
rect 349398 406046 366970 406102
rect 367026 406046 367094 406102
rect 367150 406046 367218 406102
rect 367274 406046 367342 406102
rect 367398 406046 402970 406102
rect 403026 406046 403094 406102
rect 403150 406046 403218 406102
rect 403274 406046 403342 406102
rect 403398 406046 420970 406102
rect 421026 406046 421094 406102
rect 421150 406046 421218 406102
rect 421274 406046 421342 406102
rect 421398 406046 438970 406102
rect 439026 406046 439094 406102
rect 439150 406046 439218 406102
rect 439274 406046 439342 406102
rect 439398 406046 456970 406102
rect 457026 406046 457094 406102
rect 457150 406046 457218 406102
rect 457274 406046 457342 406102
rect 457398 406046 492970 406102
rect 493026 406046 493094 406102
rect 493150 406046 493218 406102
rect 493274 406046 493342 406102
rect 493398 406046 510970 406102
rect 511026 406046 511094 406102
rect 511150 406046 511218 406102
rect 511274 406046 511342 406102
rect 511398 406046 528970 406102
rect 529026 406046 529094 406102
rect 529150 406046 529218 406102
rect 529274 406046 529342 406102
rect 529398 406046 546970 406102
rect 547026 406046 547094 406102
rect 547150 406046 547218 406102
rect 547274 406046 547342 406102
rect 547398 406046 568058 406102
rect 568114 406046 568182 406102
rect 568238 406046 574862 406102
rect 574918 406046 574986 406102
rect 575042 406046 581666 406102
rect 581722 406046 581790 406102
rect 581846 406046 588470 406102
rect 588526 406046 588594 406102
rect 588650 406046 597456 406102
rect 597512 406046 597580 406102
rect 597636 406046 597704 406102
rect 597760 406046 597828 406102
rect 597884 406046 597980 406102
rect -1916 405978 597980 406046
rect -1916 405922 -1820 405978
rect -1764 405922 -1696 405978
rect -1640 405922 -1572 405978
rect -1516 405922 -1448 405978
rect -1392 405922 6970 405978
rect 7026 405922 7094 405978
rect 7150 405922 7218 405978
rect 7274 405922 7342 405978
rect 7398 405922 24970 405978
rect 25026 405922 25094 405978
rect 25150 405922 25218 405978
rect 25274 405922 25342 405978
rect 25398 405922 42970 405978
rect 43026 405922 43094 405978
rect 43150 405922 43218 405978
rect 43274 405922 43342 405978
rect 43398 405922 60970 405978
rect 61026 405922 61094 405978
rect 61150 405922 61218 405978
rect 61274 405922 61342 405978
rect 61398 405922 78970 405978
rect 79026 405922 79094 405978
rect 79150 405922 79218 405978
rect 79274 405922 79342 405978
rect 79398 405922 96970 405978
rect 97026 405922 97094 405978
rect 97150 405922 97218 405978
rect 97274 405922 97342 405978
rect 97398 405922 132970 405978
rect 133026 405922 133094 405978
rect 133150 405922 133218 405978
rect 133274 405922 133342 405978
rect 133398 405922 150970 405978
rect 151026 405922 151094 405978
rect 151150 405922 151218 405978
rect 151274 405922 151342 405978
rect 151398 405922 168970 405978
rect 169026 405922 169094 405978
rect 169150 405922 169218 405978
rect 169274 405922 169342 405978
rect 169398 405922 186970 405978
rect 187026 405922 187094 405978
rect 187150 405922 187218 405978
rect 187274 405922 187342 405978
rect 187398 405922 222970 405978
rect 223026 405922 223094 405978
rect 223150 405922 223218 405978
rect 223274 405922 223342 405978
rect 223398 405922 240970 405978
rect 241026 405922 241094 405978
rect 241150 405922 241218 405978
rect 241274 405922 241342 405978
rect 241398 405922 258970 405978
rect 259026 405922 259094 405978
rect 259150 405922 259218 405978
rect 259274 405922 259342 405978
rect 259398 405922 276970 405978
rect 277026 405922 277094 405978
rect 277150 405922 277218 405978
rect 277274 405922 277342 405978
rect 277398 405922 312970 405978
rect 313026 405922 313094 405978
rect 313150 405922 313218 405978
rect 313274 405922 313342 405978
rect 313398 405922 330970 405978
rect 331026 405922 331094 405978
rect 331150 405922 331218 405978
rect 331274 405922 331342 405978
rect 331398 405922 348970 405978
rect 349026 405922 349094 405978
rect 349150 405922 349218 405978
rect 349274 405922 349342 405978
rect 349398 405922 366970 405978
rect 367026 405922 367094 405978
rect 367150 405922 367218 405978
rect 367274 405922 367342 405978
rect 367398 405922 402970 405978
rect 403026 405922 403094 405978
rect 403150 405922 403218 405978
rect 403274 405922 403342 405978
rect 403398 405922 420970 405978
rect 421026 405922 421094 405978
rect 421150 405922 421218 405978
rect 421274 405922 421342 405978
rect 421398 405922 438970 405978
rect 439026 405922 439094 405978
rect 439150 405922 439218 405978
rect 439274 405922 439342 405978
rect 439398 405922 456970 405978
rect 457026 405922 457094 405978
rect 457150 405922 457218 405978
rect 457274 405922 457342 405978
rect 457398 405922 492970 405978
rect 493026 405922 493094 405978
rect 493150 405922 493218 405978
rect 493274 405922 493342 405978
rect 493398 405922 510970 405978
rect 511026 405922 511094 405978
rect 511150 405922 511218 405978
rect 511274 405922 511342 405978
rect 511398 405922 528970 405978
rect 529026 405922 529094 405978
rect 529150 405922 529218 405978
rect 529274 405922 529342 405978
rect 529398 405922 546970 405978
rect 547026 405922 547094 405978
rect 547150 405922 547218 405978
rect 547274 405922 547342 405978
rect 547398 405922 568058 405978
rect 568114 405922 568182 405978
rect 568238 405922 574862 405978
rect 574918 405922 574986 405978
rect 575042 405922 581666 405978
rect 581722 405922 581790 405978
rect 581846 405922 588470 405978
rect 588526 405922 588594 405978
rect 588650 405922 597456 405978
rect 597512 405922 597580 405978
rect 597636 405922 597704 405978
rect 597760 405922 597828 405978
rect 597884 405922 597980 405978
rect -1916 405826 597980 405922
rect -1916 400350 597980 400446
rect -1916 400294 -860 400350
rect -804 400294 -736 400350
rect -680 400294 -612 400350
rect -556 400294 -488 400350
rect -432 400294 3250 400350
rect 3306 400294 3374 400350
rect 3430 400294 3498 400350
rect 3554 400294 3622 400350
rect 3678 400294 21250 400350
rect 21306 400294 21374 400350
rect 21430 400294 21498 400350
rect 21554 400294 21622 400350
rect 21678 400294 39250 400350
rect 39306 400294 39374 400350
rect 39430 400294 39498 400350
rect 39554 400294 39622 400350
rect 39678 400294 57250 400350
rect 57306 400294 57374 400350
rect 57430 400294 57498 400350
rect 57554 400294 57622 400350
rect 57678 400294 93250 400350
rect 93306 400294 93374 400350
rect 93430 400294 93498 400350
rect 93554 400294 93622 400350
rect 93678 400294 111250 400350
rect 111306 400294 111374 400350
rect 111430 400294 111498 400350
rect 111554 400294 111622 400350
rect 111678 400294 129250 400350
rect 129306 400294 129374 400350
rect 129430 400294 129498 400350
rect 129554 400294 129622 400350
rect 129678 400294 147250 400350
rect 147306 400294 147374 400350
rect 147430 400294 147498 400350
rect 147554 400294 147622 400350
rect 147678 400294 183250 400350
rect 183306 400294 183374 400350
rect 183430 400294 183498 400350
rect 183554 400294 183622 400350
rect 183678 400294 201250 400350
rect 201306 400294 201374 400350
rect 201430 400294 201498 400350
rect 201554 400294 201622 400350
rect 201678 400294 219250 400350
rect 219306 400294 219374 400350
rect 219430 400294 219498 400350
rect 219554 400294 219622 400350
rect 219678 400294 237250 400350
rect 237306 400294 237374 400350
rect 237430 400294 237498 400350
rect 237554 400294 237622 400350
rect 237678 400294 273250 400350
rect 273306 400294 273374 400350
rect 273430 400294 273498 400350
rect 273554 400294 273622 400350
rect 273678 400294 291250 400350
rect 291306 400294 291374 400350
rect 291430 400294 291498 400350
rect 291554 400294 291622 400350
rect 291678 400294 309250 400350
rect 309306 400294 309374 400350
rect 309430 400294 309498 400350
rect 309554 400294 309622 400350
rect 309678 400294 327250 400350
rect 327306 400294 327374 400350
rect 327430 400294 327498 400350
rect 327554 400294 327622 400350
rect 327678 400294 363250 400350
rect 363306 400294 363374 400350
rect 363430 400294 363498 400350
rect 363554 400294 363622 400350
rect 363678 400294 381250 400350
rect 381306 400294 381374 400350
rect 381430 400294 381498 400350
rect 381554 400294 381622 400350
rect 381678 400294 399250 400350
rect 399306 400294 399374 400350
rect 399430 400294 399498 400350
rect 399554 400294 399622 400350
rect 399678 400294 417250 400350
rect 417306 400294 417374 400350
rect 417430 400294 417498 400350
rect 417554 400294 417622 400350
rect 417678 400294 453250 400350
rect 453306 400294 453374 400350
rect 453430 400294 453498 400350
rect 453554 400294 453622 400350
rect 453678 400294 471250 400350
rect 471306 400294 471374 400350
rect 471430 400294 471498 400350
rect 471554 400294 471622 400350
rect 471678 400294 489250 400350
rect 489306 400294 489374 400350
rect 489430 400294 489498 400350
rect 489554 400294 489622 400350
rect 489678 400294 507250 400350
rect 507306 400294 507374 400350
rect 507430 400294 507498 400350
rect 507554 400294 507622 400350
rect 507678 400294 543250 400350
rect 543306 400294 543374 400350
rect 543430 400294 543498 400350
rect 543554 400294 543622 400350
rect 543678 400294 564656 400350
rect 564712 400294 564780 400350
rect 564836 400294 571460 400350
rect 571516 400294 571584 400350
rect 571640 400294 578264 400350
rect 578320 400294 578388 400350
rect 578444 400294 585068 400350
rect 585124 400294 585192 400350
rect 585248 400294 596496 400350
rect 596552 400294 596620 400350
rect 596676 400294 596744 400350
rect 596800 400294 596868 400350
rect 596924 400294 597980 400350
rect -1916 400226 597980 400294
rect -1916 400170 -860 400226
rect -804 400170 -736 400226
rect -680 400170 -612 400226
rect -556 400170 -488 400226
rect -432 400170 3250 400226
rect 3306 400170 3374 400226
rect 3430 400170 3498 400226
rect 3554 400170 3622 400226
rect 3678 400170 21250 400226
rect 21306 400170 21374 400226
rect 21430 400170 21498 400226
rect 21554 400170 21622 400226
rect 21678 400170 39250 400226
rect 39306 400170 39374 400226
rect 39430 400170 39498 400226
rect 39554 400170 39622 400226
rect 39678 400170 57250 400226
rect 57306 400170 57374 400226
rect 57430 400170 57498 400226
rect 57554 400170 57622 400226
rect 57678 400170 93250 400226
rect 93306 400170 93374 400226
rect 93430 400170 93498 400226
rect 93554 400170 93622 400226
rect 93678 400170 111250 400226
rect 111306 400170 111374 400226
rect 111430 400170 111498 400226
rect 111554 400170 111622 400226
rect 111678 400170 129250 400226
rect 129306 400170 129374 400226
rect 129430 400170 129498 400226
rect 129554 400170 129622 400226
rect 129678 400170 147250 400226
rect 147306 400170 147374 400226
rect 147430 400170 147498 400226
rect 147554 400170 147622 400226
rect 147678 400170 183250 400226
rect 183306 400170 183374 400226
rect 183430 400170 183498 400226
rect 183554 400170 183622 400226
rect 183678 400170 201250 400226
rect 201306 400170 201374 400226
rect 201430 400170 201498 400226
rect 201554 400170 201622 400226
rect 201678 400170 219250 400226
rect 219306 400170 219374 400226
rect 219430 400170 219498 400226
rect 219554 400170 219622 400226
rect 219678 400170 237250 400226
rect 237306 400170 237374 400226
rect 237430 400170 237498 400226
rect 237554 400170 237622 400226
rect 237678 400170 273250 400226
rect 273306 400170 273374 400226
rect 273430 400170 273498 400226
rect 273554 400170 273622 400226
rect 273678 400170 291250 400226
rect 291306 400170 291374 400226
rect 291430 400170 291498 400226
rect 291554 400170 291622 400226
rect 291678 400170 309250 400226
rect 309306 400170 309374 400226
rect 309430 400170 309498 400226
rect 309554 400170 309622 400226
rect 309678 400170 327250 400226
rect 327306 400170 327374 400226
rect 327430 400170 327498 400226
rect 327554 400170 327622 400226
rect 327678 400170 363250 400226
rect 363306 400170 363374 400226
rect 363430 400170 363498 400226
rect 363554 400170 363622 400226
rect 363678 400170 381250 400226
rect 381306 400170 381374 400226
rect 381430 400170 381498 400226
rect 381554 400170 381622 400226
rect 381678 400170 399250 400226
rect 399306 400170 399374 400226
rect 399430 400170 399498 400226
rect 399554 400170 399622 400226
rect 399678 400170 417250 400226
rect 417306 400170 417374 400226
rect 417430 400170 417498 400226
rect 417554 400170 417622 400226
rect 417678 400170 453250 400226
rect 453306 400170 453374 400226
rect 453430 400170 453498 400226
rect 453554 400170 453622 400226
rect 453678 400170 471250 400226
rect 471306 400170 471374 400226
rect 471430 400170 471498 400226
rect 471554 400170 471622 400226
rect 471678 400170 489250 400226
rect 489306 400170 489374 400226
rect 489430 400170 489498 400226
rect 489554 400170 489622 400226
rect 489678 400170 507250 400226
rect 507306 400170 507374 400226
rect 507430 400170 507498 400226
rect 507554 400170 507622 400226
rect 507678 400170 543250 400226
rect 543306 400170 543374 400226
rect 543430 400170 543498 400226
rect 543554 400170 543622 400226
rect 543678 400170 564656 400226
rect 564712 400170 564780 400226
rect 564836 400170 571460 400226
rect 571516 400170 571584 400226
rect 571640 400170 578264 400226
rect 578320 400170 578388 400226
rect 578444 400170 585068 400226
rect 585124 400170 585192 400226
rect 585248 400170 596496 400226
rect 596552 400170 596620 400226
rect 596676 400170 596744 400226
rect 596800 400170 596868 400226
rect 596924 400170 597980 400226
rect -1916 400102 597980 400170
rect -1916 400046 -860 400102
rect -804 400046 -736 400102
rect -680 400046 -612 400102
rect -556 400046 -488 400102
rect -432 400046 3250 400102
rect 3306 400046 3374 400102
rect 3430 400046 3498 400102
rect 3554 400046 3622 400102
rect 3678 400046 21250 400102
rect 21306 400046 21374 400102
rect 21430 400046 21498 400102
rect 21554 400046 21622 400102
rect 21678 400046 39250 400102
rect 39306 400046 39374 400102
rect 39430 400046 39498 400102
rect 39554 400046 39622 400102
rect 39678 400046 57250 400102
rect 57306 400046 57374 400102
rect 57430 400046 57498 400102
rect 57554 400046 57622 400102
rect 57678 400046 93250 400102
rect 93306 400046 93374 400102
rect 93430 400046 93498 400102
rect 93554 400046 93622 400102
rect 93678 400046 111250 400102
rect 111306 400046 111374 400102
rect 111430 400046 111498 400102
rect 111554 400046 111622 400102
rect 111678 400046 129250 400102
rect 129306 400046 129374 400102
rect 129430 400046 129498 400102
rect 129554 400046 129622 400102
rect 129678 400046 147250 400102
rect 147306 400046 147374 400102
rect 147430 400046 147498 400102
rect 147554 400046 147622 400102
rect 147678 400046 183250 400102
rect 183306 400046 183374 400102
rect 183430 400046 183498 400102
rect 183554 400046 183622 400102
rect 183678 400046 201250 400102
rect 201306 400046 201374 400102
rect 201430 400046 201498 400102
rect 201554 400046 201622 400102
rect 201678 400046 219250 400102
rect 219306 400046 219374 400102
rect 219430 400046 219498 400102
rect 219554 400046 219622 400102
rect 219678 400046 237250 400102
rect 237306 400046 237374 400102
rect 237430 400046 237498 400102
rect 237554 400046 237622 400102
rect 237678 400046 273250 400102
rect 273306 400046 273374 400102
rect 273430 400046 273498 400102
rect 273554 400046 273622 400102
rect 273678 400046 291250 400102
rect 291306 400046 291374 400102
rect 291430 400046 291498 400102
rect 291554 400046 291622 400102
rect 291678 400046 309250 400102
rect 309306 400046 309374 400102
rect 309430 400046 309498 400102
rect 309554 400046 309622 400102
rect 309678 400046 327250 400102
rect 327306 400046 327374 400102
rect 327430 400046 327498 400102
rect 327554 400046 327622 400102
rect 327678 400046 363250 400102
rect 363306 400046 363374 400102
rect 363430 400046 363498 400102
rect 363554 400046 363622 400102
rect 363678 400046 381250 400102
rect 381306 400046 381374 400102
rect 381430 400046 381498 400102
rect 381554 400046 381622 400102
rect 381678 400046 399250 400102
rect 399306 400046 399374 400102
rect 399430 400046 399498 400102
rect 399554 400046 399622 400102
rect 399678 400046 417250 400102
rect 417306 400046 417374 400102
rect 417430 400046 417498 400102
rect 417554 400046 417622 400102
rect 417678 400046 453250 400102
rect 453306 400046 453374 400102
rect 453430 400046 453498 400102
rect 453554 400046 453622 400102
rect 453678 400046 471250 400102
rect 471306 400046 471374 400102
rect 471430 400046 471498 400102
rect 471554 400046 471622 400102
rect 471678 400046 489250 400102
rect 489306 400046 489374 400102
rect 489430 400046 489498 400102
rect 489554 400046 489622 400102
rect 489678 400046 507250 400102
rect 507306 400046 507374 400102
rect 507430 400046 507498 400102
rect 507554 400046 507622 400102
rect 507678 400046 543250 400102
rect 543306 400046 543374 400102
rect 543430 400046 543498 400102
rect 543554 400046 543622 400102
rect 543678 400046 564656 400102
rect 564712 400046 564780 400102
rect 564836 400046 571460 400102
rect 571516 400046 571584 400102
rect 571640 400046 578264 400102
rect 578320 400046 578388 400102
rect 578444 400046 585068 400102
rect 585124 400046 585192 400102
rect 585248 400046 596496 400102
rect 596552 400046 596620 400102
rect 596676 400046 596744 400102
rect 596800 400046 596868 400102
rect 596924 400046 597980 400102
rect -1916 399978 597980 400046
rect -1916 399922 -860 399978
rect -804 399922 -736 399978
rect -680 399922 -612 399978
rect -556 399922 -488 399978
rect -432 399922 3250 399978
rect 3306 399922 3374 399978
rect 3430 399922 3498 399978
rect 3554 399922 3622 399978
rect 3678 399922 21250 399978
rect 21306 399922 21374 399978
rect 21430 399922 21498 399978
rect 21554 399922 21622 399978
rect 21678 399922 39250 399978
rect 39306 399922 39374 399978
rect 39430 399922 39498 399978
rect 39554 399922 39622 399978
rect 39678 399922 57250 399978
rect 57306 399922 57374 399978
rect 57430 399922 57498 399978
rect 57554 399922 57622 399978
rect 57678 399922 93250 399978
rect 93306 399922 93374 399978
rect 93430 399922 93498 399978
rect 93554 399922 93622 399978
rect 93678 399922 111250 399978
rect 111306 399922 111374 399978
rect 111430 399922 111498 399978
rect 111554 399922 111622 399978
rect 111678 399922 129250 399978
rect 129306 399922 129374 399978
rect 129430 399922 129498 399978
rect 129554 399922 129622 399978
rect 129678 399922 147250 399978
rect 147306 399922 147374 399978
rect 147430 399922 147498 399978
rect 147554 399922 147622 399978
rect 147678 399922 183250 399978
rect 183306 399922 183374 399978
rect 183430 399922 183498 399978
rect 183554 399922 183622 399978
rect 183678 399922 201250 399978
rect 201306 399922 201374 399978
rect 201430 399922 201498 399978
rect 201554 399922 201622 399978
rect 201678 399922 219250 399978
rect 219306 399922 219374 399978
rect 219430 399922 219498 399978
rect 219554 399922 219622 399978
rect 219678 399922 237250 399978
rect 237306 399922 237374 399978
rect 237430 399922 237498 399978
rect 237554 399922 237622 399978
rect 237678 399922 273250 399978
rect 273306 399922 273374 399978
rect 273430 399922 273498 399978
rect 273554 399922 273622 399978
rect 273678 399922 291250 399978
rect 291306 399922 291374 399978
rect 291430 399922 291498 399978
rect 291554 399922 291622 399978
rect 291678 399922 309250 399978
rect 309306 399922 309374 399978
rect 309430 399922 309498 399978
rect 309554 399922 309622 399978
rect 309678 399922 327250 399978
rect 327306 399922 327374 399978
rect 327430 399922 327498 399978
rect 327554 399922 327622 399978
rect 327678 399922 363250 399978
rect 363306 399922 363374 399978
rect 363430 399922 363498 399978
rect 363554 399922 363622 399978
rect 363678 399922 381250 399978
rect 381306 399922 381374 399978
rect 381430 399922 381498 399978
rect 381554 399922 381622 399978
rect 381678 399922 399250 399978
rect 399306 399922 399374 399978
rect 399430 399922 399498 399978
rect 399554 399922 399622 399978
rect 399678 399922 417250 399978
rect 417306 399922 417374 399978
rect 417430 399922 417498 399978
rect 417554 399922 417622 399978
rect 417678 399922 453250 399978
rect 453306 399922 453374 399978
rect 453430 399922 453498 399978
rect 453554 399922 453622 399978
rect 453678 399922 471250 399978
rect 471306 399922 471374 399978
rect 471430 399922 471498 399978
rect 471554 399922 471622 399978
rect 471678 399922 489250 399978
rect 489306 399922 489374 399978
rect 489430 399922 489498 399978
rect 489554 399922 489622 399978
rect 489678 399922 507250 399978
rect 507306 399922 507374 399978
rect 507430 399922 507498 399978
rect 507554 399922 507622 399978
rect 507678 399922 543250 399978
rect 543306 399922 543374 399978
rect 543430 399922 543498 399978
rect 543554 399922 543622 399978
rect 543678 399922 564656 399978
rect 564712 399922 564780 399978
rect 564836 399922 571460 399978
rect 571516 399922 571584 399978
rect 571640 399922 578264 399978
rect 578320 399922 578388 399978
rect 578444 399922 585068 399978
rect 585124 399922 585192 399978
rect 585248 399922 596496 399978
rect 596552 399922 596620 399978
rect 596676 399922 596744 399978
rect 596800 399922 596868 399978
rect 596924 399922 597980 399978
rect -1916 399826 597980 399922
rect -1916 388350 597980 388446
rect -1916 388294 -1820 388350
rect -1764 388294 -1696 388350
rect -1640 388294 -1572 388350
rect -1516 388294 -1448 388350
rect -1392 388294 6970 388350
rect 7026 388294 7094 388350
rect 7150 388294 7218 388350
rect 7274 388294 7342 388350
rect 7398 388294 24970 388350
rect 25026 388294 25094 388350
rect 25150 388294 25218 388350
rect 25274 388294 25342 388350
rect 25398 388294 42970 388350
rect 43026 388294 43094 388350
rect 43150 388294 43218 388350
rect 43274 388294 43342 388350
rect 43398 388294 60970 388350
rect 61026 388294 61094 388350
rect 61150 388294 61218 388350
rect 61274 388294 61342 388350
rect 61398 388294 78970 388350
rect 79026 388294 79094 388350
rect 79150 388294 79218 388350
rect 79274 388294 79342 388350
rect 79398 388294 96970 388350
rect 97026 388294 97094 388350
rect 97150 388294 97218 388350
rect 97274 388294 97342 388350
rect 97398 388294 132970 388350
rect 133026 388294 133094 388350
rect 133150 388294 133218 388350
rect 133274 388294 133342 388350
rect 133398 388294 150970 388350
rect 151026 388294 151094 388350
rect 151150 388294 151218 388350
rect 151274 388294 151342 388350
rect 151398 388294 168970 388350
rect 169026 388294 169094 388350
rect 169150 388294 169218 388350
rect 169274 388294 169342 388350
rect 169398 388294 186970 388350
rect 187026 388294 187094 388350
rect 187150 388294 187218 388350
rect 187274 388294 187342 388350
rect 187398 388294 222970 388350
rect 223026 388294 223094 388350
rect 223150 388294 223218 388350
rect 223274 388294 223342 388350
rect 223398 388294 240970 388350
rect 241026 388294 241094 388350
rect 241150 388294 241218 388350
rect 241274 388294 241342 388350
rect 241398 388294 258970 388350
rect 259026 388294 259094 388350
rect 259150 388294 259218 388350
rect 259274 388294 259342 388350
rect 259398 388294 276970 388350
rect 277026 388294 277094 388350
rect 277150 388294 277218 388350
rect 277274 388294 277342 388350
rect 277398 388294 312970 388350
rect 313026 388294 313094 388350
rect 313150 388294 313218 388350
rect 313274 388294 313342 388350
rect 313398 388294 330970 388350
rect 331026 388294 331094 388350
rect 331150 388294 331218 388350
rect 331274 388294 331342 388350
rect 331398 388294 348970 388350
rect 349026 388294 349094 388350
rect 349150 388294 349218 388350
rect 349274 388294 349342 388350
rect 349398 388294 366970 388350
rect 367026 388294 367094 388350
rect 367150 388294 367218 388350
rect 367274 388294 367342 388350
rect 367398 388294 402970 388350
rect 403026 388294 403094 388350
rect 403150 388294 403218 388350
rect 403274 388294 403342 388350
rect 403398 388294 420970 388350
rect 421026 388294 421094 388350
rect 421150 388294 421218 388350
rect 421274 388294 421342 388350
rect 421398 388294 438970 388350
rect 439026 388294 439094 388350
rect 439150 388294 439218 388350
rect 439274 388294 439342 388350
rect 439398 388294 456970 388350
rect 457026 388294 457094 388350
rect 457150 388294 457218 388350
rect 457274 388294 457342 388350
rect 457398 388294 492970 388350
rect 493026 388294 493094 388350
rect 493150 388294 493218 388350
rect 493274 388294 493342 388350
rect 493398 388294 510970 388350
rect 511026 388294 511094 388350
rect 511150 388294 511218 388350
rect 511274 388294 511342 388350
rect 511398 388294 528970 388350
rect 529026 388294 529094 388350
rect 529150 388294 529218 388350
rect 529274 388294 529342 388350
rect 529398 388294 546970 388350
rect 547026 388294 547094 388350
rect 547150 388294 547218 388350
rect 547274 388294 547342 388350
rect 547398 388294 568058 388350
rect 568114 388294 568182 388350
rect 568238 388294 574862 388350
rect 574918 388294 574986 388350
rect 575042 388294 581666 388350
rect 581722 388294 581790 388350
rect 581846 388294 588470 388350
rect 588526 388294 588594 388350
rect 588650 388294 597456 388350
rect 597512 388294 597580 388350
rect 597636 388294 597704 388350
rect 597760 388294 597828 388350
rect 597884 388294 597980 388350
rect -1916 388226 597980 388294
rect -1916 388170 -1820 388226
rect -1764 388170 -1696 388226
rect -1640 388170 -1572 388226
rect -1516 388170 -1448 388226
rect -1392 388170 6970 388226
rect 7026 388170 7094 388226
rect 7150 388170 7218 388226
rect 7274 388170 7342 388226
rect 7398 388170 24970 388226
rect 25026 388170 25094 388226
rect 25150 388170 25218 388226
rect 25274 388170 25342 388226
rect 25398 388170 42970 388226
rect 43026 388170 43094 388226
rect 43150 388170 43218 388226
rect 43274 388170 43342 388226
rect 43398 388170 60970 388226
rect 61026 388170 61094 388226
rect 61150 388170 61218 388226
rect 61274 388170 61342 388226
rect 61398 388170 78970 388226
rect 79026 388170 79094 388226
rect 79150 388170 79218 388226
rect 79274 388170 79342 388226
rect 79398 388170 96970 388226
rect 97026 388170 97094 388226
rect 97150 388170 97218 388226
rect 97274 388170 97342 388226
rect 97398 388170 132970 388226
rect 133026 388170 133094 388226
rect 133150 388170 133218 388226
rect 133274 388170 133342 388226
rect 133398 388170 150970 388226
rect 151026 388170 151094 388226
rect 151150 388170 151218 388226
rect 151274 388170 151342 388226
rect 151398 388170 168970 388226
rect 169026 388170 169094 388226
rect 169150 388170 169218 388226
rect 169274 388170 169342 388226
rect 169398 388170 186970 388226
rect 187026 388170 187094 388226
rect 187150 388170 187218 388226
rect 187274 388170 187342 388226
rect 187398 388170 222970 388226
rect 223026 388170 223094 388226
rect 223150 388170 223218 388226
rect 223274 388170 223342 388226
rect 223398 388170 240970 388226
rect 241026 388170 241094 388226
rect 241150 388170 241218 388226
rect 241274 388170 241342 388226
rect 241398 388170 258970 388226
rect 259026 388170 259094 388226
rect 259150 388170 259218 388226
rect 259274 388170 259342 388226
rect 259398 388170 276970 388226
rect 277026 388170 277094 388226
rect 277150 388170 277218 388226
rect 277274 388170 277342 388226
rect 277398 388170 312970 388226
rect 313026 388170 313094 388226
rect 313150 388170 313218 388226
rect 313274 388170 313342 388226
rect 313398 388170 330970 388226
rect 331026 388170 331094 388226
rect 331150 388170 331218 388226
rect 331274 388170 331342 388226
rect 331398 388170 348970 388226
rect 349026 388170 349094 388226
rect 349150 388170 349218 388226
rect 349274 388170 349342 388226
rect 349398 388170 366970 388226
rect 367026 388170 367094 388226
rect 367150 388170 367218 388226
rect 367274 388170 367342 388226
rect 367398 388170 402970 388226
rect 403026 388170 403094 388226
rect 403150 388170 403218 388226
rect 403274 388170 403342 388226
rect 403398 388170 420970 388226
rect 421026 388170 421094 388226
rect 421150 388170 421218 388226
rect 421274 388170 421342 388226
rect 421398 388170 438970 388226
rect 439026 388170 439094 388226
rect 439150 388170 439218 388226
rect 439274 388170 439342 388226
rect 439398 388170 456970 388226
rect 457026 388170 457094 388226
rect 457150 388170 457218 388226
rect 457274 388170 457342 388226
rect 457398 388170 492970 388226
rect 493026 388170 493094 388226
rect 493150 388170 493218 388226
rect 493274 388170 493342 388226
rect 493398 388170 510970 388226
rect 511026 388170 511094 388226
rect 511150 388170 511218 388226
rect 511274 388170 511342 388226
rect 511398 388170 528970 388226
rect 529026 388170 529094 388226
rect 529150 388170 529218 388226
rect 529274 388170 529342 388226
rect 529398 388170 546970 388226
rect 547026 388170 547094 388226
rect 547150 388170 547218 388226
rect 547274 388170 547342 388226
rect 547398 388170 568058 388226
rect 568114 388170 568182 388226
rect 568238 388170 574862 388226
rect 574918 388170 574986 388226
rect 575042 388170 581666 388226
rect 581722 388170 581790 388226
rect 581846 388170 588470 388226
rect 588526 388170 588594 388226
rect 588650 388170 597456 388226
rect 597512 388170 597580 388226
rect 597636 388170 597704 388226
rect 597760 388170 597828 388226
rect 597884 388170 597980 388226
rect -1916 388102 597980 388170
rect -1916 388046 -1820 388102
rect -1764 388046 -1696 388102
rect -1640 388046 -1572 388102
rect -1516 388046 -1448 388102
rect -1392 388046 6970 388102
rect 7026 388046 7094 388102
rect 7150 388046 7218 388102
rect 7274 388046 7342 388102
rect 7398 388046 24970 388102
rect 25026 388046 25094 388102
rect 25150 388046 25218 388102
rect 25274 388046 25342 388102
rect 25398 388046 42970 388102
rect 43026 388046 43094 388102
rect 43150 388046 43218 388102
rect 43274 388046 43342 388102
rect 43398 388046 60970 388102
rect 61026 388046 61094 388102
rect 61150 388046 61218 388102
rect 61274 388046 61342 388102
rect 61398 388046 78970 388102
rect 79026 388046 79094 388102
rect 79150 388046 79218 388102
rect 79274 388046 79342 388102
rect 79398 388046 96970 388102
rect 97026 388046 97094 388102
rect 97150 388046 97218 388102
rect 97274 388046 97342 388102
rect 97398 388046 132970 388102
rect 133026 388046 133094 388102
rect 133150 388046 133218 388102
rect 133274 388046 133342 388102
rect 133398 388046 150970 388102
rect 151026 388046 151094 388102
rect 151150 388046 151218 388102
rect 151274 388046 151342 388102
rect 151398 388046 168970 388102
rect 169026 388046 169094 388102
rect 169150 388046 169218 388102
rect 169274 388046 169342 388102
rect 169398 388046 186970 388102
rect 187026 388046 187094 388102
rect 187150 388046 187218 388102
rect 187274 388046 187342 388102
rect 187398 388046 222970 388102
rect 223026 388046 223094 388102
rect 223150 388046 223218 388102
rect 223274 388046 223342 388102
rect 223398 388046 240970 388102
rect 241026 388046 241094 388102
rect 241150 388046 241218 388102
rect 241274 388046 241342 388102
rect 241398 388046 258970 388102
rect 259026 388046 259094 388102
rect 259150 388046 259218 388102
rect 259274 388046 259342 388102
rect 259398 388046 276970 388102
rect 277026 388046 277094 388102
rect 277150 388046 277218 388102
rect 277274 388046 277342 388102
rect 277398 388046 312970 388102
rect 313026 388046 313094 388102
rect 313150 388046 313218 388102
rect 313274 388046 313342 388102
rect 313398 388046 330970 388102
rect 331026 388046 331094 388102
rect 331150 388046 331218 388102
rect 331274 388046 331342 388102
rect 331398 388046 348970 388102
rect 349026 388046 349094 388102
rect 349150 388046 349218 388102
rect 349274 388046 349342 388102
rect 349398 388046 366970 388102
rect 367026 388046 367094 388102
rect 367150 388046 367218 388102
rect 367274 388046 367342 388102
rect 367398 388046 402970 388102
rect 403026 388046 403094 388102
rect 403150 388046 403218 388102
rect 403274 388046 403342 388102
rect 403398 388046 420970 388102
rect 421026 388046 421094 388102
rect 421150 388046 421218 388102
rect 421274 388046 421342 388102
rect 421398 388046 438970 388102
rect 439026 388046 439094 388102
rect 439150 388046 439218 388102
rect 439274 388046 439342 388102
rect 439398 388046 456970 388102
rect 457026 388046 457094 388102
rect 457150 388046 457218 388102
rect 457274 388046 457342 388102
rect 457398 388046 492970 388102
rect 493026 388046 493094 388102
rect 493150 388046 493218 388102
rect 493274 388046 493342 388102
rect 493398 388046 510970 388102
rect 511026 388046 511094 388102
rect 511150 388046 511218 388102
rect 511274 388046 511342 388102
rect 511398 388046 528970 388102
rect 529026 388046 529094 388102
rect 529150 388046 529218 388102
rect 529274 388046 529342 388102
rect 529398 388046 546970 388102
rect 547026 388046 547094 388102
rect 547150 388046 547218 388102
rect 547274 388046 547342 388102
rect 547398 388046 568058 388102
rect 568114 388046 568182 388102
rect 568238 388046 574862 388102
rect 574918 388046 574986 388102
rect 575042 388046 581666 388102
rect 581722 388046 581790 388102
rect 581846 388046 588470 388102
rect 588526 388046 588594 388102
rect 588650 388046 597456 388102
rect 597512 388046 597580 388102
rect 597636 388046 597704 388102
rect 597760 388046 597828 388102
rect 597884 388046 597980 388102
rect -1916 387978 597980 388046
rect -1916 387922 -1820 387978
rect -1764 387922 -1696 387978
rect -1640 387922 -1572 387978
rect -1516 387922 -1448 387978
rect -1392 387922 6970 387978
rect 7026 387922 7094 387978
rect 7150 387922 7218 387978
rect 7274 387922 7342 387978
rect 7398 387922 24970 387978
rect 25026 387922 25094 387978
rect 25150 387922 25218 387978
rect 25274 387922 25342 387978
rect 25398 387922 42970 387978
rect 43026 387922 43094 387978
rect 43150 387922 43218 387978
rect 43274 387922 43342 387978
rect 43398 387922 60970 387978
rect 61026 387922 61094 387978
rect 61150 387922 61218 387978
rect 61274 387922 61342 387978
rect 61398 387922 78970 387978
rect 79026 387922 79094 387978
rect 79150 387922 79218 387978
rect 79274 387922 79342 387978
rect 79398 387922 96970 387978
rect 97026 387922 97094 387978
rect 97150 387922 97218 387978
rect 97274 387922 97342 387978
rect 97398 387922 132970 387978
rect 133026 387922 133094 387978
rect 133150 387922 133218 387978
rect 133274 387922 133342 387978
rect 133398 387922 150970 387978
rect 151026 387922 151094 387978
rect 151150 387922 151218 387978
rect 151274 387922 151342 387978
rect 151398 387922 168970 387978
rect 169026 387922 169094 387978
rect 169150 387922 169218 387978
rect 169274 387922 169342 387978
rect 169398 387922 186970 387978
rect 187026 387922 187094 387978
rect 187150 387922 187218 387978
rect 187274 387922 187342 387978
rect 187398 387922 222970 387978
rect 223026 387922 223094 387978
rect 223150 387922 223218 387978
rect 223274 387922 223342 387978
rect 223398 387922 240970 387978
rect 241026 387922 241094 387978
rect 241150 387922 241218 387978
rect 241274 387922 241342 387978
rect 241398 387922 258970 387978
rect 259026 387922 259094 387978
rect 259150 387922 259218 387978
rect 259274 387922 259342 387978
rect 259398 387922 276970 387978
rect 277026 387922 277094 387978
rect 277150 387922 277218 387978
rect 277274 387922 277342 387978
rect 277398 387922 312970 387978
rect 313026 387922 313094 387978
rect 313150 387922 313218 387978
rect 313274 387922 313342 387978
rect 313398 387922 330970 387978
rect 331026 387922 331094 387978
rect 331150 387922 331218 387978
rect 331274 387922 331342 387978
rect 331398 387922 348970 387978
rect 349026 387922 349094 387978
rect 349150 387922 349218 387978
rect 349274 387922 349342 387978
rect 349398 387922 366970 387978
rect 367026 387922 367094 387978
rect 367150 387922 367218 387978
rect 367274 387922 367342 387978
rect 367398 387922 402970 387978
rect 403026 387922 403094 387978
rect 403150 387922 403218 387978
rect 403274 387922 403342 387978
rect 403398 387922 420970 387978
rect 421026 387922 421094 387978
rect 421150 387922 421218 387978
rect 421274 387922 421342 387978
rect 421398 387922 438970 387978
rect 439026 387922 439094 387978
rect 439150 387922 439218 387978
rect 439274 387922 439342 387978
rect 439398 387922 456970 387978
rect 457026 387922 457094 387978
rect 457150 387922 457218 387978
rect 457274 387922 457342 387978
rect 457398 387922 492970 387978
rect 493026 387922 493094 387978
rect 493150 387922 493218 387978
rect 493274 387922 493342 387978
rect 493398 387922 510970 387978
rect 511026 387922 511094 387978
rect 511150 387922 511218 387978
rect 511274 387922 511342 387978
rect 511398 387922 528970 387978
rect 529026 387922 529094 387978
rect 529150 387922 529218 387978
rect 529274 387922 529342 387978
rect 529398 387922 546970 387978
rect 547026 387922 547094 387978
rect 547150 387922 547218 387978
rect 547274 387922 547342 387978
rect 547398 387922 568058 387978
rect 568114 387922 568182 387978
rect 568238 387922 574862 387978
rect 574918 387922 574986 387978
rect 575042 387922 581666 387978
rect 581722 387922 581790 387978
rect 581846 387922 588470 387978
rect 588526 387922 588594 387978
rect 588650 387922 597456 387978
rect 597512 387922 597580 387978
rect 597636 387922 597704 387978
rect 597760 387922 597828 387978
rect 597884 387922 597980 387978
rect -1916 387826 597980 387922
rect -1916 382350 597980 382446
rect -1916 382294 -860 382350
rect -804 382294 -736 382350
rect -680 382294 -612 382350
rect -556 382294 -488 382350
rect -432 382294 3250 382350
rect 3306 382294 3374 382350
rect 3430 382294 3498 382350
rect 3554 382294 3622 382350
rect 3678 382294 21250 382350
rect 21306 382294 21374 382350
rect 21430 382294 21498 382350
rect 21554 382294 21622 382350
rect 21678 382294 39250 382350
rect 39306 382294 39374 382350
rect 39430 382294 39498 382350
rect 39554 382294 39622 382350
rect 39678 382294 57250 382350
rect 57306 382294 57374 382350
rect 57430 382294 57498 382350
rect 57554 382294 57622 382350
rect 57678 382294 93250 382350
rect 93306 382294 93374 382350
rect 93430 382294 93498 382350
rect 93554 382294 93622 382350
rect 93678 382294 111250 382350
rect 111306 382294 111374 382350
rect 111430 382294 111498 382350
rect 111554 382294 111622 382350
rect 111678 382294 129250 382350
rect 129306 382294 129374 382350
rect 129430 382294 129498 382350
rect 129554 382294 129622 382350
rect 129678 382294 147250 382350
rect 147306 382294 147374 382350
rect 147430 382294 147498 382350
rect 147554 382294 147622 382350
rect 147678 382294 183250 382350
rect 183306 382294 183374 382350
rect 183430 382294 183498 382350
rect 183554 382294 183622 382350
rect 183678 382294 201250 382350
rect 201306 382294 201374 382350
rect 201430 382294 201498 382350
rect 201554 382294 201622 382350
rect 201678 382294 219250 382350
rect 219306 382294 219374 382350
rect 219430 382294 219498 382350
rect 219554 382294 219622 382350
rect 219678 382294 237250 382350
rect 237306 382294 237374 382350
rect 237430 382294 237498 382350
rect 237554 382294 237622 382350
rect 237678 382294 273250 382350
rect 273306 382294 273374 382350
rect 273430 382294 273498 382350
rect 273554 382294 273622 382350
rect 273678 382294 291250 382350
rect 291306 382294 291374 382350
rect 291430 382294 291498 382350
rect 291554 382294 291622 382350
rect 291678 382294 309250 382350
rect 309306 382294 309374 382350
rect 309430 382294 309498 382350
rect 309554 382294 309622 382350
rect 309678 382294 327250 382350
rect 327306 382294 327374 382350
rect 327430 382294 327498 382350
rect 327554 382294 327622 382350
rect 327678 382294 363250 382350
rect 363306 382294 363374 382350
rect 363430 382294 363498 382350
rect 363554 382294 363622 382350
rect 363678 382294 381250 382350
rect 381306 382294 381374 382350
rect 381430 382294 381498 382350
rect 381554 382294 381622 382350
rect 381678 382294 399250 382350
rect 399306 382294 399374 382350
rect 399430 382294 399498 382350
rect 399554 382294 399622 382350
rect 399678 382294 417250 382350
rect 417306 382294 417374 382350
rect 417430 382294 417498 382350
rect 417554 382294 417622 382350
rect 417678 382294 453250 382350
rect 453306 382294 453374 382350
rect 453430 382294 453498 382350
rect 453554 382294 453622 382350
rect 453678 382294 471250 382350
rect 471306 382294 471374 382350
rect 471430 382294 471498 382350
rect 471554 382294 471622 382350
rect 471678 382294 489250 382350
rect 489306 382294 489374 382350
rect 489430 382294 489498 382350
rect 489554 382294 489622 382350
rect 489678 382294 507250 382350
rect 507306 382294 507374 382350
rect 507430 382294 507498 382350
rect 507554 382294 507622 382350
rect 507678 382294 543250 382350
rect 543306 382294 543374 382350
rect 543430 382294 543498 382350
rect 543554 382294 543622 382350
rect 543678 382294 564656 382350
rect 564712 382294 564780 382350
rect 564836 382294 571460 382350
rect 571516 382294 571584 382350
rect 571640 382294 578264 382350
rect 578320 382294 578388 382350
rect 578444 382294 585068 382350
rect 585124 382294 585192 382350
rect 585248 382294 596496 382350
rect 596552 382294 596620 382350
rect 596676 382294 596744 382350
rect 596800 382294 596868 382350
rect 596924 382294 597980 382350
rect -1916 382226 597980 382294
rect -1916 382170 -860 382226
rect -804 382170 -736 382226
rect -680 382170 -612 382226
rect -556 382170 -488 382226
rect -432 382170 3250 382226
rect 3306 382170 3374 382226
rect 3430 382170 3498 382226
rect 3554 382170 3622 382226
rect 3678 382170 21250 382226
rect 21306 382170 21374 382226
rect 21430 382170 21498 382226
rect 21554 382170 21622 382226
rect 21678 382170 39250 382226
rect 39306 382170 39374 382226
rect 39430 382170 39498 382226
rect 39554 382170 39622 382226
rect 39678 382170 57250 382226
rect 57306 382170 57374 382226
rect 57430 382170 57498 382226
rect 57554 382170 57622 382226
rect 57678 382170 93250 382226
rect 93306 382170 93374 382226
rect 93430 382170 93498 382226
rect 93554 382170 93622 382226
rect 93678 382170 111250 382226
rect 111306 382170 111374 382226
rect 111430 382170 111498 382226
rect 111554 382170 111622 382226
rect 111678 382170 129250 382226
rect 129306 382170 129374 382226
rect 129430 382170 129498 382226
rect 129554 382170 129622 382226
rect 129678 382170 147250 382226
rect 147306 382170 147374 382226
rect 147430 382170 147498 382226
rect 147554 382170 147622 382226
rect 147678 382170 183250 382226
rect 183306 382170 183374 382226
rect 183430 382170 183498 382226
rect 183554 382170 183622 382226
rect 183678 382170 201250 382226
rect 201306 382170 201374 382226
rect 201430 382170 201498 382226
rect 201554 382170 201622 382226
rect 201678 382170 219250 382226
rect 219306 382170 219374 382226
rect 219430 382170 219498 382226
rect 219554 382170 219622 382226
rect 219678 382170 237250 382226
rect 237306 382170 237374 382226
rect 237430 382170 237498 382226
rect 237554 382170 237622 382226
rect 237678 382170 273250 382226
rect 273306 382170 273374 382226
rect 273430 382170 273498 382226
rect 273554 382170 273622 382226
rect 273678 382170 291250 382226
rect 291306 382170 291374 382226
rect 291430 382170 291498 382226
rect 291554 382170 291622 382226
rect 291678 382170 309250 382226
rect 309306 382170 309374 382226
rect 309430 382170 309498 382226
rect 309554 382170 309622 382226
rect 309678 382170 327250 382226
rect 327306 382170 327374 382226
rect 327430 382170 327498 382226
rect 327554 382170 327622 382226
rect 327678 382170 363250 382226
rect 363306 382170 363374 382226
rect 363430 382170 363498 382226
rect 363554 382170 363622 382226
rect 363678 382170 381250 382226
rect 381306 382170 381374 382226
rect 381430 382170 381498 382226
rect 381554 382170 381622 382226
rect 381678 382170 399250 382226
rect 399306 382170 399374 382226
rect 399430 382170 399498 382226
rect 399554 382170 399622 382226
rect 399678 382170 417250 382226
rect 417306 382170 417374 382226
rect 417430 382170 417498 382226
rect 417554 382170 417622 382226
rect 417678 382170 453250 382226
rect 453306 382170 453374 382226
rect 453430 382170 453498 382226
rect 453554 382170 453622 382226
rect 453678 382170 471250 382226
rect 471306 382170 471374 382226
rect 471430 382170 471498 382226
rect 471554 382170 471622 382226
rect 471678 382170 489250 382226
rect 489306 382170 489374 382226
rect 489430 382170 489498 382226
rect 489554 382170 489622 382226
rect 489678 382170 507250 382226
rect 507306 382170 507374 382226
rect 507430 382170 507498 382226
rect 507554 382170 507622 382226
rect 507678 382170 543250 382226
rect 543306 382170 543374 382226
rect 543430 382170 543498 382226
rect 543554 382170 543622 382226
rect 543678 382170 564656 382226
rect 564712 382170 564780 382226
rect 564836 382170 571460 382226
rect 571516 382170 571584 382226
rect 571640 382170 578264 382226
rect 578320 382170 578388 382226
rect 578444 382170 585068 382226
rect 585124 382170 585192 382226
rect 585248 382170 596496 382226
rect 596552 382170 596620 382226
rect 596676 382170 596744 382226
rect 596800 382170 596868 382226
rect 596924 382170 597980 382226
rect -1916 382102 597980 382170
rect -1916 382046 -860 382102
rect -804 382046 -736 382102
rect -680 382046 -612 382102
rect -556 382046 -488 382102
rect -432 382046 3250 382102
rect 3306 382046 3374 382102
rect 3430 382046 3498 382102
rect 3554 382046 3622 382102
rect 3678 382046 21250 382102
rect 21306 382046 21374 382102
rect 21430 382046 21498 382102
rect 21554 382046 21622 382102
rect 21678 382046 39250 382102
rect 39306 382046 39374 382102
rect 39430 382046 39498 382102
rect 39554 382046 39622 382102
rect 39678 382046 57250 382102
rect 57306 382046 57374 382102
rect 57430 382046 57498 382102
rect 57554 382046 57622 382102
rect 57678 382046 93250 382102
rect 93306 382046 93374 382102
rect 93430 382046 93498 382102
rect 93554 382046 93622 382102
rect 93678 382046 111250 382102
rect 111306 382046 111374 382102
rect 111430 382046 111498 382102
rect 111554 382046 111622 382102
rect 111678 382046 129250 382102
rect 129306 382046 129374 382102
rect 129430 382046 129498 382102
rect 129554 382046 129622 382102
rect 129678 382046 147250 382102
rect 147306 382046 147374 382102
rect 147430 382046 147498 382102
rect 147554 382046 147622 382102
rect 147678 382046 183250 382102
rect 183306 382046 183374 382102
rect 183430 382046 183498 382102
rect 183554 382046 183622 382102
rect 183678 382046 201250 382102
rect 201306 382046 201374 382102
rect 201430 382046 201498 382102
rect 201554 382046 201622 382102
rect 201678 382046 219250 382102
rect 219306 382046 219374 382102
rect 219430 382046 219498 382102
rect 219554 382046 219622 382102
rect 219678 382046 237250 382102
rect 237306 382046 237374 382102
rect 237430 382046 237498 382102
rect 237554 382046 237622 382102
rect 237678 382046 273250 382102
rect 273306 382046 273374 382102
rect 273430 382046 273498 382102
rect 273554 382046 273622 382102
rect 273678 382046 291250 382102
rect 291306 382046 291374 382102
rect 291430 382046 291498 382102
rect 291554 382046 291622 382102
rect 291678 382046 309250 382102
rect 309306 382046 309374 382102
rect 309430 382046 309498 382102
rect 309554 382046 309622 382102
rect 309678 382046 327250 382102
rect 327306 382046 327374 382102
rect 327430 382046 327498 382102
rect 327554 382046 327622 382102
rect 327678 382046 363250 382102
rect 363306 382046 363374 382102
rect 363430 382046 363498 382102
rect 363554 382046 363622 382102
rect 363678 382046 381250 382102
rect 381306 382046 381374 382102
rect 381430 382046 381498 382102
rect 381554 382046 381622 382102
rect 381678 382046 399250 382102
rect 399306 382046 399374 382102
rect 399430 382046 399498 382102
rect 399554 382046 399622 382102
rect 399678 382046 417250 382102
rect 417306 382046 417374 382102
rect 417430 382046 417498 382102
rect 417554 382046 417622 382102
rect 417678 382046 453250 382102
rect 453306 382046 453374 382102
rect 453430 382046 453498 382102
rect 453554 382046 453622 382102
rect 453678 382046 471250 382102
rect 471306 382046 471374 382102
rect 471430 382046 471498 382102
rect 471554 382046 471622 382102
rect 471678 382046 489250 382102
rect 489306 382046 489374 382102
rect 489430 382046 489498 382102
rect 489554 382046 489622 382102
rect 489678 382046 507250 382102
rect 507306 382046 507374 382102
rect 507430 382046 507498 382102
rect 507554 382046 507622 382102
rect 507678 382046 543250 382102
rect 543306 382046 543374 382102
rect 543430 382046 543498 382102
rect 543554 382046 543622 382102
rect 543678 382046 564656 382102
rect 564712 382046 564780 382102
rect 564836 382046 571460 382102
rect 571516 382046 571584 382102
rect 571640 382046 578264 382102
rect 578320 382046 578388 382102
rect 578444 382046 585068 382102
rect 585124 382046 585192 382102
rect 585248 382046 596496 382102
rect 596552 382046 596620 382102
rect 596676 382046 596744 382102
rect 596800 382046 596868 382102
rect 596924 382046 597980 382102
rect -1916 381978 597980 382046
rect -1916 381922 -860 381978
rect -804 381922 -736 381978
rect -680 381922 -612 381978
rect -556 381922 -488 381978
rect -432 381922 3250 381978
rect 3306 381922 3374 381978
rect 3430 381922 3498 381978
rect 3554 381922 3622 381978
rect 3678 381922 21250 381978
rect 21306 381922 21374 381978
rect 21430 381922 21498 381978
rect 21554 381922 21622 381978
rect 21678 381922 39250 381978
rect 39306 381922 39374 381978
rect 39430 381922 39498 381978
rect 39554 381922 39622 381978
rect 39678 381922 57250 381978
rect 57306 381922 57374 381978
rect 57430 381922 57498 381978
rect 57554 381922 57622 381978
rect 57678 381922 93250 381978
rect 93306 381922 93374 381978
rect 93430 381922 93498 381978
rect 93554 381922 93622 381978
rect 93678 381922 111250 381978
rect 111306 381922 111374 381978
rect 111430 381922 111498 381978
rect 111554 381922 111622 381978
rect 111678 381922 129250 381978
rect 129306 381922 129374 381978
rect 129430 381922 129498 381978
rect 129554 381922 129622 381978
rect 129678 381922 147250 381978
rect 147306 381922 147374 381978
rect 147430 381922 147498 381978
rect 147554 381922 147622 381978
rect 147678 381922 183250 381978
rect 183306 381922 183374 381978
rect 183430 381922 183498 381978
rect 183554 381922 183622 381978
rect 183678 381922 201250 381978
rect 201306 381922 201374 381978
rect 201430 381922 201498 381978
rect 201554 381922 201622 381978
rect 201678 381922 219250 381978
rect 219306 381922 219374 381978
rect 219430 381922 219498 381978
rect 219554 381922 219622 381978
rect 219678 381922 237250 381978
rect 237306 381922 237374 381978
rect 237430 381922 237498 381978
rect 237554 381922 237622 381978
rect 237678 381922 273250 381978
rect 273306 381922 273374 381978
rect 273430 381922 273498 381978
rect 273554 381922 273622 381978
rect 273678 381922 291250 381978
rect 291306 381922 291374 381978
rect 291430 381922 291498 381978
rect 291554 381922 291622 381978
rect 291678 381922 309250 381978
rect 309306 381922 309374 381978
rect 309430 381922 309498 381978
rect 309554 381922 309622 381978
rect 309678 381922 327250 381978
rect 327306 381922 327374 381978
rect 327430 381922 327498 381978
rect 327554 381922 327622 381978
rect 327678 381922 363250 381978
rect 363306 381922 363374 381978
rect 363430 381922 363498 381978
rect 363554 381922 363622 381978
rect 363678 381922 381250 381978
rect 381306 381922 381374 381978
rect 381430 381922 381498 381978
rect 381554 381922 381622 381978
rect 381678 381922 399250 381978
rect 399306 381922 399374 381978
rect 399430 381922 399498 381978
rect 399554 381922 399622 381978
rect 399678 381922 417250 381978
rect 417306 381922 417374 381978
rect 417430 381922 417498 381978
rect 417554 381922 417622 381978
rect 417678 381922 453250 381978
rect 453306 381922 453374 381978
rect 453430 381922 453498 381978
rect 453554 381922 453622 381978
rect 453678 381922 471250 381978
rect 471306 381922 471374 381978
rect 471430 381922 471498 381978
rect 471554 381922 471622 381978
rect 471678 381922 489250 381978
rect 489306 381922 489374 381978
rect 489430 381922 489498 381978
rect 489554 381922 489622 381978
rect 489678 381922 507250 381978
rect 507306 381922 507374 381978
rect 507430 381922 507498 381978
rect 507554 381922 507622 381978
rect 507678 381922 543250 381978
rect 543306 381922 543374 381978
rect 543430 381922 543498 381978
rect 543554 381922 543622 381978
rect 543678 381922 564656 381978
rect 564712 381922 564780 381978
rect 564836 381922 571460 381978
rect 571516 381922 571584 381978
rect 571640 381922 578264 381978
rect 578320 381922 578388 381978
rect 578444 381922 585068 381978
rect 585124 381922 585192 381978
rect 585248 381922 596496 381978
rect 596552 381922 596620 381978
rect 596676 381922 596744 381978
rect 596800 381922 596868 381978
rect 596924 381922 597980 381978
rect -1916 381826 597980 381922
rect -1916 370350 597980 370446
rect -1916 370294 -1820 370350
rect -1764 370294 -1696 370350
rect -1640 370294 -1572 370350
rect -1516 370294 -1448 370350
rect -1392 370294 6970 370350
rect 7026 370294 7094 370350
rect 7150 370294 7218 370350
rect 7274 370294 7342 370350
rect 7398 370294 24970 370350
rect 25026 370294 25094 370350
rect 25150 370294 25218 370350
rect 25274 370294 25342 370350
rect 25398 370294 42970 370350
rect 43026 370294 43094 370350
rect 43150 370294 43218 370350
rect 43274 370294 43342 370350
rect 43398 370294 60970 370350
rect 61026 370294 61094 370350
rect 61150 370294 61218 370350
rect 61274 370294 61342 370350
rect 61398 370294 78970 370350
rect 79026 370294 79094 370350
rect 79150 370294 79218 370350
rect 79274 370294 79342 370350
rect 79398 370294 96970 370350
rect 97026 370294 97094 370350
rect 97150 370294 97218 370350
rect 97274 370294 97342 370350
rect 97398 370294 132970 370350
rect 133026 370294 133094 370350
rect 133150 370294 133218 370350
rect 133274 370294 133342 370350
rect 133398 370294 150970 370350
rect 151026 370294 151094 370350
rect 151150 370294 151218 370350
rect 151274 370294 151342 370350
rect 151398 370294 168970 370350
rect 169026 370294 169094 370350
rect 169150 370294 169218 370350
rect 169274 370294 169342 370350
rect 169398 370294 186970 370350
rect 187026 370294 187094 370350
rect 187150 370294 187218 370350
rect 187274 370294 187342 370350
rect 187398 370294 222970 370350
rect 223026 370294 223094 370350
rect 223150 370294 223218 370350
rect 223274 370294 223342 370350
rect 223398 370294 240970 370350
rect 241026 370294 241094 370350
rect 241150 370294 241218 370350
rect 241274 370294 241342 370350
rect 241398 370294 258970 370350
rect 259026 370294 259094 370350
rect 259150 370294 259218 370350
rect 259274 370294 259342 370350
rect 259398 370294 276970 370350
rect 277026 370294 277094 370350
rect 277150 370294 277218 370350
rect 277274 370294 277342 370350
rect 277398 370294 312970 370350
rect 313026 370294 313094 370350
rect 313150 370294 313218 370350
rect 313274 370294 313342 370350
rect 313398 370294 330970 370350
rect 331026 370294 331094 370350
rect 331150 370294 331218 370350
rect 331274 370294 331342 370350
rect 331398 370294 348970 370350
rect 349026 370294 349094 370350
rect 349150 370294 349218 370350
rect 349274 370294 349342 370350
rect 349398 370294 366970 370350
rect 367026 370294 367094 370350
rect 367150 370294 367218 370350
rect 367274 370294 367342 370350
rect 367398 370294 402970 370350
rect 403026 370294 403094 370350
rect 403150 370294 403218 370350
rect 403274 370294 403342 370350
rect 403398 370294 420970 370350
rect 421026 370294 421094 370350
rect 421150 370294 421218 370350
rect 421274 370294 421342 370350
rect 421398 370294 438970 370350
rect 439026 370294 439094 370350
rect 439150 370294 439218 370350
rect 439274 370294 439342 370350
rect 439398 370294 456970 370350
rect 457026 370294 457094 370350
rect 457150 370294 457218 370350
rect 457274 370294 457342 370350
rect 457398 370294 492970 370350
rect 493026 370294 493094 370350
rect 493150 370294 493218 370350
rect 493274 370294 493342 370350
rect 493398 370294 510970 370350
rect 511026 370294 511094 370350
rect 511150 370294 511218 370350
rect 511274 370294 511342 370350
rect 511398 370294 528970 370350
rect 529026 370294 529094 370350
rect 529150 370294 529218 370350
rect 529274 370294 529342 370350
rect 529398 370294 546970 370350
rect 547026 370294 547094 370350
rect 547150 370294 547218 370350
rect 547274 370294 547342 370350
rect 547398 370294 564970 370350
rect 565026 370294 565094 370350
rect 565150 370294 565218 370350
rect 565274 370294 565342 370350
rect 565398 370294 582970 370350
rect 583026 370294 583094 370350
rect 583150 370294 583218 370350
rect 583274 370294 583342 370350
rect 583398 370294 597456 370350
rect 597512 370294 597580 370350
rect 597636 370294 597704 370350
rect 597760 370294 597828 370350
rect 597884 370294 597980 370350
rect -1916 370226 597980 370294
rect -1916 370170 -1820 370226
rect -1764 370170 -1696 370226
rect -1640 370170 -1572 370226
rect -1516 370170 -1448 370226
rect -1392 370170 6970 370226
rect 7026 370170 7094 370226
rect 7150 370170 7218 370226
rect 7274 370170 7342 370226
rect 7398 370170 24970 370226
rect 25026 370170 25094 370226
rect 25150 370170 25218 370226
rect 25274 370170 25342 370226
rect 25398 370170 42970 370226
rect 43026 370170 43094 370226
rect 43150 370170 43218 370226
rect 43274 370170 43342 370226
rect 43398 370170 60970 370226
rect 61026 370170 61094 370226
rect 61150 370170 61218 370226
rect 61274 370170 61342 370226
rect 61398 370170 78970 370226
rect 79026 370170 79094 370226
rect 79150 370170 79218 370226
rect 79274 370170 79342 370226
rect 79398 370170 96970 370226
rect 97026 370170 97094 370226
rect 97150 370170 97218 370226
rect 97274 370170 97342 370226
rect 97398 370170 132970 370226
rect 133026 370170 133094 370226
rect 133150 370170 133218 370226
rect 133274 370170 133342 370226
rect 133398 370170 150970 370226
rect 151026 370170 151094 370226
rect 151150 370170 151218 370226
rect 151274 370170 151342 370226
rect 151398 370170 168970 370226
rect 169026 370170 169094 370226
rect 169150 370170 169218 370226
rect 169274 370170 169342 370226
rect 169398 370170 186970 370226
rect 187026 370170 187094 370226
rect 187150 370170 187218 370226
rect 187274 370170 187342 370226
rect 187398 370170 222970 370226
rect 223026 370170 223094 370226
rect 223150 370170 223218 370226
rect 223274 370170 223342 370226
rect 223398 370170 240970 370226
rect 241026 370170 241094 370226
rect 241150 370170 241218 370226
rect 241274 370170 241342 370226
rect 241398 370170 258970 370226
rect 259026 370170 259094 370226
rect 259150 370170 259218 370226
rect 259274 370170 259342 370226
rect 259398 370170 276970 370226
rect 277026 370170 277094 370226
rect 277150 370170 277218 370226
rect 277274 370170 277342 370226
rect 277398 370170 312970 370226
rect 313026 370170 313094 370226
rect 313150 370170 313218 370226
rect 313274 370170 313342 370226
rect 313398 370170 330970 370226
rect 331026 370170 331094 370226
rect 331150 370170 331218 370226
rect 331274 370170 331342 370226
rect 331398 370170 348970 370226
rect 349026 370170 349094 370226
rect 349150 370170 349218 370226
rect 349274 370170 349342 370226
rect 349398 370170 366970 370226
rect 367026 370170 367094 370226
rect 367150 370170 367218 370226
rect 367274 370170 367342 370226
rect 367398 370170 402970 370226
rect 403026 370170 403094 370226
rect 403150 370170 403218 370226
rect 403274 370170 403342 370226
rect 403398 370170 420970 370226
rect 421026 370170 421094 370226
rect 421150 370170 421218 370226
rect 421274 370170 421342 370226
rect 421398 370170 438970 370226
rect 439026 370170 439094 370226
rect 439150 370170 439218 370226
rect 439274 370170 439342 370226
rect 439398 370170 456970 370226
rect 457026 370170 457094 370226
rect 457150 370170 457218 370226
rect 457274 370170 457342 370226
rect 457398 370170 492970 370226
rect 493026 370170 493094 370226
rect 493150 370170 493218 370226
rect 493274 370170 493342 370226
rect 493398 370170 510970 370226
rect 511026 370170 511094 370226
rect 511150 370170 511218 370226
rect 511274 370170 511342 370226
rect 511398 370170 528970 370226
rect 529026 370170 529094 370226
rect 529150 370170 529218 370226
rect 529274 370170 529342 370226
rect 529398 370170 546970 370226
rect 547026 370170 547094 370226
rect 547150 370170 547218 370226
rect 547274 370170 547342 370226
rect 547398 370170 564970 370226
rect 565026 370170 565094 370226
rect 565150 370170 565218 370226
rect 565274 370170 565342 370226
rect 565398 370170 582970 370226
rect 583026 370170 583094 370226
rect 583150 370170 583218 370226
rect 583274 370170 583342 370226
rect 583398 370170 597456 370226
rect 597512 370170 597580 370226
rect 597636 370170 597704 370226
rect 597760 370170 597828 370226
rect 597884 370170 597980 370226
rect -1916 370102 597980 370170
rect -1916 370046 -1820 370102
rect -1764 370046 -1696 370102
rect -1640 370046 -1572 370102
rect -1516 370046 -1448 370102
rect -1392 370046 6970 370102
rect 7026 370046 7094 370102
rect 7150 370046 7218 370102
rect 7274 370046 7342 370102
rect 7398 370046 24970 370102
rect 25026 370046 25094 370102
rect 25150 370046 25218 370102
rect 25274 370046 25342 370102
rect 25398 370046 42970 370102
rect 43026 370046 43094 370102
rect 43150 370046 43218 370102
rect 43274 370046 43342 370102
rect 43398 370046 60970 370102
rect 61026 370046 61094 370102
rect 61150 370046 61218 370102
rect 61274 370046 61342 370102
rect 61398 370046 78970 370102
rect 79026 370046 79094 370102
rect 79150 370046 79218 370102
rect 79274 370046 79342 370102
rect 79398 370046 96970 370102
rect 97026 370046 97094 370102
rect 97150 370046 97218 370102
rect 97274 370046 97342 370102
rect 97398 370046 132970 370102
rect 133026 370046 133094 370102
rect 133150 370046 133218 370102
rect 133274 370046 133342 370102
rect 133398 370046 150970 370102
rect 151026 370046 151094 370102
rect 151150 370046 151218 370102
rect 151274 370046 151342 370102
rect 151398 370046 168970 370102
rect 169026 370046 169094 370102
rect 169150 370046 169218 370102
rect 169274 370046 169342 370102
rect 169398 370046 186970 370102
rect 187026 370046 187094 370102
rect 187150 370046 187218 370102
rect 187274 370046 187342 370102
rect 187398 370046 222970 370102
rect 223026 370046 223094 370102
rect 223150 370046 223218 370102
rect 223274 370046 223342 370102
rect 223398 370046 240970 370102
rect 241026 370046 241094 370102
rect 241150 370046 241218 370102
rect 241274 370046 241342 370102
rect 241398 370046 258970 370102
rect 259026 370046 259094 370102
rect 259150 370046 259218 370102
rect 259274 370046 259342 370102
rect 259398 370046 276970 370102
rect 277026 370046 277094 370102
rect 277150 370046 277218 370102
rect 277274 370046 277342 370102
rect 277398 370046 312970 370102
rect 313026 370046 313094 370102
rect 313150 370046 313218 370102
rect 313274 370046 313342 370102
rect 313398 370046 330970 370102
rect 331026 370046 331094 370102
rect 331150 370046 331218 370102
rect 331274 370046 331342 370102
rect 331398 370046 348970 370102
rect 349026 370046 349094 370102
rect 349150 370046 349218 370102
rect 349274 370046 349342 370102
rect 349398 370046 366970 370102
rect 367026 370046 367094 370102
rect 367150 370046 367218 370102
rect 367274 370046 367342 370102
rect 367398 370046 402970 370102
rect 403026 370046 403094 370102
rect 403150 370046 403218 370102
rect 403274 370046 403342 370102
rect 403398 370046 420970 370102
rect 421026 370046 421094 370102
rect 421150 370046 421218 370102
rect 421274 370046 421342 370102
rect 421398 370046 438970 370102
rect 439026 370046 439094 370102
rect 439150 370046 439218 370102
rect 439274 370046 439342 370102
rect 439398 370046 456970 370102
rect 457026 370046 457094 370102
rect 457150 370046 457218 370102
rect 457274 370046 457342 370102
rect 457398 370046 492970 370102
rect 493026 370046 493094 370102
rect 493150 370046 493218 370102
rect 493274 370046 493342 370102
rect 493398 370046 510970 370102
rect 511026 370046 511094 370102
rect 511150 370046 511218 370102
rect 511274 370046 511342 370102
rect 511398 370046 528970 370102
rect 529026 370046 529094 370102
rect 529150 370046 529218 370102
rect 529274 370046 529342 370102
rect 529398 370046 546970 370102
rect 547026 370046 547094 370102
rect 547150 370046 547218 370102
rect 547274 370046 547342 370102
rect 547398 370046 564970 370102
rect 565026 370046 565094 370102
rect 565150 370046 565218 370102
rect 565274 370046 565342 370102
rect 565398 370046 582970 370102
rect 583026 370046 583094 370102
rect 583150 370046 583218 370102
rect 583274 370046 583342 370102
rect 583398 370046 597456 370102
rect 597512 370046 597580 370102
rect 597636 370046 597704 370102
rect 597760 370046 597828 370102
rect 597884 370046 597980 370102
rect -1916 369978 597980 370046
rect -1916 369922 -1820 369978
rect -1764 369922 -1696 369978
rect -1640 369922 -1572 369978
rect -1516 369922 -1448 369978
rect -1392 369922 6970 369978
rect 7026 369922 7094 369978
rect 7150 369922 7218 369978
rect 7274 369922 7342 369978
rect 7398 369922 24970 369978
rect 25026 369922 25094 369978
rect 25150 369922 25218 369978
rect 25274 369922 25342 369978
rect 25398 369922 42970 369978
rect 43026 369922 43094 369978
rect 43150 369922 43218 369978
rect 43274 369922 43342 369978
rect 43398 369922 60970 369978
rect 61026 369922 61094 369978
rect 61150 369922 61218 369978
rect 61274 369922 61342 369978
rect 61398 369922 78970 369978
rect 79026 369922 79094 369978
rect 79150 369922 79218 369978
rect 79274 369922 79342 369978
rect 79398 369922 96970 369978
rect 97026 369922 97094 369978
rect 97150 369922 97218 369978
rect 97274 369922 97342 369978
rect 97398 369922 132970 369978
rect 133026 369922 133094 369978
rect 133150 369922 133218 369978
rect 133274 369922 133342 369978
rect 133398 369922 150970 369978
rect 151026 369922 151094 369978
rect 151150 369922 151218 369978
rect 151274 369922 151342 369978
rect 151398 369922 168970 369978
rect 169026 369922 169094 369978
rect 169150 369922 169218 369978
rect 169274 369922 169342 369978
rect 169398 369922 186970 369978
rect 187026 369922 187094 369978
rect 187150 369922 187218 369978
rect 187274 369922 187342 369978
rect 187398 369922 222970 369978
rect 223026 369922 223094 369978
rect 223150 369922 223218 369978
rect 223274 369922 223342 369978
rect 223398 369922 240970 369978
rect 241026 369922 241094 369978
rect 241150 369922 241218 369978
rect 241274 369922 241342 369978
rect 241398 369922 258970 369978
rect 259026 369922 259094 369978
rect 259150 369922 259218 369978
rect 259274 369922 259342 369978
rect 259398 369922 276970 369978
rect 277026 369922 277094 369978
rect 277150 369922 277218 369978
rect 277274 369922 277342 369978
rect 277398 369922 312970 369978
rect 313026 369922 313094 369978
rect 313150 369922 313218 369978
rect 313274 369922 313342 369978
rect 313398 369922 330970 369978
rect 331026 369922 331094 369978
rect 331150 369922 331218 369978
rect 331274 369922 331342 369978
rect 331398 369922 348970 369978
rect 349026 369922 349094 369978
rect 349150 369922 349218 369978
rect 349274 369922 349342 369978
rect 349398 369922 366970 369978
rect 367026 369922 367094 369978
rect 367150 369922 367218 369978
rect 367274 369922 367342 369978
rect 367398 369922 402970 369978
rect 403026 369922 403094 369978
rect 403150 369922 403218 369978
rect 403274 369922 403342 369978
rect 403398 369922 420970 369978
rect 421026 369922 421094 369978
rect 421150 369922 421218 369978
rect 421274 369922 421342 369978
rect 421398 369922 438970 369978
rect 439026 369922 439094 369978
rect 439150 369922 439218 369978
rect 439274 369922 439342 369978
rect 439398 369922 456970 369978
rect 457026 369922 457094 369978
rect 457150 369922 457218 369978
rect 457274 369922 457342 369978
rect 457398 369922 492970 369978
rect 493026 369922 493094 369978
rect 493150 369922 493218 369978
rect 493274 369922 493342 369978
rect 493398 369922 510970 369978
rect 511026 369922 511094 369978
rect 511150 369922 511218 369978
rect 511274 369922 511342 369978
rect 511398 369922 528970 369978
rect 529026 369922 529094 369978
rect 529150 369922 529218 369978
rect 529274 369922 529342 369978
rect 529398 369922 546970 369978
rect 547026 369922 547094 369978
rect 547150 369922 547218 369978
rect 547274 369922 547342 369978
rect 547398 369922 564970 369978
rect 565026 369922 565094 369978
rect 565150 369922 565218 369978
rect 565274 369922 565342 369978
rect 565398 369922 582970 369978
rect 583026 369922 583094 369978
rect 583150 369922 583218 369978
rect 583274 369922 583342 369978
rect 583398 369922 597456 369978
rect 597512 369922 597580 369978
rect 597636 369922 597704 369978
rect 597760 369922 597828 369978
rect 597884 369922 597980 369978
rect -1916 369826 597980 369922
rect -1916 364350 597980 364446
rect -1916 364294 -860 364350
rect -804 364294 -736 364350
rect -680 364294 -612 364350
rect -556 364294 -488 364350
rect -432 364294 3250 364350
rect 3306 364294 3374 364350
rect 3430 364294 3498 364350
rect 3554 364294 3622 364350
rect 3678 364294 21250 364350
rect 21306 364294 21374 364350
rect 21430 364294 21498 364350
rect 21554 364294 21622 364350
rect 21678 364294 39250 364350
rect 39306 364294 39374 364350
rect 39430 364294 39498 364350
rect 39554 364294 39622 364350
rect 39678 364294 57250 364350
rect 57306 364294 57374 364350
rect 57430 364294 57498 364350
rect 57554 364294 57622 364350
rect 57678 364294 93250 364350
rect 93306 364294 93374 364350
rect 93430 364294 93498 364350
rect 93554 364294 93622 364350
rect 93678 364294 111250 364350
rect 111306 364294 111374 364350
rect 111430 364294 111498 364350
rect 111554 364294 111622 364350
rect 111678 364294 129250 364350
rect 129306 364294 129374 364350
rect 129430 364294 129498 364350
rect 129554 364294 129622 364350
rect 129678 364294 147250 364350
rect 147306 364294 147374 364350
rect 147430 364294 147498 364350
rect 147554 364294 147622 364350
rect 147678 364294 183250 364350
rect 183306 364294 183374 364350
rect 183430 364294 183498 364350
rect 183554 364294 183622 364350
rect 183678 364294 201250 364350
rect 201306 364294 201374 364350
rect 201430 364294 201498 364350
rect 201554 364294 201622 364350
rect 201678 364294 219250 364350
rect 219306 364294 219374 364350
rect 219430 364294 219498 364350
rect 219554 364294 219622 364350
rect 219678 364294 237250 364350
rect 237306 364294 237374 364350
rect 237430 364294 237498 364350
rect 237554 364294 237622 364350
rect 237678 364294 273250 364350
rect 273306 364294 273374 364350
rect 273430 364294 273498 364350
rect 273554 364294 273622 364350
rect 273678 364294 291250 364350
rect 291306 364294 291374 364350
rect 291430 364294 291498 364350
rect 291554 364294 291622 364350
rect 291678 364294 309250 364350
rect 309306 364294 309374 364350
rect 309430 364294 309498 364350
rect 309554 364294 309622 364350
rect 309678 364294 327250 364350
rect 327306 364294 327374 364350
rect 327430 364294 327498 364350
rect 327554 364294 327622 364350
rect 327678 364294 363250 364350
rect 363306 364294 363374 364350
rect 363430 364294 363498 364350
rect 363554 364294 363622 364350
rect 363678 364294 381250 364350
rect 381306 364294 381374 364350
rect 381430 364294 381498 364350
rect 381554 364294 381622 364350
rect 381678 364294 399250 364350
rect 399306 364294 399374 364350
rect 399430 364294 399498 364350
rect 399554 364294 399622 364350
rect 399678 364294 417250 364350
rect 417306 364294 417374 364350
rect 417430 364294 417498 364350
rect 417554 364294 417622 364350
rect 417678 364294 453250 364350
rect 453306 364294 453374 364350
rect 453430 364294 453498 364350
rect 453554 364294 453622 364350
rect 453678 364294 471250 364350
rect 471306 364294 471374 364350
rect 471430 364294 471498 364350
rect 471554 364294 471622 364350
rect 471678 364294 489250 364350
rect 489306 364294 489374 364350
rect 489430 364294 489498 364350
rect 489554 364294 489622 364350
rect 489678 364294 507250 364350
rect 507306 364294 507374 364350
rect 507430 364294 507498 364350
rect 507554 364294 507622 364350
rect 507678 364294 543250 364350
rect 543306 364294 543374 364350
rect 543430 364294 543498 364350
rect 543554 364294 543622 364350
rect 543678 364294 561250 364350
rect 561306 364294 561374 364350
rect 561430 364294 561498 364350
rect 561554 364294 561622 364350
rect 561678 364294 579250 364350
rect 579306 364294 579374 364350
rect 579430 364294 579498 364350
rect 579554 364294 579622 364350
rect 579678 364294 596496 364350
rect 596552 364294 596620 364350
rect 596676 364294 596744 364350
rect 596800 364294 596868 364350
rect 596924 364294 597980 364350
rect -1916 364226 597980 364294
rect -1916 364170 -860 364226
rect -804 364170 -736 364226
rect -680 364170 -612 364226
rect -556 364170 -488 364226
rect -432 364170 3250 364226
rect 3306 364170 3374 364226
rect 3430 364170 3498 364226
rect 3554 364170 3622 364226
rect 3678 364170 21250 364226
rect 21306 364170 21374 364226
rect 21430 364170 21498 364226
rect 21554 364170 21622 364226
rect 21678 364170 39250 364226
rect 39306 364170 39374 364226
rect 39430 364170 39498 364226
rect 39554 364170 39622 364226
rect 39678 364170 57250 364226
rect 57306 364170 57374 364226
rect 57430 364170 57498 364226
rect 57554 364170 57622 364226
rect 57678 364170 93250 364226
rect 93306 364170 93374 364226
rect 93430 364170 93498 364226
rect 93554 364170 93622 364226
rect 93678 364170 111250 364226
rect 111306 364170 111374 364226
rect 111430 364170 111498 364226
rect 111554 364170 111622 364226
rect 111678 364170 129250 364226
rect 129306 364170 129374 364226
rect 129430 364170 129498 364226
rect 129554 364170 129622 364226
rect 129678 364170 147250 364226
rect 147306 364170 147374 364226
rect 147430 364170 147498 364226
rect 147554 364170 147622 364226
rect 147678 364170 183250 364226
rect 183306 364170 183374 364226
rect 183430 364170 183498 364226
rect 183554 364170 183622 364226
rect 183678 364170 201250 364226
rect 201306 364170 201374 364226
rect 201430 364170 201498 364226
rect 201554 364170 201622 364226
rect 201678 364170 219250 364226
rect 219306 364170 219374 364226
rect 219430 364170 219498 364226
rect 219554 364170 219622 364226
rect 219678 364170 237250 364226
rect 237306 364170 237374 364226
rect 237430 364170 237498 364226
rect 237554 364170 237622 364226
rect 237678 364170 273250 364226
rect 273306 364170 273374 364226
rect 273430 364170 273498 364226
rect 273554 364170 273622 364226
rect 273678 364170 291250 364226
rect 291306 364170 291374 364226
rect 291430 364170 291498 364226
rect 291554 364170 291622 364226
rect 291678 364170 309250 364226
rect 309306 364170 309374 364226
rect 309430 364170 309498 364226
rect 309554 364170 309622 364226
rect 309678 364170 327250 364226
rect 327306 364170 327374 364226
rect 327430 364170 327498 364226
rect 327554 364170 327622 364226
rect 327678 364170 363250 364226
rect 363306 364170 363374 364226
rect 363430 364170 363498 364226
rect 363554 364170 363622 364226
rect 363678 364170 381250 364226
rect 381306 364170 381374 364226
rect 381430 364170 381498 364226
rect 381554 364170 381622 364226
rect 381678 364170 399250 364226
rect 399306 364170 399374 364226
rect 399430 364170 399498 364226
rect 399554 364170 399622 364226
rect 399678 364170 417250 364226
rect 417306 364170 417374 364226
rect 417430 364170 417498 364226
rect 417554 364170 417622 364226
rect 417678 364170 453250 364226
rect 453306 364170 453374 364226
rect 453430 364170 453498 364226
rect 453554 364170 453622 364226
rect 453678 364170 471250 364226
rect 471306 364170 471374 364226
rect 471430 364170 471498 364226
rect 471554 364170 471622 364226
rect 471678 364170 489250 364226
rect 489306 364170 489374 364226
rect 489430 364170 489498 364226
rect 489554 364170 489622 364226
rect 489678 364170 507250 364226
rect 507306 364170 507374 364226
rect 507430 364170 507498 364226
rect 507554 364170 507622 364226
rect 507678 364170 543250 364226
rect 543306 364170 543374 364226
rect 543430 364170 543498 364226
rect 543554 364170 543622 364226
rect 543678 364170 561250 364226
rect 561306 364170 561374 364226
rect 561430 364170 561498 364226
rect 561554 364170 561622 364226
rect 561678 364170 579250 364226
rect 579306 364170 579374 364226
rect 579430 364170 579498 364226
rect 579554 364170 579622 364226
rect 579678 364170 596496 364226
rect 596552 364170 596620 364226
rect 596676 364170 596744 364226
rect 596800 364170 596868 364226
rect 596924 364170 597980 364226
rect -1916 364102 597980 364170
rect -1916 364046 -860 364102
rect -804 364046 -736 364102
rect -680 364046 -612 364102
rect -556 364046 -488 364102
rect -432 364046 3250 364102
rect 3306 364046 3374 364102
rect 3430 364046 3498 364102
rect 3554 364046 3622 364102
rect 3678 364046 21250 364102
rect 21306 364046 21374 364102
rect 21430 364046 21498 364102
rect 21554 364046 21622 364102
rect 21678 364046 39250 364102
rect 39306 364046 39374 364102
rect 39430 364046 39498 364102
rect 39554 364046 39622 364102
rect 39678 364046 57250 364102
rect 57306 364046 57374 364102
rect 57430 364046 57498 364102
rect 57554 364046 57622 364102
rect 57678 364046 93250 364102
rect 93306 364046 93374 364102
rect 93430 364046 93498 364102
rect 93554 364046 93622 364102
rect 93678 364046 111250 364102
rect 111306 364046 111374 364102
rect 111430 364046 111498 364102
rect 111554 364046 111622 364102
rect 111678 364046 129250 364102
rect 129306 364046 129374 364102
rect 129430 364046 129498 364102
rect 129554 364046 129622 364102
rect 129678 364046 147250 364102
rect 147306 364046 147374 364102
rect 147430 364046 147498 364102
rect 147554 364046 147622 364102
rect 147678 364046 183250 364102
rect 183306 364046 183374 364102
rect 183430 364046 183498 364102
rect 183554 364046 183622 364102
rect 183678 364046 201250 364102
rect 201306 364046 201374 364102
rect 201430 364046 201498 364102
rect 201554 364046 201622 364102
rect 201678 364046 219250 364102
rect 219306 364046 219374 364102
rect 219430 364046 219498 364102
rect 219554 364046 219622 364102
rect 219678 364046 237250 364102
rect 237306 364046 237374 364102
rect 237430 364046 237498 364102
rect 237554 364046 237622 364102
rect 237678 364046 273250 364102
rect 273306 364046 273374 364102
rect 273430 364046 273498 364102
rect 273554 364046 273622 364102
rect 273678 364046 291250 364102
rect 291306 364046 291374 364102
rect 291430 364046 291498 364102
rect 291554 364046 291622 364102
rect 291678 364046 309250 364102
rect 309306 364046 309374 364102
rect 309430 364046 309498 364102
rect 309554 364046 309622 364102
rect 309678 364046 327250 364102
rect 327306 364046 327374 364102
rect 327430 364046 327498 364102
rect 327554 364046 327622 364102
rect 327678 364046 363250 364102
rect 363306 364046 363374 364102
rect 363430 364046 363498 364102
rect 363554 364046 363622 364102
rect 363678 364046 381250 364102
rect 381306 364046 381374 364102
rect 381430 364046 381498 364102
rect 381554 364046 381622 364102
rect 381678 364046 399250 364102
rect 399306 364046 399374 364102
rect 399430 364046 399498 364102
rect 399554 364046 399622 364102
rect 399678 364046 417250 364102
rect 417306 364046 417374 364102
rect 417430 364046 417498 364102
rect 417554 364046 417622 364102
rect 417678 364046 453250 364102
rect 453306 364046 453374 364102
rect 453430 364046 453498 364102
rect 453554 364046 453622 364102
rect 453678 364046 471250 364102
rect 471306 364046 471374 364102
rect 471430 364046 471498 364102
rect 471554 364046 471622 364102
rect 471678 364046 489250 364102
rect 489306 364046 489374 364102
rect 489430 364046 489498 364102
rect 489554 364046 489622 364102
rect 489678 364046 507250 364102
rect 507306 364046 507374 364102
rect 507430 364046 507498 364102
rect 507554 364046 507622 364102
rect 507678 364046 543250 364102
rect 543306 364046 543374 364102
rect 543430 364046 543498 364102
rect 543554 364046 543622 364102
rect 543678 364046 561250 364102
rect 561306 364046 561374 364102
rect 561430 364046 561498 364102
rect 561554 364046 561622 364102
rect 561678 364046 579250 364102
rect 579306 364046 579374 364102
rect 579430 364046 579498 364102
rect 579554 364046 579622 364102
rect 579678 364046 596496 364102
rect 596552 364046 596620 364102
rect 596676 364046 596744 364102
rect 596800 364046 596868 364102
rect 596924 364046 597980 364102
rect -1916 363978 597980 364046
rect -1916 363922 -860 363978
rect -804 363922 -736 363978
rect -680 363922 -612 363978
rect -556 363922 -488 363978
rect -432 363922 3250 363978
rect 3306 363922 3374 363978
rect 3430 363922 3498 363978
rect 3554 363922 3622 363978
rect 3678 363922 21250 363978
rect 21306 363922 21374 363978
rect 21430 363922 21498 363978
rect 21554 363922 21622 363978
rect 21678 363922 39250 363978
rect 39306 363922 39374 363978
rect 39430 363922 39498 363978
rect 39554 363922 39622 363978
rect 39678 363922 57250 363978
rect 57306 363922 57374 363978
rect 57430 363922 57498 363978
rect 57554 363922 57622 363978
rect 57678 363922 93250 363978
rect 93306 363922 93374 363978
rect 93430 363922 93498 363978
rect 93554 363922 93622 363978
rect 93678 363922 111250 363978
rect 111306 363922 111374 363978
rect 111430 363922 111498 363978
rect 111554 363922 111622 363978
rect 111678 363922 129250 363978
rect 129306 363922 129374 363978
rect 129430 363922 129498 363978
rect 129554 363922 129622 363978
rect 129678 363922 147250 363978
rect 147306 363922 147374 363978
rect 147430 363922 147498 363978
rect 147554 363922 147622 363978
rect 147678 363922 183250 363978
rect 183306 363922 183374 363978
rect 183430 363922 183498 363978
rect 183554 363922 183622 363978
rect 183678 363922 201250 363978
rect 201306 363922 201374 363978
rect 201430 363922 201498 363978
rect 201554 363922 201622 363978
rect 201678 363922 219250 363978
rect 219306 363922 219374 363978
rect 219430 363922 219498 363978
rect 219554 363922 219622 363978
rect 219678 363922 237250 363978
rect 237306 363922 237374 363978
rect 237430 363922 237498 363978
rect 237554 363922 237622 363978
rect 237678 363922 273250 363978
rect 273306 363922 273374 363978
rect 273430 363922 273498 363978
rect 273554 363922 273622 363978
rect 273678 363922 291250 363978
rect 291306 363922 291374 363978
rect 291430 363922 291498 363978
rect 291554 363922 291622 363978
rect 291678 363922 309250 363978
rect 309306 363922 309374 363978
rect 309430 363922 309498 363978
rect 309554 363922 309622 363978
rect 309678 363922 327250 363978
rect 327306 363922 327374 363978
rect 327430 363922 327498 363978
rect 327554 363922 327622 363978
rect 327678 363922 363250 363978
rect 363306 363922 363374 363978
rect 363430 363922 363498 363978
rect 363554 363922 363622 363978
rect 363678 363922 381250 363978
rect 381306 363922 381374 363978
rect 381430 363922 381498 363978
rect 381554 363922 381622 363978
rect 381678 363922 399250 363978
rect 399306 363922 399374 363978
rect 399430 363922 399498 363978
rect 399554 363922 399622 363978
rect 399678 363922 417250 363978
rect 417306 363922 417374 363978
rect 417430 363922 417498 363978
rect 417554 363922 417622 363978
rect 417678 363922 453250 363978
rect 453306 363922 453374 363978
rect 453430 363922 453498 363978
rect 453554 363922 453622 363978
rect 453678 363922 471250 363978
rect 471306 363922 471374 363978
rect 471430 363922 471498 363978
rect 471554 363922 471622 363978
rect 471678 363922 489250 363978
rect 489306 363922 489374 363978
rect 489430 363922 489498 363978
rect 489554 363922 489622 363978
rect 489678 363922 507250 363978
rect 507306 363922 507374 363978
rect 507430 363922 507498 363978
rect 507554 363922 507622 363978
rect 507678 363922 543250 363978
rect 543306 363922 543374 363978
rect 543430 363922 543498 363978
rect 543554 363922 543622 363978
rect 543678 363922 561250 363978
rect 561306 363922 561374 363978
rect 561430 363922 561498 363978
rect 561554 363922 561622 363978
rect 561678 363922 579250 363978
rect 579306 363922 579374 363978
rect 579430 363922 579498 363978
rect 579554 363922 579622 363978
rect 579678 363922 596496 363978
rect 596552 363922 596620 363978
rect 596676 363922 596744 363978
rect 596800 363922 596868 363978
rect 596924 363922 597980 363978
rect -1916 363826 597980 363922
rect -1916 352350 597980 352446
rect -1916 352294 -1820 352350
rect -1764 352294 -1696 352350
rect -1640 352294 -1572 352350
rect -1516 352294 -1448 352350
rect -1392 352294 6970 352350
rect 7026 352294 7094 352350
rect 7150 352294 7218 352350
rect 7274 352294 7342 352350
rect 7398 352294 24970 352350
rect 25026 352294 25094 352350
rect 25150 352294 25218 352350
rect 25274 352294 25342 352350
rect 25398 352294 42970 352350
rect 43026 352294 43094 352350
rect 43150 352294 43218 352350
rect 43274 352294 43342 352350
rect 43398 352294 60970 352350
rect 61026 352294 61094 352350
rect 61150 352294 61218 352350
rect 61274 352294 61342 352350
rect 61398 352294 78970 352350
rect 79026 352294 79094 352350
rect 79150 352294 79218 352350
rect 79274 352294 79342 352350
rect 79398 352294 96970 352350
rect 97026 352294 97094 352350
rect 97150 352294 97218 352350
rect 97274 352294 97342 352350
rect 97398 352294 132970 352350
rect 133026 352294 133094 352350
rect 133150 352294 133218 352350
rect 133274 352294 133342 352350
rect 133398 352294 150970 352350
rect 151026 352294 151094 352350
rect 151150 352294 151218 352350
rect 151274 352294 151342 352350
rect 151398 352294 168970 352350
rect 169026 352294 169094 352350
rect 169150 352294 169218 352350
rect 169274 352294 169342 352350
rect 169398 352294 186970 352350
rect 187026 352294 187094 352350
rect 187150 352294 187218 352350
rect 187274 352294 187342 352350
rect 187398 352294 222970 352350
rect 223026 352294 223094 352350
rect 223150 352294 223218 352350
rect 223274 352294 223342 352350
rect 223398 352294 240970 352350
rect 241026 352294 241094 352350
rect 241150 352294 241218 352350
rect 241274 352294 241342 352350
rect 241398 352294 258970 352350
rect 259026 352294 259094 352350
rect 259150 352294 259218 352350
rect 259274 352294 259342 352350
rect 259398 352294 276970 352350
rect 277026 352294 277094 352350
rect 277150 352294 277218 352350
rect 277274 352294 277342 352350
rect 277398 352294 312970 352350
rect 313026 352294 313094 352350
rect 313150 352294 313218 352350
rect 313274 352294 313342 352350
rect 313398 352294 330970 352350
rect 331026 352294 331094 352350
rect 331150 352294 331218 352350
rect 331274 352294 331342 352350
rect 331398 352294 348970 352350
rect 349026 352294 349094 352350
rect 349150 352294 349218 352350
rect 349274 352294 349342 352350
rect 349398 352294 366970 352350
rect 367026 352294 367094 352350
rect 367150 352294 367218 352350
rect 367274 352294 367342 352350
rect 367398 352294 402970 352350
rect 403026 352294 403094 352350
rect 403150 352294 403218 352350
rect 403274 352294 403342 352350
rect 403398 352294 420970 352350
rect 421026 352294 421094 352350
rect 421150 352294 421218 352350
rect 421274 352294 421342 352350
rect 421398 352294 438970 352350
rect 439026 352294 439094 352350
rect 439150 352294 439218 352350
rect 439274 352294 439342 352350
rect 439398 352294 456970 352350
rect 457026 352294 457094 352350
rect 457150 352294 457218 352350
rect 457274 352294 457342 352350
rect 457398 352294 492970 352350
rect 493026 352294 493094 352350
rect 493150 352294 493218 352350
rect 493274 352294 493342 352350
rect 493398 352294 510970 352350
rect 511026 352294 511094 352350
rect 511150 352294 511218 352350
rect 511274 352294 511342 352350
rect 511398 352294 528970 352350
rect 529026 352294 529094 352350
rect 529150 352294 529218 352350
rect 529274 352294 529342 352350
rect 529398 352294 546970 352350
rect 547026 352294 547094 352350
rect 547150 352294 547218 352350
rect 547274 352294 547342 352350
rect 547398 352294 564970 352350
rect 565026 352294 565094 352350
rect 565150 352294 565218 352350
rect 565274 352294 565342 352350
rect 565398 352294 582970 352350
rect 583026 352294 583094 352350
rect 583150 352294 583218 352350
rect 583274 352294 583342 352350
rect 583398 352294 597456 352350
rect 597512 352294 597580 352350
rect 597636 352294 597704 352350
rect 597760 352294 597828 352350
rect 597884 352294 597980 352350
rect -1916 352226 597980 352294
rect -1916 352170 -1820 352226
rect -1764 352170 -1696 352226
rect -1640 352170 -1572 352226
rect -1516 352170 -1448 352226
rect -1392 352170 6970 352226
rect 7026 352170 7094 352226
rect 7150 352170 7218 352226
rect 7274 352170 7342 352226
rect 7398 352170 24970 352226
rect 25026 352170 25094 352226
rect 25150 352170 25218 352226
rect 25274 352170 25342 352226
rect 25398 352170 42970 352226
rect 43026 352170 43094 352226
rect 43150 352170 43218 352226
rect 43274 352170 43342 352226
rect 43398 352170 60970 352226
rect 61026 352170 61094 352226
rect 61150 352170 61218 352226
rect 61274 352170 61342 352226
rect 61398 352170 78970 352226
rect 79026 352170 79094 352226
rect 79150 352170 79218 352226
rect 79274 352170 79342 352226
rect 79398 352170 96970 352226
rect 97026 352170 97094 352226
rect 97150 352170 97218 352226
rect 97274 352170 97342 352226
rect 97398 352170 132970 352226
rect 133026 352170 133094 352226
rect 133150 352170 133218 352226
rect 133274 352170 133342 352226
rect 133398 352170 150970 352226
rect 151026 352170 151094 352226
rect 151150 352170 151218 352226
rect 151274 352170 151342 352226
rect 151398 352170 168970 352226
rect 169026 352170 169094 352226
rect 169150 352170 169218 352226
rect 169274 352170 169342 352226
rect 169398 352170 186970 352226
rect 187026 352170 187094 352226
rect 187150 352170 187218 352226
rect 187274 352170 187342 352226
rect 187398 352170 222970 352226
rect 223026 352170 223094 352226
rect 223150 352170 223218 352226
rect 223274 352170 223342 352226
rect 223398 352170 240970 352226
rect 241026 352170 241094 352226
rect 241150 352170 241218 352226
rect 241274 352170 241342 352226
rect 241398 352170 258970 352226
rect 259026 352170 259094 352226
rect 259150 352170 259218 352226
rect 259274 352170 259342 352226
rect 259398 352170 276970 352226
rect 277026 352170 277094 352226
rect 277150 352170 277218 352226
rect 277274 352170 277342 352226
rect 277398 352170 312970 352226
rect 313026 352170 313094 352226
rect 313150 352170 313218 352226
rect 313274 352170 313342 352226
rect 313398 352170 330970 352226
rect 331026 352170 331094 352226
rect 331150 352170 331218 352226
rect 331274 352170 331342 352226
rect 331398 352170 348970 352226
rect 349026 352170 349094 352226
rect 349150 352170 349218 352226
rect 349274 352170 349342 352226
rect 349398 352170 366970 352226
rect 367026 352170 367094 352226
rect 367150 352170 367218 352226
rect 367274 352170 367342 352226
rect 367398 352170 402970 352226
rect 403026 352170 403094 352226
rect 403150 352170 403218 352226
rect 403274 352170 403342 352226
rect 403398 352170 420970 352226
rect 421026 352170 421094 352226
rect 421150 352170 421218 352226
rect 421274 352170 421342 352226
rect 421398 352170 438970 352226
rect 439026 352170 439094 352226
rect 439150 352170 439218 352226
rect 439274 352170 439342 352226
rect 439398 352170 456970 352226
rect 457026 352170 457094 352226
rect 457150 352170 457218 352226
rect 457274 352170 457342 352226
rect 457398 352170 492970 352226
rect 493026 352170 493094 352226
rect 493150 352170 493218 352226
rect 493274 352170 493342 352226
rect 493398 352170 510970 352226
rect 511026 352170 511094 352226
rect 511150 352170 511218 352226
rect 511274 352170 511342 352226
rect 511398 352170 528970 352226
rect 529026 352170 529094 352226
rect 529150 352170 529218 352226
rect 529274 352170 529342 352226
rect 529398 352170 546970 352226
rect 547026 352170 547094 352226
rect 547150 352170 547218 352226
rect 547274 352170 547342 352226
rect 547398 352170 564970 352226
rect 565026 352170 565094 352226
rect 565150 352170 565218 352226
rect 565274 352170 565342 352226
rect 565398 352170 582970 352226
rect 583026 352170 583094 352226
rect 583150 352170 583218 352226
rect 583274 352170 583342 352226
rect 583398 352170 597456 352226
rect 597512 352170 597580 352226
rect 597636 352170 597704 352226
rect 597760 352170 597828 352226
rect 597884 352170 597980 352226
rect -1916 352102 597980 352170
rect -1916 352046 -1820 352102
rect -1764 352046 -1696 352102
rect -1640 352046 -1572 352102
rect -1516 352046 -1448 352102
rect -1392 352046 6970 352102
rect 7026 352046 7094 352102
rect 7150 352046 7218 352102
rect 7274 352046 7342 352102
rect 7398 352046 24970 352102
rect 25026 352046 25094 352102
rect 25150 352046 25218 352102
rect 25274 352046 25342 352102
rect 25398 352046 42970 352102
rect 43026 352046 43094 352102
rect 43150 352046 43218 352102
rect 43274 352046 43342 352102
rect 43398 352046 60970 352102
rect 61026 352046 61094 352102
rect 61150 352046 61218 352102
rect 61274 352046 61342 352102
rect 61398 352046 78970 352102
rect 79026 352046 79094 352102
rect 79150 352046 79218 352102
rect 79274 352046 79342 352102
rect 79398 352046 96970 352102
rect 97026 352046 97094 352102
rect 97150 352046 97218 352102
rect 97274 352046 97342 352102
rect 97398 352046 132970 352102
rect 133026 352046 133094 352102
rect 133150 352046 133218 352102
rect 133274 352046 133342 352102
rect 133398 352046 150970 352102
rect 151026 352046 151094 352102
rect 151150 352046 151218 352102
rect 151274 352046 151342 352102
rect 151398 352046 168970 352102
rect 169026 352046 169094 352102
rect 169150 352046 169218 352102
rect 169274 352046 169342 352102
rect 169398 352046 186970 352102
rect 187026 352046 187094 352102
rect 187150 352046 187218 352102
rect 187274 352046 187342 352102
rect 187398 352046 222970 352102
rect 223026 352046 223094 352102
rect 223150 352046 223218 352102
rect 223274 352046 223342 352102
rect 223398 352046 240970 352102
rect 241026 352046 241094 352102
rect 241150 352046 241218 352102
rect 241274 352046 241342 352102
rect 241398 352046 258970 352102
rect 259026 352046 259094 352102
rect 259150 352046 259218 352102
rect 259274 352046 259342 352102
rect 259398 352046 276970 352102
rect 277026 352046 277094 352102
rect 277150 352046 277218 352102
rect 277274 352046 277342 352102
rect 277398 352046 312970 352102
rect 313026 352046 313094 352102
rect 313150 352046 313218 352102
rect 313274 352046 313342 352102
rect 313398 352046 330970 352102
rect 331026 352046 331094 352102
rect 331150 352046 331218 352102
rect 331274 352046 331342 352102
rect 331398 352046 348970 352102
rect 349026 352046 349094 352102
rect 349150 352046 349218 352102
rect 349274 352046 349342 352102
rect 349398 352046 366970 352102
rect 367026 352046 367094 352102
rect 367150 352046 367218 352102
rect 367274 352046 367342 352102
rect 367398 352046 402970 352102
rect 403026 352046 403094 352102
rect 403150 352046 403218 352102
rect 403274 352046 403342 352102
rect 403398 352046 420970 352102
rect 421026 352046 421094 352102
rect 421150 352046 421218 352102
rect 421274 352046 421342 352102
rect 421398 352046 438970 352102
rect 439026 352046 439094 352102
rect 439150 352046 439218 352102
rect 439274 352046 439342 352102
rect 439398 352046 456970 352102
rect 457026 352046 457094 352102
rect 457150 352046 457218 352102
rect 457274 352046 457342 352102
rect 457398 352046 492970 352102
rect 493026 352046 493094 352102
rect 493150 352046 493218 352102
rect 493274 352046 493342 352102
rect 493398 352046 510970 352102
rect 511026 352046 511094 352102
rect 511150 352046 511218 352102
rect 511274 352046 511342 352102
rect 511398 352046 528970 352102
rect 529026 352046 529094 352102
rect 529150 352046 529218 352102
rect 529274 352046 529342 352102
rect 529398 352046 546970 352102
rect 547026 352046 547094 352102
rect 547150 352046 547218 352102
rect 547274 352046 547342 352102
rect 547398 352046 564970 352102
rect 565026 352046 565094 352102
rect 565150 352046 565218 352102
rect 565274 352046 565342 352102
rect 565398 352046 582970 352102
rect 583026 352046 583094 352102
rect 583150 352046 583218 352102
rect 583274 352046 583342 352102
rect 583398 352046 597456 352102
rect 597512 352046 597580 352102
rect 597636 352046 597704 352102
rect 597760 352046 597828 352102
rect 597884 352046 597980 352102
rect -1916 351978 597980 352046
rect -1916 351922 -1820 351978
rect -1764 351922 -1696 351978
rect -1640 351922 -1572 351978
rect -1516 351922 -1448 351978
rect -1392 351922 6970 351978
rect 7026 351922 7094 351978
rect 7150 351922 7218 351978
rect 7274 351922 7342 351978
rect 7398 351922 24970 351978
rect 25026 351922 25094 351978
rect 25150 351922 25218 351978
rect 25274 351922 25342 351978
rect 25398 351922 42970 351978
rect 43026 351922 43094 351978
rect 43150 351922 43218 351978
rect 43274 351922 43342 351978
rect 43398 351922 60970 351978
rect 61026 351922 61094 351978
rect 61150 351922 61218 351978
rect 61274 351922 61342 351978
rect 61398 351922 78970 351978
rect 79026 351922 79094 351978
rect 79150 351922 79218 351978
rect 79274 351922 79342 351978
rect 79398 351922 96970 351978
rect 97026 351922 97094 351978
rect 97150 351922 97218 351978
rect 97274 351922 97342 351978
rect 97398 351922 132970 351978
rect 133026 351922 133094 351978
rect 133150 351922 133218 351978
rect 133274 351922 133342 351978
rect 133398 351922 150970 351978
rect 151026 351922 151094 351978
rect 151150 351922 151218 351978
rect 151274 351922 151342 351978
rect 151398 351922 168970 351978
rect 169026 351922 169094 351978
rect 169150 351922 169218 351978
rect 169274 351922 169342 351978
rect 169398 351922 186970 351978
rect 187026 351922 187094 351978
rect 187150 351922 187218 351978
rect 187274 351922 187342 351978
rect 187398 351922 222970 351978
rect 223026 351922 223094 351978
rect 223150 351922 223218 351978
rect 223274 351922 223342 351978
rect 223398 351922 240970 351978
rect 241026 351922 241094 351978
rect 241150 351922 241218 351978
rect 241274 351922 241342 351978
rect 241398 351922 258970 351978
rect 259026 351922 259094 351978
rect 259150 351922 259218 351978
rect 259274 351922 259342 351978
rect 259398 351922 276970 351978
rect 277026 351922 277094 351978
rect 277150 351922 277218 351978
rect 277274 351922 277342 351978
rect 277398 351922 312970 351978
rect 313026 351922 313094 351978
rect 313150 351922 313218 351978
rect 313274 351922 313342 351978
rect 313398 351922 330970 351978
rect 331026 351922 331094 351978
rect 331150 351922 331218 351978
rect 331274 351922 331342 351978
rect 331398 351922 348970 351978
rect 349026 351922 349094 351978
rect 349150 351922 349218 351978
rect 349274 351922 349342 351978
rect 349398 351922 366970 351978
rect 367026 351922 367094 351978
rect 367150 351922 367218 351978
rect 367274 351922 367342 351978
rect 367398 351922 402970 351978
rect 403026 351922 403094 351978
rect 403150 351922 403218 351978
rect 403274 351922 403342 351978
rect 403398 351922 420970 351978
rect 421026 351922 421094 351978
rect 421150 351922 421218 351978
rect 421274 351922 421342 351978
rect 421398 351922 438970 351978
rect 439026 351922 439094 351978
rect 439150 351922 439218 351978
rect 439274 351922 439342 351978
rect 439398 351922 456970 351978
rect 457026 351922 457094 351978
rect 457150 351922 457218 351978
rect 457274 351922 457342 351978
rect 457398 351922 492970 351978
rect 493026 351922 493094 351978
rect 493150 351922 493218 351978
rect 493274 351922 493342 351978
rect 493398 351922 510970 351978
rect 511026 351922 511094 351978
rect 511150 351922 511218 351978
rect 511274 351922 511342 351978
rect 511398 351922 528970 351978
rect 529026 351922 529094 351978
rect 529150 351922 529218 351978
rect 529274 351922 529342 351978
rect 529398 351922 546970 351978
rect 547026 351922 547094 351978
rect 547150 351922 547218 351978
rect 547274 351922 547342 351978
rect 547398 351922 564970 351978
rect 565026 351922 565094 351978
rect 565150 351922 565218 351978
rect 565274 351922 565342 351978
rect 565398 351922 582970 351978
rect 583026 351922 583094 351978
rect 583150 351922 583218 351978
rect 583274 351922 583342 351978
rect 583398 351922 597456 351978
rect 597512 351922 597580 351978
rect 597636 351922 597704 351978
rect 597760 351922 597828 351978
rect 597884 351922 597980 351978
rect -1916 351826 597980 351922
rect -1916 346350 597980 346446
rect -1916 346294 -860 346350
rect -804 346294 -736 346350
rect -680 346294 -612 346350
rect -556 346294 -488 346350
rect -432 346294 3250 346350
rect 3306 346294 3374 346350
rect 3430 346294 3498 346350
rect 3554 346294 3622 346350
rect 3678 346294 21250 346350
rect 21306 346294 21374 346350
rect 21430 346294 21498 346350
rect 21554 346294 21622 346350
rect 21678 346294 39250 346350
rect 39306 346294 39374 346350
rect 39430 346294 39498 346350
rect 39554 346294 39622 346350
rect 39678 346294 57250 346350
rect 57306 346294 57374 346350
rect 57430 346294 57498 346350
rect 57554 346294 57622 346350
rect 57678 346294 93250 346350
rect 93306 346294 93374 346350
rect 93430 346294 93498 346350
rect 93554 346294 93622 346350
rect 93678 346294 111250 346350
rect 111306 346294 111374 346350
rect 111430 346294 111498 346350
rect 111554 346294 111622 346350
rect 111678 346294 129250 346350
rect 129306 346294 129374 346350
rect 129430 346294 129498 346350
rect 129554 346294 129622 346350
rect 129678 346294 147250 346350
rect 147306 346294 147374 346350
rect 147430 346294 147498 346350
rect 147554 346294 147622 346350
rect 147678 346294 183250 346350
rect 183306 346294 183374 346350
rect 183430 346294 183498 346350
rect 183554 346294 183622 346350
rect 183678 346294 201250 346350
rect 201306 346294 201374 346350
rect 201430 346294 201498 346350
rect 201554 346294 201622 346350
rect 201678 346294 219250 346350
rect 219306 346294 219374 346350
rect 219430 346294 219498 346350
rect 219554 346294 219622 346350
rect 219678 346294 237250 346350
rect 237306 346294 237374 346350
rect 237430 346294 237498 346350
rect 237554 346294 237622 346350
rect 237678 346294 273250 346350
rect 273306 346294 273374 346350
rect 273430 346294 273498 346350
rect 273554 346294 273622 346350
rect 273678 346294 291250 346350
rect 291306 346294 291374 346350
rect 291430 346294 291498 346350
rect 291554 346294 291622 346350
rect 291678 346294 309250 346350
rect 309306 346294 309374 346350
rect 309430 346294 309498 346350
rect 309554 346294 309622 346350
rect 309678 346294 327250 346350
rect 327306 346294 327374 346350
rect 327430 346294 327498 346350
rect 327554 346294 327622 346350
rect 327678 346294 363250 346350
rect 363306 346294 363374 346350
rect 363430 346294 363498 346350
rect 363554 346294 363622 346350
rect 363678 346294 381250 346350
rect 381306 346294 381374 346350
rect 381430 346294 381498 346350
rect 381554 346294 381622 346350
rect 381678 346294 399250 346350
rect 399306 346294 399374 346350
rect 399430 346294 399498 346350
rect 399554 346294 399622 346350
rect 399678 346294 417250 346350
rect 417306 346294 417374 346350
rect 417430 346294 417498 346350
rect 417554 346294 417622 346350
rect 417678 346294 453250 346350
rect 453306 346294 453374 346350
rect 453430 346294 453498 346350
rect 453554 346294 453622 346350
rect 453678 346294 471250 346350
rect 471306 346294 471374 346350
rect 471430 346294 471498 346350
rect 471554 346294 471622 346350
rect 471678 346294 489250 346350
rect 489306 346294 489374 346350
rect 489430 346294 489498 346350
rect 489554 346294 489622 346350
rect 489678 346294 507250 346350
rect 507306 346294 507374 346350
rect 507430 346294 507498 346350
rect 507554 346294 507622 346350
rect 507678 346294 543250 346350
rect 543306 346294 543374 346350
rect 543430 346294 543498 346350
rect 543554 346294 543622 346350
rect 543678 346294 561250 346350
rect 561306 346294 561374 346350
rect 561430 346294 561498 346350
rect 561554 346294 561622 346350
rect 561678 346294 579250 346350
rect 579306 346294 579374 346350
rect 579430 346294 579498 346350
rect 579554 346294 579622 346350
rect 579678 346294 596496 346350
rect 596552 346294 596620 346350
rect 596676 346294 596744 346350
rect 596800 346294 596868 346350
rect 596924 346294 597980 346350
rect -1916 346226 597980 346294
rect -1916 346170 -860 346226
rect -804 346170 -736 346226
rect -680 346170 -612 346226
rect -556 346170 -488 346226
rect -432 346170 3250 346226
rect 3306 346170 3374 346226
rect 3430 346170 3498 346226
rect 3554 346170 3622 346226
rect 3678 346170 21250 346226
rect 21306 346170 21374 346226
rect 21430 346170 21498 346226
rect 21554 346170 21622 346226
rect 21678 346170 39250 346226
rect 39306 346170 39374 346226
rect 39430 346170 39498 346226
rect 39554 346170 39622 346226
rect 39678 346170 57250 346226
rect 57306 346170 57374 346226
rect 57430 346170 57498 346226
rect 57554 346170 57622 346226
rect 57678 346170 93250 346226
rect 93306 346170 93374 346226
rect 93430 346170 93498 346226
rect 93554 346170 93622 346226
rect 93678 346170 111250 346226
rect 111306 346170 111374 346226
rect 111430 346170 111498 346226
rect 111554 346170 111622 346226
rect 111678 346170 129250 346226
rect 129306 346170 129374 346226
rect 129430 346170 129498 346226
rect 129554 346170 129622 346226
rect 129678 346170 147250 346226
rect 147306 346170 147374 346226
rect 147430 346170 147498 346226
rect 147554 346170 147622 346226
rect 147678 346170 183250 346226
rect 183306 346170 183374 346226
rect 183430 346170 183498 346226
rect 183554 346170 183622 346226
rect 183678 346170 201250 346226
rect 201306 346170 201374 346226
rect 201430 346170 201498 346226
rect 201554 346170 201622 346226
rect 201678 346170 219250 346226
rect 219306 346170 219374 346226
rect 219430 346170 219498 346226
rect 219554 346170 219622 346226
rect 219678 346170 237250 346226
rect 237306 346170 237374 346226
rect 237430 346170 237498 346226
rect 237554 346170 237622 346226
rect 237678 346170 273250 346226
rect 273306 346170 273374 346226
rect 273430 346170 273498 346226
rect 273554 346170 273622 346226
rect 273678 346170 291250 346226
rect 291306 346170 291374 346226
rect 291430 346170 291498 346226
rect 291554 346170 291622 346226
rect 291678 346170 309250 346226
rect 309306 346170 309374 346226
rect 309430 346170 309498 346226
rect 309554 346170 309622 346226
rect 309678 346170 327250 346226
rect 327306 346170 327374 346226
rect 327430 346170 327498 346226
rect 327554 346170 327622 346226
rect 327678 346170 363250 346226
rect 363306 346170 363374 346226
rect 363430 346170 363498 346226
rect 363554 346170 363622 346226
rect 363678 346170 381250 346226
rect 381306 346170 381374 346226
rect 381430 346170 381498 346226
rect 381554 346170 381622 346226
rect 381678 346170 399250 346226
rect 399306 346170 399374 346226
rect 399430 346170 399498 346226
rect 399554 346170 399622 346226
rect 399678 346170 417250 346226
rect 417306 346170 417374 346226
rect 417430 346170 417498 346226
rect 417554 346170 417622 346226
rect 417678 346170 453250 346226
rect 453306 346170 453374 346226
rect 453430 346170 453498 346226
rect 453554 346170 453622 346226
rect 453678 346170 471250 346226
rect 471306 346170 471374 346226
rect 471430 346170 471498 346226
rect 471554 346170 471622 346226
rect 471678 346170 489250 346226
rect 489306 346170 489374 346226
rect 489430 346170 489498 346226
rect 489554 346170 489622 346226
rect 489678 346170 507250 346226
rect 507306 346170 507374 346226
rect 507430 346170 507498 346226
rect 507554 346170 507622 346226
rect 507678 346170 543250 346226
rect 543306 346170 543374 346226
rect 543430 346170 543498 346226
rect 543554 346170 543622 346226
rect 543678 346170 561250 346226
rect 561306 346170 561374 346226
rect 561430 346170 561498 346226
rect 561554 346170 561622 346226
rect 561678 346170 579250 346226
rect 579306 346170 579374 346226
rect 579430 346170 579498 346226
rect 579554 346170 579622 346226
rect 579678 346170 596496 346226
rect 596552 346170 596620 346226
rect 596676 346170 596744 346226
rect 596800 346170 596868 346226
rect 596924 346170 597980 346226
rect -1916 346102 597980 346170
rect -1916 346046 -860 346102
rect -804 346046 -736 346102
rect -680 346046 -612 346102
rect -556 346046 -488 346102
rect -432 346046 3250 346102
rect 3306 346046 3374 346102
rect 3430 346046 3498 346102
rect 3554 346046 3622 346102
rect 3678 346046 21250 346102
rect 21306 346046 21374 346102
rect 21430 346046 21498 346102
rect 21554 346046 21622 346102
rect 21678 346046 39250 346102
rect 39306 346046 39374 346102
rect 39430 346046 39498 346102
rect 39554 346046 39622 346102
rect 39678 346046 57250 346102
rect 57306 346046 57374 346102
rect 57430 346046 57498 346102
rect 57554 346046 57622 346102
rect 57678 346046 93250 346102
rect 93306 346046 93374 346102
rect 93430 346046 93498 346102
rect 93554 346046 93622 346102
rect 93678 346046 111250 346102
rect 111306 346046 111374 346102
rect 111430 346046 111498 346102
rect 111554 346046 111622 346102
rect 111678 346046 129250 346102
rect 129306 346046 129374 346102
rect 129430 346046 129498 346102
rect 129554 346046 129622 346102
rect 129678 346046 147250 346102
rect 147306 346046 147374 346102
rect 147430 346046 147498 346102
rect 147554 346046 147622 346102
rect 147678 346046 183250 346102
rect 183306 346046 183374 346102
rect 183430 346046 183498 346102
rect 183554 346046 183622 346102
rect 183678 346046 201250 346102
rect 201306 346046 201374 346102
rect 201430 346046 201498 346102
rect 201554 346046 201622 346102
rect 201678 346046 219250 346102
rect 219306 346046 219374 346102
rect 219430 346046 219498 346102
rect 219554 346046 219622 346102
rect 219678 346046 237250 346102
rect 237306 346046 237374 346102
rect 237430 346046 237498 346102
rect 237554 346046 237622 346102
rect 237678 346046 273250 346102
rect 273306 346046 273374 346102
rect 273430 346046 273498 346102
rect 273554 346046 273622 346102
rect 273678 346046 291250 346102
rect 291306 346046 291374 346102
rect 291430 346046 291498 346102
rect 291554 346046 291622 346102
rect 291678 346046 309250 346102
rect 309306 346046 309374 346102
rect 309430 346046 309498 346102
rect 309554 346046 309622 346102
rect 309678 346046 327250 346102
rect 327306 346046 327374 346102
rect 327430 346046 327498 346102
rect 327554 346046 327622 346102
rect 327678 346046 363250 346102
rect 363306 346046 363374 346102
rect 363430 346046 363498 346102
rect 363554 346046 363622 346102
rect 363678 346046 381250 346102
rect 381306 346046 381374 346102
rect 381430 346046 381498 346102
rect 381554 346046 381622 346102
rect 381678 346046 399250 346102
rect 399306 346046 399374 346102
rect 399430 346046 399498 346102
rect 399554 346046 399622 346102
rect 399678 346046 417250 346102
rect 417306 346046 417374 346102
rect 417430 346046 417498 346102
rect 417554 346046 417622 346102
rect 417678 346046 453250 346102
rect 453306 346046 453374 346102
rect 453430 346046 453498 346102
rect 453554 346046 453622 346102
rect 453678 346046 471250 346102
rect 471306 346046 471374 346102
rect 471430 346046 471498 346102
rect 471554 346046 471622 346102
rect 471678 346046 489250 346102
rect 489306 346046 489374 346102
rect 489430 346046 489498 346102
rect 489554 346046 489622 346102
rect 489678 346046 507250 346102
rect 507306 346046 507374 346102
rect 507430 346046 507498 346102
rect 507554 346046 507622 346102
rect 507678 346046 543250 346102
rect 543306 346046 543374 346102
rect 543430 346046 543498 346102
rect 543554 346046 543622 346102
rect 543678 346046 561250 346102
rect 561306 346046 561374 346102
rect 561430 346046 561498 346102
rect 561554 346046 561622 346102
rect 561678 346046 579250 346102
rect 579306 346046 579374 346102
rect 579430 346046 579498 346102
rect 579554 346046 579622 346102
rect 579678 346046 596496 346102
rect 596552 346046 596620 346102
rect 596676 346046 596744 346102
rect 596800 346046 596868 346102
rect 596924 346046 597980 346102
rect -1916 345978 597980 346046
rect -1916 345922 -860 345978
rect -804 345922 -736 345978
rect -680 345922 -612 345978
rect -556 345922 -488 345978
rect -432 345922 3250 345978
rect 3306 345922 3374 345978
rect 3430 345922 3498 345978
rect 3554 345922 3622 345978
rect 3678 345922 21250 345978
rect 21306 345922 21374 345978
rect 21430 345922 21498 345978
rect 21554 345922 21622 345978
rect 21678 345922 39250 345978
rect 39306 345922 39374 345978
rect 39430 345922 39498 345978
rect 39554 345922 39622 345978
rect 39678 345922 57250 345978
rect 57306 345922 57374 345978
rect 57430 345922 57498 345978
rect 57554 345922 57622 345978
rect 57678 345922 93250 345978
rect 93306 345922 93374 345978
rect 93430 345922 93498 345978
rect 93554 345922 93622 345978
rect 93678 345922 111250 345978
rect 111306 345922 111374 345978
rect 111430 345922 111498 345978
rect 111554 345922 111622 345978
rect 111678 345922 129250 345978
rect 129306 345922 129374 345978
rect 129430 345922 129498 345978
rect 129554 345922 129622 345978
rect 129678 345922 147250 345978
rect 147306 345922 147374 345978
rect 147430 345922 147498 345978
rect 147554 345922 147622 345978
rect 147678 345922 183250 345978
rect 183306 345922 183374 345978
rect 183430 345922 183498 345978
rect 183554 345922 183622 345978
rect 183678 345922 201250 345978
rect 201306 345922 201374 345978
rect 201430 345922 201498 345978
rect 201554 345922 201622 345978
rect 201678 345922 219250 345978
rect 219306 345922 219374 345978
rect 219430 345922 219498 345978
rect 219554 345922 219622 345978
rect 219678 345922 237250 345978
rect 237306 345922 237374 345978
rect 237430 345922 237498 345978
rect 237554 345922 237622 345978
rect 237678 345922 273250 345978
rect 273306 345922 273374 345978
rect 273430 345922 273498 345978
rect 273554 345922 273622 345978
rect 273678 345922 291250 345978
rect 291306 345922 291374 345978
rect 291430 345922 291498 345978
rect 291554 345922 291622 345978
rect 291678 345922 309250 345978
rect 309306 345922 309374 345978
rect 309430 345922 309498 345978
rect 309554 345922 309622 345978
rect 309678 345922 327250 345978
rect 327306 345922 327374 345978
rect 327430 345922 327498 345978
rect 327554 345922 327622 345978
rect 327678 345922 363250 345978
rect 363306 345922 363374 345978
rect 363430 345922 363498 345978
rect 363554 345922 363622 345978
rect 363678 345922 381250 345978
rect 381306 345922 381374 345978
rect 381430 345922 381498 345978
rect 381554 345922 381622 345978
rect 381678 345922 399250 345978
rect 399306 345922 399374 345978
rect 399430 345922 399498 345978
rect 399554 345922 399622 345978
rect 399678 345922 417250 345978
rect 417306 345922 417374 345978
rect 417430 345922 417498 345978
rect 417554 345922 417622 345978
rect 417678 345922 453250 345978
rect 453306 345922 453374 345978
rect 453430 345922 453498 345978
rect 453554 345922 453622 345978
rect 453678 345922 471250 345978
rect 471306 345922 471374 345978
rect 471430 345922 471498 345978
rect 471554 345922 471622 345978
rect 471678 345922 489250 345978
rect 489306 345922 489374 345978
rect 489430 345922 489498 345978
rect 489554 345922 489622 345978
rect 489678 345922 507250 345978
rect 507306 345922 507374 345978
rect 507430 345922 507498 345978
rect 507554 345922 507622 345978
rect 507678 345922 543250 345978
rect 543306 345922 543374 345978
rect 543430 345922 543498 345978
rect 543554 345922 543622 345978
rect 543678 345922 561250 345978
rect 561306 345922 561374 345978
rect 561430 345922 561498 345978
rect 561554 345922 561622 345978
rect 561678 345922 579250 345978
rect 579306 345922 579374 345978
rect 579430 345922 579498 345978
rect 579554 345922 579622 345978
rect 579678 345922 596496 345978
rect 596552 345922 596620 345978
rect 596676 345922 596744 345978
rect 596800 345922 596868 345978
rect 596924 345922 597980 345978
rect -1916 345826 597980 345922
rect -1916 334350 597980 334446
rect -1916 334294 -1820 334350
rect -1764 334294 -1696 334350
rect -1640 334294 -1572 334350
rect -1516 334294 -1448 334350
rect -1392 334294 6970 334350
rect 7026 334294 7094 334350
rect 7150 334294 7218 334350
rect 7274 334294 7342 334350
rect 7398 334294 24970 334350
rect 25026 334294 25094 334350
rect 25150 334294 25218 334350
rect 25274 334294 25342 334350
rect 25398 334294 42970 334350
rect 43026 334294 43094 334350
rect 43150 334294 43218 334350
rect 43274 334294 43342 334350
rect 43398 334294 60970 334350
rect 61026 334294 61094 334350
rect 61150 334294 61218 334350
rect 61274 334294 61342 334350
rect 61398 334294 78970 334350
rect 79026 334294 79094 334350
rect 79150 334294 79218 334350
rect 79274 334294 79342 334350
rect 79398 334294 96970 334350
rect 97026 334294 97094 334350
rect 97150 334294 97218 334350
rect 97274 334294 97342 334350
rect 97398 334294 132970 334350
rect 133026 334294 133094 334350
rect 133150 334294 133218 334350
rect 133274 334294 133342 334350
rect 133398 334294 150970 334350
rect 151026 334294 151094 334350
rect 151150 334294 151218 334350
rect 151274 334294 151342 334350
rect 151398 334294 168970 334350
rect 169026 334294 169094 334350
rect 169150 334294 169218 334350
rect 169274 334294 169342 334350
rect 169398 334294 186970 334350
rect 187026 334294 187094 334350
rect 187150 334294 187218 334350
rect 187274 334294 187342 334350
rect 187398 334294 222970 334350
rect 223026 334294 223094 334350
rect 223150 334294 223218 334350
rect 223274 334294 223342 334350
rect 223398 334294 240970 334350
rect 241026 334294 241094 334350
rect 241150 334294 241218 334350
rect 241274 334294 241342 334350
rect 241398 334294 258970 334350
rect 259026 334294 259094 334350
rect 259150 334294 259218 334350
rect 259274 334294 259342 334350
rect 259398 334294 276970 334350
rect 277026 334294 277094 334350
rect 277150 334294 277218 334350
rect 277274 334294 277342 334350
rect 277398 334294 312970 334350
rect 313026 334294 313094 334350
rect 313150 334294 313218 334350
rect 313274 334294 313342 334350
rect 313398 334294 330970 334350
rect 331026 334294 331094 334350
rect 331150 334294 331218 334350
rect 331274 334294 331342 334350
rect 331398 334294 348970 334350
rect 349026 334294 349094 334350
rect 349150 334294 349218 334350
rect 349274 334294 349342 334350
rect 349398 334294 366970 334350
rect 367026 334294 367094 334350
rect 367150 334294 367218 334350
rect 367274 334294 367342 334350
rect 367398 334294 402970 334350
rect 403026 334294 403094 334350
rect 403150 334294 403218 334350
rect 403274 334294 403342 334350
rect 403398 334294 420970 334350
rect 421026 334294 421094 334350
rect 421150 334294 421218 334350
rect 421274 334294 421342 334350
rect 421398 334294 438970 334350
rect 439026 334294 439094 334350
rect 439150 334294 439218 334350
rect 439274 334294 439342 334350
rect 439398 334294 456970 334350
rect 457026 334294 457094 334350
rect 457150 334294 457218 334350
rect 457274 334294 457342 334350
rect 457398 334294 492970 334350
rect 493026 334294 493094 334350
rect 493150 334294 493218 334350
rect 493274 334294 493342 334350
rect 493398 334294 510970 334350
rect 511026 334294 511094 334350
rect 511150 334294 511218 334350
rect 511274 334294 511342 334350
rect 511398 334294 528970 334350
rect 529026 334294 529094 334350
rect 529150 334294 529218 334350
rect 529274 334294 529342 334350
rect 529398 334294 546970 334350
rect 547026 334294 547094 334350
rect 547150 334294 547218 334350
rect 547274 334294 547342 334350
rect 547398 334294 564970 334350
rect 565026 334294 565094 334350
rect 565150 334294 565218 334350
rect 565274 334294 565342 334350
rect 565398 334294 582970 334350
rect 583026 334294 583094 334350
rect 583150 334294 583218 334350
rect 583274 334294 583342 334350
rect 583398 334294 597456 334350
rect 597512 334294 597580 334350
rect 597636 334294 597704 334350
rect 597760 334294 597828 334350
rect 597884 334294 597980 334350
rect -1916 334226 597980 334294
rect -1916 334170 -1820 334226
rect -1764 334170 -1696 334226
rect -1640 334170 -1572 334226
rect -1516 334170 -1448 334226
rect -1392 334170 6970 334226
rect 7026 334170 7094 334226
rect 7150 334170 7218 334226
rect 7274 334170 7342 334226
rect 7398 334170 24970 334226
rect 25026 334170 25094 334226
rect 25150 334170 25218 334226
rect 25274 334170 25342 334226
rect 25398 334170 42970 334226
rect 43026 334170 43094 334226
rect 43150 334170 43218 334226
rect 43274 334170 43342 334226
rect 43398 334170 60970 334226
rect 61026 334170 61094 334226
rect 61150 334170 61218 334226
rect 61274 334170 61342 334226
rect 61398 334170 78970 334226
rect 79026 334170 79094 334226
rect 79150 334170 79218 334226
rect 79274 334170 79342 334226
rect 79398 334170 96970 334226
rect 97026 334170 97094 334226
rect 97150 334170 97218 334226
rect 97274 334170 97342 334226
rect 97398 334170 132970 334226
rect 133026 334170 133094 334226
rect 133150 334170 133218 334226
rect 133274 334170 133342 334226
rect 133398 334170 150970 334226
rect 151026 334170 151094 334226
rect 151150 334170 151218 334226
rect 151274 334170 151342 334226
rect 151398 334170 168970 334226
rect 169026 334170 169094 334226
rect 169150 334170 169218 334226
rect 169274 334170 169342 334226
rect 169398 334170 186970 334226
rect 187026 334170 187094 334226
rect 187150 334170 187218 334226
rect 187274 334170 187342 334226
rect 187398 334170 222970 334226
rect 223026 334170 223094 334226
rect 223150 334170 223218 334226
rect 223274 334170 223342 334226
rect 223398 334170 240970 334226
rect 241026 334170 241094 334226
rect 241150 334170 241218 334226
rect 241274 334170 241342 334226
rect 241398 334170 258970 334226
rect 259026 334170 259094 334226
rect 259150 334170 259218 334226
rect 259274 334170 259342 334226
rect 259398 334170 276970 334226
rect 277026 334170 277094 334226
rect 277150 334170 277218 334226
rect 277274 334170 277342 334226
rect 277398 334170 312970 334226
rect 313026 334170 313094 334226
rect 313150 334170 313218 334226
rect 313274 334170 313342 334226
rect 313398 334170 330970 334226
rect 331026 334170 331094 334226
rect 331150 334170 331218 334226
rect 331274 334170 331342 334226
rect 331398 334170 348970 334226
rect 349026 334170 349094 334226
rect 349150 334170 349218 334226
rect 349274 334170 349342 334226
rect 349398 334170 366970 334226
rect 367026 334170 367094 334226
rect 367150 334170 367218 334226
rect 367274 334170 367342 334226
rect 367398 334170 402970 334226
rect 403026 334170 403094 334226
rect 403150 334170 403218 334226
rect 403274 334170 403342 334226
rect 403398 334170 420970 334226
rect 421026 334170 421094 334226
rect 421150 334170 421218 334226
rect 421274 334170 421342 334226
rect 421398 334170 438970 334226
rect 439026 334170 439094 334226
rect 439150 334170 439218 334226
rect 439274 334170 439342 334226
rect 439398 334170 456970 334226
rect 457026 334170 457094 334226
rect 457150 334170 457218 334226
rect 457274 334170 457342 334226
rect 457398 334170 492970 334226
rect 493026 334170 493094 334226
rect 493150 334170 493218 334226
rect 493274 334170 493342 334226
rect 493398 334170 510970 334226
rect 511026 334170 511094 334226
rect 511150 334170 511218 334226
rect 511274 334170 511342 334226
rect 511398 334170 528970 334226
rect 529026 334170 529094 334226
rect 529150 334170 529218 334226
rect 529274 334170 529342 334226
rect 529398 334170 546970 334226
rect 547026 334170 547094 334226
rect 547150 334170 547218 334226
rect 547274 334170 547342 334226
rect 547398 334170 564970 334226
rect 565026 334170 565094 334226
rect 565150 334170 565218 334226
rect 565274 334170 565342 334226
rect 565398 334170 582970 334226
rect 583026 334170 583094 334226
rect 583150 334170 583218 334226
rect 583274 334170 583342 334226
rect 583398 334170 597456 334226
rect 597512 334170 597580 334226
rect 597636 334170 597704 334226
rect 597760 334170 597828 334226
rect 597884 334170 597980 334226
rect -1916 334102 597980 334170
rect -1916 334046 -1820 334102
rect -1764 334046 -1696 334102
rect -1640 334046 -1572 334102
rect -1516 334046 -1448 334102
rect -1392 334046 6970 334102
rect 7026 334046 7094 334102
rect 7150 334046 7218 334102
rect 7274 334046 7342 334102
rect 7398 334046 24970 334102
rect 25026 334046 25094 334102
rect 25150 334046 25218 334102
rect 25274 334046 25342 334102
rect 25398 334046 42970 334102
rect 43026 334046 43094 334102
rect 43150 334046 43218 334102
rect 43274 334046 43342 334102
rect 43398 334046 60970 334102
rect 61026 334046 61094 334102
rect 61150 334046 61218 334102
rect 61274 334046 61342 334102
rect 61398 334046 78970 334102
rect 79026 334046 79094 334102
rect 79150 334046 79218 334102
rect 79274 334046 79342 334102
rect 79398 334046 96970 334102
rect 97026 334046 97094 334102
rect 97150 334046 97218 334102
rect 97274 334046 97342 334102
rect 97398 334046 132970 334102
rect 133026 334046 133094 334102
rect 133150 334046 133218 334102
rect 133274 334046 133342 334102
rect 133398 334046 150970 334102
rect 151026 334046 151094 334102
rect 151150 334046 151218 334102
rect 151274 334046 151342 334102
rect 151398 334046 168970 334102
rect 169026 334046 169094 334102
rect 169150 334046 169218 334102
rect 169274 334046 169342 334102
rect 169398 334046 186970 334102
rect 187026 334046 187094 334102
rect 187150 334046 187218 334102
rect 187274 334046 187342 334102
rect 187398 334046 222970 334102
rect 223026 334046 223094 334102
rect 223150 334046 223218 334102
rect 223274 334046 223342 334102
rect 223398 334046 240970 334102
rect 241026 334046 241094 334102
rect 241150 334046 241218 334102
rect 241274 334046 241342 334102
rect 241398 334046 258970 334102
rect 259026 334046 259094 334102
rect 259150 334046 259218 334102
rect 259274 334046 259342 334102
rect 259398 334046 276970 334102
rect 277026 334046 277094 334102
rect 277150 334046 277218 334102
rect 277274 334046 277342 334102
rect 277398 334046 312970 334102
rect 313026 334046 313094 334102
rect 313150 334046 313218 334102
rect 313274 334046 313342 334102
rect 313398 334046 330970 334102
rect 331026 334046 331094 334102
rect 331150 334046 331218 334102
rect 331274 334046 331342 334102
rect 331398 334046 348970 334102
rect 349026 334046 349094 334102
rect 349150 334046 349218 334102
rect 349274 334046 349342 334102
rect 349398 334046 366970 334102
rect 367026 334046 367094 334102
rect 367150 334046 367218 334102
rect 367274 334046 367342 334102
rect 367398 334046 402970 334102
rect 403026 334046 403094 334102
rect 403150 334046 403218 334102
rect 403274 334046 403342 334102
rect 403398 334046 420970 334102
rect 421026 334046 421094 334102
rect 421150 334046 421218 334102
rect 421274 334046 421342 334102
rect 421398 334046 438970 334102
rect 439026 334046 439094 334102
rect 439150 334046 439218 334102
rect 439274 334046 439342 334102
rect 439398 334046 456970 334102
rect 457026 334046 457094 334102
rect 457150 334046 457218 334102
rect 457274 334046 457342 334102
rect 457398 334046 492970 334102
rect 493026 334046 493094 334102
rect 493150 334046 493218 334102
rect 493274 334046 493342 334102
rect 493398 334046 510970 334102
rect 511026 334046 511094 334102
rect 511150 334046 511218 334102
rect 511274 334046 511342 334102
rect 511398 334046 528970 334102
rect 529026 334046 529094 334102
rect 529150 334046 529218 334102
rect 529274 334046 529342 334102
rect 529398 334046 546970 334102
rect 547026 334046 547094 334102
rect 547150 334046 547218 334102
rect 547274 334046 547342 334102
rect 547398 334046 564970 334102
rect 565026 334046 565094 334102
rect 565150 334046 565218 334102
rect 565274 334046 565342 334102
rect 565398 334046 582970 334102
rect 583026 334046 583094 334102
rect 583150 334046 583218 334102
rect 583274 334046 583342 334102
rect 583398 334046 597456 334102
rect 597512 334046 597580 334102
rect 597636 334046 597704 334102
rect 597760 334046 597828 334102
rect 597884 334046 597980 334102
rect -1916 333978 597980 334046
rect -1916 333922 -1820 333978
rect -1764 333922 -1696 333978
rect -1640 333922 -1572 333978
rect -1516 333922 -1448 333978
rect -1392 333922 6970 333978
rect 7026 333922 7094 333978
rect 7150 333922 7218 333978
rect 7274 333922 7342 333978
rect 7398 333922 24970 333978
rect 25026 333922 25094 333978
rect 25150 333922 25218 333978
rect 25274 333922 25342 333978
rect 25398 333922 42970 333978
rect 43026 333922 43094 333978
rect 43150 333922 43218 333978
rect 43274 333922 43342 333978
rect 43398 333922 60970 333978
rect 61026 333922 61094 333978
rect 61150 333922 61218 333978
rect 61274 333922 61342 333978
rect 61398 333922 78970 333978
rect 79026 333922 79094 333978
rect 79150 333922 79218 333978
rect 79274 333922 79342 333978
rect 79398 333922 96970 333978
rect 97026 333922 97094 333978
rect 97150 333922 97218 333978
rect 97274 333922 97342 333978
rect 97398 333922 132970 333978
rect 133026 333922 133094 333978
rect 133150 333922 133218 333978
rect 133274 333922 133342 333978
rect 133398 333922 150970 333978
rect 151026 333922 151094 333978
rect 151150 333922 151218 333978
rect 151274 333922 151342 333978
rect 151398 333922 168970 333978
rect 169026 333922 169094 333978
rect 169150 333922 169218 333978
rect 169274 333922 169342 333978
rect 169398 333922 186970 333978
rect 187026 333922 187094 333978
rect 187150 333922 187218 333978
rect 187274 333922 187342 333978
rect 187398 333922 222970 333978
rect 223026 333922 223094 333978
rect 223150 333922 223218 333978
rect 223274 333922 223342 333978
rect 223398 333922 240970 333978
rect 241026 333922 241094 333978
rect 241150 333922 241218 333978
rect 241274 333922 241342 333978
rect 241398 333922 258970 333978
rect 259026 333922 259094 333978
rect 259150 333922 259218 333978
rect 259274 333922 259342 333978
rect 259398 333922 276970 333978
rect 277026 333922 277094 333978
rect 277150 333922 277218 333978
rect 277274 333922 277342 333978
rect 277398 333922 312970 333978
rect 313026 333922 313094 333978
rect 313150 333922 313218 333978
rect 313274 333922 313342 333978
rect 313398 333922 330970 333978
rect 331026 333922 331094 333978
rect 331150 333922 331218 333978
rect 331274 333922 331342 333978
rect 331398 333922 348970 333978
rect 349026 333922 349094 333978
rect 349150 333922 349218 333978
rect 349274 333922 349342 333978
rect 349398 333922 366970 333978
rect 367026 333922 367094 333978
rect 367150 333922 367218 333978
rect 367274 333922 367342 333978
rect 367398 333922 402970 333978
rect 403026 333922 403094 333978
rect 403150 333922 403218 333978
rect 403274 333922 403342 333978
rect 403398 333922 420970 333978
rect 421026 333922 421094 333978
rect 421150 333922 421218 333978
rect 421274 333922 421342 333978
rect 421398 333922 438970 333978
rect 439026 333922 439094 333978
rect 439150 333922 439218 333978
rect 439274 333922 439342 333978
rect 439398 333922 456970 333978
rect 457026 333922 457094 333978
rect 457150 333922 457218 333978
rect 457274 333922 457342 333978
rect 457398 333922 492970 333978
rect 493026 333922 493094 333978
rect 493150 333922 493218 333978
rect 493274 333922 493342 333978
rect 493398 333922 510970 333978
rect 511026 333922 511094 333978
rect 511150 333922 511218 333978
rect 511274 333922 511342 333978
rect 511398 333922 528970 333978
rect 529026 333922 529094 333978
rect 529150 333922 529218 333978
rect 529274 333922 529342 333978
rect 529398 333922 546970 333978
rect 547026 333922 547094 333978
rect 547150 333922 547218 333978
rect 547274 333922 547342 333978
rect 547398 333922 564970 333978
rect 565026 333922 565094 333978
rect 565150 333922 565218 333978
rect 565274 333922 565342 333978
rect 565398 333922 582970 333978
rect 583026 333922 583094 333978
rect 583150 333922 583218 333978
rect 583274 333922 583342 333978
rect 583398 333922 597456 333978
rect 597512 333922 597580 333978
rect 597636 333922 597704 333978
rect 597760 333922 597828 333978
rect 597884 333922 597980 333978
rect -1916 333826 597980 333922
rect -1916 328350 597980 328446
rect -1916 328294 -860 328350
rect -804 328294 -736 328350
rect -680 328294 -612 328350
rect -556 328294 -488 328350
rect -432 328294 3250 328350
rect 3306 328294 3374 328350
rect 3430 328294 3498 328350
rect 3554 328294 3622 328350
rect 3678 328294 21250 328350
rect 21306 328294 21374 328350
rect 21430 328294 21498 328350
rect 21554 328294 21622 328350
rect 21678 328294 39250 328350
rect 39306 328294 39374 328350
rect 39430 328294 39498 328350
rect 39554 328294 39622 328350
rect 39678 328294 57250 328350
rect 57306 328294 57374 328350
rect 57430 328294 57498 328350
rect 57554 328294 57622 328350
rect 57678 328294 93250 328350
rect 93306 328294 93374 328350
rect 93430 328294 93498 328350
rect 93554 328294 93622 328350
rect 93678 328294 111250 328350
rect 111306 328294 111374 328350
rect 111430 328294 111498 328350
rect 111554 328294 111622 328350
rect 111678 328294 129250 328350
rect 129306 328294 129374 328350
rect 129430 328294 129498 328350
rect 129554 328294 129622 328350
rect 129678 328294 147250 328350
rect 147306 328294 147374 328350
rect 147430 328294 147498 328350
rect 147554 328294 147622 328350
rect 147678 328294 183250 328350
rect 183306 328294 183374 328350
rect 183430 328294 183498 328350
rect 183554 328294 183622 328350
rect 183678 328294 201250 328350
rect 201306 328294 201374 328350
rect 201430 328294 201498 328350
rect 201554 328294 201622 328350
rect 201678 328294 219250 328350
rect 219306 328294 219374 328350
rect 219430 328294 219498 328350
rect 219554 328294 219622 328350
rect 219678 328294 237250 328350
rect 237306 328294 237374 328350
rect 237430 328294 237498 328350
rect 237554 328294 237622 328350
rect 237678 328294 273250 328350
rect 273306 328294 273374 328350
rect 273430 328294 273498 328350
rect 273554 328294 273622 328350
rect 273678 328294 291250 328350
rect 291306 328294 291374 328350
rect 291430 328294 291498 328350
rect 291554 328294 291622 328350
rect 291678 328294 309250 328350
rect 309306 328294 309374 328350
rect 309430 328294 309498 328350
rect 309554 328294 309622 328350
rect 309678 328294 327250 328350
rect 327306 328294 327374 328350
rect 327430 328294 327498 328350
rect 327554 328294 327622 328350
rect 327678 328294 363250 328350
rect 363306 328294 363374 328350
rect 363430 328294 363498 328350
rect 363554 328294 363622 328350
rect 363678 328294 381250 328350
rect 381306 328294 381374 328350
rect 381430 328294 381498 328350
rect 381554 328294 381622 328350
rect 381678 328294 399250 328350
rect 399306 328294 399374 328350
rect 399430 328294 399498 328350
rect 399554 328294 399622 328350
rect 399678 328294 417250 328350
rect 417306 328294 417374 328350
rect 417430 328294 417498 328350
rect 417554 328294 417622 328350
rect 417678 328294 453250 328350
rect 453306 328294 453374 328350
rect 453430 328294 453498 328350
rect 453554 328294 453622 328350
rect 453678 328294 471250 328350
rect 471306 328294 471374 328350
rect 471430 328294 471498 328350
rect 471554 328294 471622 328350
rect 471678 328294 489250 328350
rect 489306 328294 489374 328350
rect 489430 328294 489498 328350
rect 489554 328294 489622 328350
rect 489678 328294 507250 328350
rect 507306 328294 507374 328350
rect 507430 328294 507498 328350
rect 507554 328294 507622 328350
rect 507678 328294 543250 328350
rect 543306 328294 543374 328350
rect 543430 328294 543498 328350
rect 543554 328294 543622 328350
rect 543678 328294 561250 328350
rect 561306 328294 561374 328350
rect 561430 328294 561498 328350
rect 561554 328294 561622 328350
rect 561678 328294 579250 328350
rect 579306 328294 579374 328350
rect 579430 328294 579498 328350
rect 579554 328294 579622 328350
rect 579678 328294 596496 328350
rect 596552 328294 596620 328350
rect 596676 328294 596744 328350
rect 596800 328294 596868 328350
rect 596924 328294 597980 328350
rect -1916 328226 597980 328294
rect -1916 328170 -860 328226
rect -804 328170 -736 328226
rect -680 328170 -612 328226
rect -556 328170 -488 328226
rect -432 328170 3250 328226
rect 3306 328170 3374 328226
rect 3430 328170 3498 328226
rect 3554 328170 3622 328226
rect 3678 328170 21250 328226
rect 21306 328170 21374 328226
rect 21430 328170 21498 328226
rect 21554 328170 21622 328226
rect 21678 328170 39250 328226
rect 39306 328170 39374 328226
rect 39430 328170 39498 328226
rect 39554 328170 39622 328226
rect 39678 328170 57250 328226
rect 57306 328170 57374 328226
rect 57430 328170 57498 328226
rect 57554 328170 57622 328226
rect 57678 328170 93250 328226
rect 93306 328170 93374 328226
rect 93430 328170 93498 328226
rect 93554 328170 93622 328226
rect 93678 328170 111250 328226
rect 111306 328170 111374 328226
rect 111430 328170 111498 328226
rect 111554 328170 111622 328226
rect 111678 328170 129250 328226
rect 129306 328170 129374 328226
rect 129430 328170 129498 328226
rect 129554 328170 129622 328226
rect 129678 328170 147250 328226
rect 147306 328170 147374 328226
rect 147430 328170 147498 328226
rect 147554 328170 147622 328226
rect 147678 328170 183250 328226
rect 183306 328170 183374 328226
rect 183430 328170 183498 328226
rect 183554 328170 183622 328226
rect 183678 328170 201250 328226
rect 201306 328170 201374 328226
rect 201430 328170 201498 328226
rect 201554 328170 201622 328226
rect 201678 328170 219250 328226
rect 219306 328170 219374 328226
rect 219430 328170 219498 328226
rect 219554 328170 219622 328226
rect 219678 328170 237250 328226
rect 237306 328170 237374 328226
rect 237430 328170 237498 328226
rect 237554 328170 237622 328226
rect 237678 328170 273250 328226
rect 273306 328170 273374 328226
rect 273430 328170 273498 328226
rect 273554 328170 273622 328226
rect 273678 328170 291250 328226
rect 291306 328170 291374 328226
rect 291430 328170 291498 328226
rect 291554 328170 291622 328226
rect 291678 328170 309250 328226
rect 309306 328170 309374 328226
rect 309430 328170 309498 328226
rect 309554 328170 309622 328226
rect 309678 328170 327250 328226
rect 327306 328170 327374 328226
rect 327430 328170 327498 328226
rect 327554 328170 327622 328226
rect 327678 328170 363250 328226
rect 363306 328170 363374 328226
rect 363430 328170 363498 328226
rect 363554 328170 363622 328226
rect 363678 328170 381250 328226
rect 381306 328170 381374 328226
rect 381430 328170 381498 328226
rect 381554 328170 381622 328226
rect 381678 328170 399250 328226
rect 399306 328170 399374 328226
rect 399430 328170 399498 328226
rect 399554 328170 399622 328226
rect 399678 328170 417250 328226
rect 417306 328170 417374 328226
rect 417430 328170 417498 328226
rect 417554 328170 417622 328226
rect 417678 328170 453250 328226
rect 453306 328170 453374 328226
rect 453430 328170 453498 328226
rect 453554 328170 453622 328226
rect 453678 328170 471250 328226
rect 471306 328170 471374 328226
rect 471430 328170 471498 328226
rect 471554 328170 471622 328226
rect 471678 328170 489250 328226
rect 489306 328170 489374 328226
rect 489430 328170 489498 328226
rect 489554 328170 489622 328226
rect 489678 328170 507250 328226
rect 507306 328170 507374 328226
rect 507430 328170 507498 328226
rect 507554 328170 507622 328226
rect 507678 328170 543250 328226
rect 543306 328170 543374 328226
rect 543430 328170 543498 328226
rect 543554 328170 543622 328226
rect 543678 328170 561250 328226
rect 561306 328170 561374 328226
rect 561430 328170 561498 328226
rect 561554 328170 561622 328226
rect 561678 328170 579250 328226
rect 579306 328170 579374 328226
rect 579430 328170 579498 328226
rect 579554 328170 579622 328226
rect 579678 328170 596496 328226
rect 596552 328170 596620 328226
rect 596676 328170 596744 328226
rect 596800 328170 596868 328226
rect 596924 328170 597980 328226
rect -1916 328102 597980 328170
rect -1916 328046 -860 328102
rect -804 328046 -736 328102
rect -680 328046 -612 328102
rect -556 328046 -488 328102
rect -432 328046 3250 328102
rect 3306 328046 3374 328102
rect 3430 328046 3498 328102
rect 3554 328046 3622 328102
rect 3678 328046 21250 328102
rect 21306 328046 21374 328102
rect 21430 328046 21498 328102
rect 21554 328046 21622 328102
rect 21678 328046 39250 328102
rect 39306 328046 39374 328102
rect 39430 328046 39498 328102
rect 39554 328046 39622 328102
rect 39678 328046 57250 328102
rect 57306 328046 57374 328102
rect 57430 328046 57498 328102
rect 57554 328046 57622 328102
rect 57678 328046 93250 328102
rect 93306 328046 93374 328102
rect 93430 328046 93498 328102
rect 93554 328046 93622 328102
rect 93678 328046 111250 328102
rect 111306 328046 111374 328102
rect 111430 328046 111498 328102
rect 111554 328046 111622 328102
rect 111678 328046 129250 328102
rect 129306 328046 129374 328102
rect 129430 328046 129498 328102
rect 129554 328046 129622 328102
rect 129678 328046 147250 328102
rect 147306 328046 147374 328102
rect 147430 328046 147498 328102
rect 147554 328046 147622 328102
rect 147678 328046 183250 328102
rect 183306 328046 183374 328102
rect 183430 328046 183498 328102
rect 183554 328046 183622 328102
rect 183678 328046 201250 328102
rect 201306 328046 201374 328102
rect 201430 328046 201498 328102
rect 201554 328046 201622 328102
rect 201678 328046 219250 328102
rect 219306 328046 219374 328102
rect 219430 328046 219498 328102
rect 219554 328046 219622 328102
rect 219678 328046 237250 328102
rect 237306 328046 237374 328102
rect 237430 328046 237498 328102
rect 237554 328046 237622 328102
rect 237678 328046 273250 328102
rect 273306 328046 273374 328102
rect 273430 328046 273498 328102
rect 273554 328046 273622 328102
rect 273678 328046 291250 328102
rect 291306 328046 291374 328102
rect 291430 328046 291498 328102
rect 291554 328046 291622 328102
rect 291678 328046 309250 328102
rect 309306 328046 309374 328102
rect 309430 328046 309498 328102
rect 309554 328046 309622 328102
rect 309678 328046 327250 328102
rect 327306 328046 327374 328102
rect 327430 328046 327498 328102
rect 327554 328046 327622 328102
rect 327678 328046 363250 328102
rect 363306 328046 363374 328102
rect 363430 328046 363498 328102
rect 363554 328046 363622 328102
rect 363678 328046 381250 328102
rect 381306 328046 381374 328102
rect 381430 328046 381498 328102
rect 381554 328046 381622 328102
rect 381678 328046 399250 328102
rect 399306 328046 399374 328102
rect 399430 328046 399498 328102
rect 399554 328046 399622 328102
rect 399678 328046 417250 328102
rect 417306 328046 417374 328102
rect 417430 328046 417498 328102
rect 417554 328046 417622 328102
rect 417678 328046 453250 328102
rect 453306 328046 453374 328102
rect 453430 328046 453498 328102
rect 453554 328046 453622 328102
rect 453678 328046 471250 328102
rect 471306 328046 471374 328102
rect 471430 328046 471498 328102
rect 471554 328046 471622 328102
rect 471678 328046 489250 328102
rect 489306 328046 489374 328102
rect 489430 328046 489498 328102
rect 489554 328046 489622 328102
rect 489678 328046 507250 328102
rect 507306 328046 507374 328102
rect 507430 328046 507498 328102
rect 507554 328046 507622 328102
rect 507678 328046 543250 328102
rect 543306 328046 543374 328102
rect 543430 328046 543498 328102
rect 543554 328046 543622 328102
rect 543678 328046 561250 328102
rect 561306 328046 561374 328102
rect 561430 328046 561498 328102
rect 561554 328046 561622 328102
rect 561678 328046 579250 328102
rect 579306 328046 579374 328102
rect 579430 328046 579498 328102
rect 579554 328046 579622 328102
rect 579678 328046 596496 328102
rect 596552 328046 596620 328102
rect 596676 328046 596744 328102
rect 596800 328046 596868 328102
rect 596924 328046 597980 328102
rect -1916 327978 597980 328046
rect -1916 327922 -860 327978
rect -804 327922 -736 327978
rect -680 327922 -612 327978
rect -556 327922 -488 327978
rect -432 327922 3250 327978
rect 3306 327922 3374 327978
rect 3430 327922 3498 327978
rect 3554 327922 3622 327978
rect 3678 327922 21250 327978
rect 21306 327922 21374 327978
rect 21430 327922 21498 327978
rect 21554 327922 21622 327978
rect 21678 327922 39250 327978
rect 39306 327922 39374 327978
rect 39430 327922 39498 327978
rect 39554 327922 39622 327978
rect 39678 327922 57250 327978
rect 57306 327922 57374 327978
rect 57430 327922 57498 327978
rect 57554 327922 57622 327978
rect 57678 327922 93250 327978
rect 93306 327922 93374 327978
rect 93430 327922 93498 327978
rect 93554 327922 93622 327978
rect 93678 327922 111250 327978
rect 111306 327922 111374 327978
rect 111430 327922 111498 327978
rect 111554 327922 111622 327978
rect 111678 327922 129250 327978
rect 129306 327922 129374 327978
rect 129430 327922 129498 327978
rect 129554 327922 129622 327978
rect 129678 327922 147250 327978
rect 147306 327922 147374 327978
rect 147430 327922 147498 327978
rect 147554 327922 147622 327978
rect 147678 327922 183250 327978
rect 183306 327922 183374 327978
rect 183430 327922 183498 327978
rect 183554 327922 183622 327978
rect 183678 327922 201250 327978
rect 201306 327922 201374 327978
rect 201430 327922 201498 327978
rect 201554 327922 201622 327978
rect 201678 327922 219250 327978
rect 219306 327922 219374 327978
rect 219430 327922 219498 327978
rect 219554 327922 219622 327978
rect 219678 327922 237250 327978
rect 237306 327922 237374 327978
rect 237430 327922 237498 327978
rect 237554 327922 237622 327978
rect 237678 327922 273250 327978
rect 273306 327922 273374 327978
rect 273430 327922 273498 327978
rect 273554 327922 273622 327978
rect 273678 327922 291250 327978
rect 291306 327922 291374 327978
rect 291430 327922 291498 327978
rect 291554 327922 291622 327978
rect 291678 327922 309250 327978
rect 309306 327922 309374 327978
rect 309430 327922 309498 327978
rect 309554 327922 309622 327978
rect 309678 327922 327250 327978
rect 327306 327922 327374 327978
rect 327430 327922 327498 327978
rect 327554 327922 327622 327978
rect 327678 327922 363250 327978
rect 363306 327922 363374 327978
rect 363430 327922 363498 327978
rect 363554 327922 363622 327978
rect 363678 327922 381250 327978
rect 381306 327922 381374 327978
rect 381430 327922 381498 327978
rect 381554 327922 381622 327978
rect 381678 327922 399250 327978
rect 399306 327922 399374 327978
rect 399430 327922 399498 327978
rect 399554 327922 399622 327978
rect 399678 327922 417250 327978
rect 417306 327922 417374 327978
rect 417430 327922 417498 327978
rect 417554 327922 417622 327978
rect 417678 327922 453250 327978
rect 453306 327922 453374 327978
rect 453430 327922 453498 327978
rect 453554 327922 453622 327978
rect 453678 327922 471250 327978
rect 471306 327922 471374 327978
rect 471430 327922 471498 327978
rect 471554 327922 471622 327978
rect 471678 327922 489250 327978
rect 489306 327922 489374 327978
rect 489430 327922 489498 327978
rect 489554 327922 489622 327978
rect 489678 327922 507250 327978
rect 507306 327922 507374 327978
rect 507430 327922 507498 327978
rect 507554 327922 507622 327978
rect 507678 327922 543250 327978
rect 543306 327922 543374 327978
rect 543430 327922 543498 327978
rect 543554 327922 543622 327978
rect 543678 327922 561250 327978
rect 561306 327922 561374 327978
rect 561430 327922 561498 327978
rect 561554 327922 561622 327978
rect 561678 327922 579250 327978
rect 579306 327922 579374 327978
rect 579430 327922 579498 327978
rect 579554 327922 579622 327978
rect 579678 327922 596496 327978
rect 596552 327922 596620 327978
rect 596676 327922 596744 327978
rect 596800 327922 596868 327978
rect 596924 327922 597980 327978
rect -1916 327826 597980 327922
rect -1916 316350 597980 316446
rect -1916 316294 -1820 316350
rect -1764 316294 -1696 316350
rect -1640 316294 -1572 316350
rect -1516 316294 -1448 316350
rect -1392 316294 6970 316350
rect 7026 316294 7094 316350
rect 7150 316294 7218 316350
rect 7274 316294 7342 316350
rect 7398 316294 24970 316350
rect 25026 316294 25094 316350
rect 25150 316294 25218 316350
rect 25274 316294 25342 316350
rect 25398 316294 42970 316350
rect 43026 316294 43094 316350
rect 43150 316294 43218 316350
rect 43274 316294 43342 316350
rect 43398 316294 60970 316350
rect 61026 316294 61094 316350
rect 61150 316294 61218 316350
rect 61274 316294 61342 316350
rect 61398 316294 78970 316350
rect 79026 316294 79094 316350
rect 79150 316294 79218 316350
rect 79274 316294 79342 316350
rect 79398 316294 96970 316350
rect 97026 316294 97094 316350
rect 97150 316294 97218 316350
rect 97274 316294 97342 316350
rect 97398 316294 132970 316350
rect 133026 316294 133094 316350
rect 133150 316294 133218 316350
rect 133274 316294 133342 316350
rect 133398 316294 150970 316350
rect 151026 316294 151094 316350
rect 151150 316294 151218 316350
rect 151274 316294 151342 316350
rect 151398 316294 168970 316350
rect 169026 316294 169094 316350
rect 169150 316294 169218 316350
rect 169274 316294 169342 316350
rect 169398 316294 186970 316350
rect 187026 316294 187094 316350
rect 187150 316294 187218 316350
rect 187274 316294 187342 316350
rect 187398 316294 222970 316350
rect 223026 316294 223094 316350
rect 223150 316294 223218 316350
rect 223274 316294 223342 316350
rect 223398 316294 240970 316350
rect 241026 316294 241094 316350
rect 241150 316294 241218 316350
rect 241274 316294 241342 316350
rect 241398 316294 258970 316350
rect 259026 316294 259094 316350
rect 259150 316294 259218 316350
rect 259274 316294 259342 316350
rect 259398 316294 276970 316350
rect 277026 316294 277094 316350
rect 277150 316294 277218 316350
rect 277274 316294 277342 316350
rect 277398 316294 312970 316350
rect 313026 316294 313094 316350
rect 313150 316294 313218 316350
rect 313274 316294 313342 316350
rect 313398 316294 330970 316350
rect 331026 316294 331094 316350
rect 331150 316294 331218 316350
rect 331274 316294 331342 316350
rect 331398 316294 348970 316350
rect 349026 316294 349094 316350
rect 349150 316294 349218 316350
rect 349274 316294 349342 316350
rect 349398 316294 366970 316350
rect 367026 316294 367094 316350
rect 367150 316294 367218 316350
rect 367274 316294 367342 316350
rect 367398 316294 402970 316350
rect 403026 316294 403094 316350
rect 403150 316294 403218 316350
rect 403274 316294 403342 316350
rect 403398 316294 420970 316350
rect 421026 316294 421094 316350
rect 421150 316294 421218 316350
rect 421274 316294 421342 316350
rect 421398 316294 438970 316350
rect 439026 316294 439094 316350
rect 439150 316294 439218 316350
rect 439274 316294 439342 316350
rect 439398 316294 456970 316350
rect 457026 316294 457094 316350
rect 457150 316294 457218 316350
rect 457274 316294 457342 316350
rect 457398 316294 492970 316350
rect 493026 316294 493094 316350
rect 493150 316294 493218 316350
rect 493274 316294 493342 316350
rect 493398 316294 510970 316350
rect 511026 316294 511094 316350
rect 511150 316294 511218 316350
rect 511274 316294 511342 316350
rect 511398 316294 528970 316350
rect 529026 316294 529094 316350
rect 529150 316294 529218 316350
rect 529274 316294 529342 316350
rect 529398 316294 546970 316350
rect 547026 316294 547094 316350
rect 547150 316294 547218 316350
rect 547274 316294 547342 316350
rect 547398 316294 564970 316350
rect 565026 316294 565094 316350
rect 565150 316294 565218 316350
rect 565274 316294 565342 316350
rect 565398 316294 582970 316350
rect 583026 316294 583094 316350
rect 583150 316294 583218 316350
rect 583274 316294 583342 316350
rect 583398 316294 597456 316350
rect 597512 316294 597580 316350
rect 597636 316294 597704 316350
rect 597760 316294 597828 316350
rect 597884 316294 597980 316350
rect -1916 316226 597980 316294
rect -1916 316170 -1820 316226
rect -1764 316170 -1696 316226
rect -1640 316170 -1572 316226
rect -1516 316170 -1448 316226
rect -1392 316170 6970 316226
rect 7026 316170 7094 316226
rect 7150 316170 7218 316226
rect 7274 316170 7342 316226
rect 7398 316170 24970 316226
rect 25026 316170 25094 316226
rect 25150 316170 25218 316226
rect 25274 316170 25342 316226
rect 25398 316170 42970 316226
rect 43026 316170 43094 316226
rect 43150 316170 43218 316226
rect 43274 316170 43342 316226
rect 43398 316170 60970 316226
rect 61026 316170 61094 316226
rect 61150 316170 61218 316226
rect 61274 316170 61342 316226
rect 61398 316170 78970 316226
rect 79026 316170 79094 316226
rect 79150 316170 79218 316226
rect 79274 316170 79342 316226
rect 79398 316170 96970 316226
rect 97026 316170 97094 316226
rect 97150 316170 97218 316226
rect 97274 316170 97342 316226
rect 97398 316170 132970 316226
rect 133026 316170 133094 316226
rect 133150 316170 133218 316226
rect 133274 316170 133342 316226
rect 133398 316170 150970 316226
rect 151026 316170 151094 316226
rect 151150 316170 151218 316226
rect 151274 316170 151342 316226
rect 151398 316170 168970 316226
rect 169026 316170 169094 316226
rect 169150 316170 169218 316226
rect 169274 316170 169342 316226
rect 169398 316170 186970 316226
rect 187026 316170 187094 316226
rect 187150 316170 187218 316226
rect 187274 316170 187342 316226
rect 187398 316170 222970 316226
rect 223026 316170 223094 316226
rect 223150 316170 223218 316226
rect 223274 316170 223342 316226
rect 223398 316170 240970 316226
rect 241026 316170 241094 316226
rect 241150 316170 241218 316226
rect 241274 316170 241342 316226
rect 241398 316170 258970 316226
rect 259026 316170 259094 316226
rect 259150 316170 259218 316226
rect 259274 316170 259342 316226
rect 259398 316170 276970 316226
rect 277026 316170 277094 316226
rect 277150 316170 277218 316226
rect 277274 316170 277342 316226
rect 277398 316170 312970 316226
rect 313026 316170 313094 316226
rect 313150 316170 313218 316226
rect 313274 316170 313342 316226
rect 313398 316170 330970 316226
rect 331026 316170 331094 316226
rect 331150 316170 331218 316226
rect 331274 316170 331342 316226
rect 331398 316170 348970 316226
rect 349026 316170 349094 316226
rect 349150 316170 349218 316226
rect 349274 316170 349342 316226
rect 349398 316170 366970 316226
rect 367026 316170 367094 316226
rect 367150 316170 367218 316226
rect 367274 316170 367342 316226
rect 367398 316170 402970 316226
rect 403026 316170 403094 316226
rect 403150 316170 403218 316226
rect 403274 316170 403342 316226
rect 403398 316170 420970 316226
rect 421026 316170 421094 316226
rect 421150 316170 421218 316226
rect 421274 316170 421342 316226
rect 421398 316170 438970 316226
rect 439026 316170 439094 316226
rect 439150 316170 439218 316226
rect 439274 316170 439342 316226
rect 439398 316170 456970 316226
rect 457026 316170 457094 316226
rect 457150 316170 457218 316226
rect 457274 316170 457342 316226
rect 457398 316170 492970 316226
rect 493026 316170 493094 316226
rect 493150 316170 493218 316226
rect 493274 316170 493342 316226
rect 493398 316170 510970 316226
rect 511026 316170 511094 316226
rect 511150 316170 511218 316226
rect 511274 316170 511342 316226
rect 511398 316170 528970 316226
rect 529026 316170 529094 316226
rect 529150 316170 529218 316226
rect 529274 316170 529342 316226
rect 529398 316170 546970 316226
rect 547026 316170 547094 316226
rect 547150 316170 547218 316226
rect 547274 316170 547342 316226
rect 547398 316170 564970 316226
rect 565026 316170 565094 316226
rect 565150 316170 565218 316226
rect 565274 316170 565342 316226
rect 565398 316170 582970 316226
rect 583026 316170 583094 316226
rect 583150 316170 583218 316226
rect 583274 316170 583342 316226
rect 583398 316170 597456 316226
rect 597512 316170 597580 316226
rect 597636 316170 597704 316226
rect 597760 316170 597828 316226
rect 597884 316170 597980 316226
rect -1916 316102 597980 316170
rect -1916 316046 -1820 316102
rect -1764 316046 -1696 316102
rect -1640 316046 -1572 316102
rect -1516 316046 -1448 316102
rect -1392 316046 6970 316102
rect 7026 316046 7094 316102
rect 7150 316046 7218 316102
rect 7274 316046 7342 316102
rect 7398 316046 24970 316102
rect 25026 316046 25094 316102
rect 25150 316046 25218 316102
rect 25274 316046 25342 316102
rect 25398 316046 42970 316102
rect 43026 316046 43094 316102
rect 43150 316046 43218 316102
rect 43274 316046 43342 316102
rect 43398 316046 60970 316102
rect 61026 316046 61094 316102
rect 61150 316046 61218 316102
rect 61274 316046 61342 316102
rect 61398 316046 78970 316102
rect 79026 316046 79094 316102
rect 79150 316046 79218 316102
rect 79274 316046 79342 316102
rect 79398 316046 96970 316102
rect 97026 316046 97094 316102
rect 97150 316046 97218 316102
rect 97274 316046 97342 316102
rect 97398 316046 132970 316102
rect 133026 316046 133094 316102
rect 133150 316046 133218 316102
rect 133274 316046 133342 316102
rect 133398 316046 150970 316102
rect 151026 316046 151094 316102
rect 151150 316046 151218 316102
rect 151274 316046 151342 316102
rect 151398 316046 168970 316102
rect 169026 316046 169094 316102
rect 169150 316046 169218 316102
rect 169274 316046 169342 316102
rect 169398 316046 186970 316102
rect 187026 316046 187094 316102
rect 187150 316046 187218 316102
rect 187274 316046 187342 316102
rect 187398 316046 222970 316102
rect 223026 316046 223094 316102
rect 223150 316046 223218 316102
rect 223274 316046 223342 316102
rect 223398 316046 240970 316102
rect 241026 316046 241094 316102
rect 241150 316046 241218 316102
rect 241274 316046 241342 316102
rect 241398 316046 258970 316102
rect 259026 316046 259094 316102
rect 259150 316046 259218 316102
rect 259274 316046 259342 316102
rect 259398 316046 276970 316102
rect 277026 316046 277094 316102
rect 277150 316046 277218 316102
rect 277274 316046 277342 316102
rect 277398 316046 312970 316102
rect 313026 316046 313094 316102
rect 313150 316046 313218 316102
rect 313274 316046 313342 316102
rect 313398 316046 330970 316102
rect 331026 316046 331094 316102
rect 331150 316046 331218 316102
rect 331274 316046 331342 316102
rect 331398 316046 348970 316102
rect 349026 316046 349094 316102
rect 349150 316046 349218 316102
rect 349274 316046 349342 316102
rect 349398 316046 366970 316102
rect 367026 316046 367094 316102
rect 367150 316046 367218 316102
rect 367274 316046 367342 316102
rect 367398 316046 402970 316102
rect 403026 316046 403094 316102
rect 403150 316046 403218 316102
rect 403274 316046 403342 316102
rect 403398 316046 420970 316102
rect 421026 316046 421094 316102
rect 421150 316046 421218 316102
rect 421274 316046 421342 316102
rect 421398 316046 438970 316102
rect 439026 316046 439094 316102
rect 439150 316046 439218 316102
rect 439274 316046 439342 316102
rect 439398 316046 456970 316102
rect 457026 316046 457094 316102
rect 457150 316046 457218 316102
rect 457274 316046 457342 316102
rect 457398 316046 492970 316102
rect 493026 316046 493094 316102
rect 493150 316046 493218 316102
rect 493274 316046 493342 316102
rect 493398 316046 510970 316102
rect 511026 316046 511094 316102
rect 511150 316046 511218 316102
rect 511274 316046 511342 316102
rect 511398 316046 528970 316102
rect 529026 316046 529094 316102
rect 529150 316046 529218 316102
rect 529274 316046 529342 316102
rect 529398 316046 546970 316102
rect 547026 316046 547094 316102
rect 547150 316046 547218 316102
rect 547274 316046 547342 316102
rect 547398 316046 564970 316102
rect 565026 316046 565094 316102
rect 565150 316046 565218 316102
rect 565274 316046 565342 316102
rect 565398 316046 582970 316102
rect 583026 316046 583094 316102
rect 583150 316046 583218 316102
rect 583274 316046 583342 316102
rect 583398 316046 597456 316102
rect 597512 316046 597580 316102
rect 597636 316046 597704 316102
rect 597760 316046 597828 316102
rect 597884 316046 597980 316102
rect -1916 315978 597980 316046
rect -1916 315922 -1820 315978
rect -1764 315922 -1696 315978
rect -1640 315922 -1572 315978
rect -1516 315922 -1448 315978
rect -1392 315922 6970 315978
rect 7026 315922 7094 315978
rect 7150 315922 7218 315978
rect 7274 315922 7342 315978
rect 7398 315922 24970 315978
rect 25026 315922 25094 315978
rect 25150 315922 25218 315978
rect 25274 315922 25342 315978
rect 25398 315922 42970 315978
rect 43026 315922 43094 315978
rect 43150 315922 43218 315978
rect 43274 315922 43342 315978
rect 43398 315922 60970 315978
rect 61026 315922 61094 315978
rect 61150 315922 61218 315978
rect 61274 315922 61342 315978
rect 61398 315922 78970 315978
rect 79026 315922 79094 315978
rect 79150 315922 79218 315978
rect 79274 315922 79342 315978
rect 79398 315922 96970 315978
rect 97026 315922 97094 315978
rect 97150 315922 97218 315978
rect 97274 315922 97342 315978
rect 97398 315922 132970 315978
rect 133026 315922 133094 315978
rect 133150 315922 133218 315978
rect 133274 315922 133342 315978
rect 133398 315922 150970 315978
rect 151026 315922 151094 315978
rect 151150 315922 151218 315978
rect 151274 315922 151342 315978
rect 151398 315922 168970 315978
rect 169026 315922 169094 315978
rect 169150 315922 169218 315978
rect 169274 315922 169342 315978
rect 169398 315922 186970 315978
rect 187026 315922 187094 315978
rect 187150 315922 187218 315978
rect 187274 315922 187342 315978
rect 187398 315922 222970 315978
rect 223026 315922 223094 315978
rect 223150 315922 223218 315978
rect 223274 315922 223342 315978
rect 223398 315922 240970 315978
rect 241026 315922 241094 315978
rect 241150 315922 241218 315978
rect 241274 315922 241342 315978
rect 241398 315922 258970 315978
rect 259026 315922 259094 315978
rect 259150 315922 259218 315978
rect 259274 315922 259342 315978
rect 259398 315922 276970 315978
rect 277026 315922 277094 315978
rect 277150 315922 277218 315978
rect 277274 315922 277342 315978
rect 277398 315922 312970 315978
rect 313026 315922 313094 315978
rect 313150 315922 313218 315978
rect 313274 315922 313342 315978
rect 313398 315922 330970 315978
rect 331026 315922 331094 315978
rect 331150 315922 331218 315978
rect 331274 315922 331342 315978
rect 331398 315922 348970 315978
rect 349026 315922 349094 315978
rect 349150 315922 349218 315978
rect 349274 315922 349342 315978
rect 349398 315922 366970 315978
rect 367026 315922 367094 315978
rect 367150 315922 367218 315978
rect 367274 315922 367342 315978
rect 367398 315922 402970 315978
rect 403026 315922 403094 315978
rect 403150 315922 403218 315978
rect 403274 315922 403342 315978
rect 403398 315922 420970 315978
rect 421026 315922 421094 315978
rect 421150 315922 421218 315978
rect 421274 315922 421342 315978
rect 421398 315922 438970 315978
rect 439026 315922 439094 315978
rect 439150 315922 439218 315978
rect 439274 315922 439342 315978
rect 439398 315922 456970 315978
rect 457026 315922 457094 315978
rect 457150 315922 457218 315978
rect 457274 315922 457342 315978
rect 457398 315922 492970 315978
rect 493026 315922 493094 315978
rect 493150 315922 493218 315978
rect 493274 315922 493342 315978
rect 493398 315922 510970 315978
rect 511026 315922 511094 315978
rect 511150 315922 511218 315978
rect 511274 315922 511342 315978
rect 511398 315922 528970 315978
rect 529026 315922 529094 315978
rect 529150 315922 529218 315978
rect 529274 315922 529342 315978
rect 529398 315922 546970 315978
rect 547026 315922 547094 315978
rect 547150 315922 547218 315978
rect 547274 315922 547342 315978
rect 547398 315922 564970 315978
rect 565026 315922 565094 315978
rect 565150 315922 565218 315978
rect 565274 315922 565342 315978
rect 565398 315922 582970 315978
rect 583026 315922 583094 315978
rect 583150 315922 583218 315978
rect 583274 315922 583342 315978
rect 583398 315922 597456 315978
rect 597512 315922 597580 315978
rect 597636 315922 597704 315978
rect 597760 315922 597828 315978
rect 597884 315922 597980 315978
rect -1916 315826 597980 315922
rect -1916 310350 597980 310446
rect -1916 310294 -860 310350
rect -804 310294 -736 310350
rect -680 310294 -612 310350
rect -556 310294 -488 310350
rect -432 310294 3250 310350
rect 3306 310294 3374 310350
rect 3430 310294 3498 310350
rect 3554 310294 3622 310350
rect 3678 310294 21250 310350
rect 21306 310294 21374 310350
rect 21430 310294 21498 310350
rect 21554 310294 21622 310350
rect 21678 310294 39250 310350
rect 39306 310294 39374 310350
rect 39430 310294 39498 310350
rect 39554 310294 39622 310350
rect 39678 310294 57250 310350
rect 57306 310294 57374 310350
rect 57430 310294 57498 310350
rect 57554 310294 57622 310350
rect 57678 310294 93250 310350
rect 93306 310294 93374 310350
rect 93430 310294 93498 310350
rect 93554 310294 93622 310350
rect 93678 310294 111250 310350
rect 111306 310294 111374 310350
rect 111430 310294 111498 310350
rect 111554 310294 111622 310350
rect 111678 310294 129250 310350
rect 129306 310294 129374 310350
rect 129430 310294 129498 310350
rect 129554 310294 129622 310350
rect 129678 310294 147250 310350
rect 147306 310294 147374 310350
rect 147430 310294 147498 310350
rect 147554 310294 147622 310350
rect 147678 310294 183250 310350
rect 183306 310294 183374 310350
rect 183430 310294 183498 310350
rect 183554 310294 183622 310350
rect 183678 310294 201250 310350
rect 201306 310294 201374 310350
rect 201430 310294 201498 310350
rect 201554 310294 201622 310350
rect 201678 310294 219250 310350
rect 219306 310294 219374 310350
rect 219430 310294 219498 310350
rect 219554 310294 219622 310350
rect 219678 310294 237250 310350
rect 237306 310294 237374 310350
rect 237430 310294 237498 310350
rect 237554 310294 237622 310350
rect 237678 310294 273250 310350
rect 273306 310294 273374 310350
rect 273430 310294 273498 310350
rect 273554 310294 273622 310350
rect 273678 310294 291250 310350
rect 291306 310294 291374 310350
rect 291430 310294 291498 310350
rect 291554 310294 291622 310350
rect 291678 310294 309250 310350
rect 309306 310294 309374 310350
rect 309430 310294 309498 310350
rect 309554 310294 309622 310350
rect 309678 310294 327250 310350
rect 327306 310294 327374 310350
rect 327430 310294 327498 310350
rect 327554 310294 327622 310350
rect 327678 310294 363250 310350
rect 363306 310294 363374 310350
rect 363430 310294 363498 310350
rect 363554 310294 363622 310350
rect 363678 310294 381250 310350
rect 381306 310294 381374 310350
rect 381430 310294 381498 310350
rect 381554 310294 381622 310350
rect 381678 310294 399250 310350
rect 399306 310294 399374 310350
rect 399430 310294 399498 310350
rect 399554 310294 399622 310350
rect 399678 310294 417250 310350
rect 417306 310294 417374 310350
rect 417430 310294 417498 310350
rect 417554 310294 417622 310350
rect 417678 310294 453250 310350
rect 453306 310294 453374 310350
rect 453430 310294 453498 310350
rect 453554 310294 453622 310350
rect 453678 310294 471250 310350
rect 471306 310294 471374 310350
rect 471430 310294 471498 310350
rect 471554 310294 471622 310350
rect 471678 310294 489250 310350
rect 489306 310294 489374 310350
rect 489430 310294 489498 310350
rect 489554 310294 489622 310350
rect 489678 310294 507250 310350
rect 507306 310294 507374 310350
rect 507430 310294 507498 310350
rect 507554 310294 507622 310350
rect 507678 310294 543250 310350
rect 543306 310294 543374 310350
rect 543430 310294 543498 310350
rect 543554 310294 543622 310350
rect 543678 310294 561250 310350
rect 561306 310294 561374 310350
rect 561430 310294 561498 310350
rect 561554 310294 561622 310350
rect 561678 310294 579250 310350
rect 579306 310294 579374 310350
rect 579430 310294 579498 310350
rect 579554 310294 579622 310350
rect 579678 310294 596496 310350
rect 596552 310294 596620 310350
rect 596676 310294 596744 310350
rect 596800 310294 596868 310350
rect 596924 310294 597980 310350
rect -1916 310226 597980 310294
rect -1916 310170 -860 310226
rect -804 310170 -736 310226
rect -680 310170 -612 310226
rect -556 310170 -488 310226
rect -432 310170 3250 310226
rect 3306 310170 3374 310226
rect 3430 310170 3498 310226
rect 3554 310170 3622 310226
rect 3678 310170 21250 310226
rect 21306 310170 21374 310226
rect 21430 310170 21498 310226
rect 21554 310170 21622 310226
rect 21678 310170 39250 310226
rect 39306 310170 39374 310226
rect 39430 310170 39498 310226
rect 39554 310170 39622 310226
rect 39678 310170 57250 310226
rect 57306 310170 57374 310226
rect 57430 310170 57498 310226
rect 57554 310170 57622 310226
rect 57678 310170 93250 310226
rect 93306 310170 93374 310226
rect 93430 310170 93498 310226
rect 93554 310170 93622 310226
rect 93678 310170 111250 310226
rect 111306 310170 111374 310226
rect 111430 310170 111498 310226
rect 111554 310170 111622 310226
rect 111678 310170 129250 310226
rect 129306 310170 129374 310226
rect 129430 310170 129498 310226
rect 129554 310170 129622 310226
rect 129678 310170 147250 310226
rect 147306 310170 147374 310226
rect 147430 310170 147498 310226
rect 147554 310170 147622 310226
rect 147678 310170 183250 310226
rect 183306 310170 183374 310226
rect 183430 310170 183498 310226
rect 183554 310170 183622 310226
rect 183678 310170 201250 310226
rect 201306 310170 201374 310226
rect 201430 310170 201498 310226
rect 201554 310170 201622 310226
rect 201678 310170 219250 310226
rect 219306 310170 219374 310226
rect 219430 310170 219498 310226
rect 219554 310170 219622 310226
rect 219678 310170 237250 310226
rect 237306 310170 237374 310226
rect 237430 310170 237498 310226
rect 237554 310170 237622 310226
rect 237678 310170 273250 310226
rect 273306 310170 273374 310226
rect 273430 310170 273498 310226
rect 273554 310170 273622 310226
rect 273678 310170 291250 310226
rect 291306 310170 291374 310226
rect 291430 310170 291498 310226
rect 291554 310170 291622 310226
rect 291678 310170 309250 310226
rect 309306 310170 309374 310226
rect 309430 310170 309498 310226
rect 309554 310170 309622 310226
rect 309678 310170 327250 310226
rect 327306 310170 327374 310226
rect 327430 310170 327498 310226
rect 327554 310170 327622 310226
rect 327678 310170 363250 310226
rect 363306 310170 363374 310226
rect 363430 310170 363498 310226
rect 363554 310170 363622 310226
rect 363678 310170 381250 310226
rect 381306 310170 381374 310226
rect 381430 310170 381498 310226
rect 381554 310170 381622 310226
rect 381678 310170 399250 310226
rect 399306 310170 399374 310226
rect 399430 310170 399498 310226
rect 399554 310170 399622 310226
rect 399678 310170 417250 310226
rect 417306 310170 417374 310226
rect 417430 310170 417498 310226
rect 417554 310170 417622 310226
rect 417678 310170 453250 310226
rect 453306 310170 453374 310226
rect 453430 310170 453498 310226
rect 453554 310170 453622 310226
rect 453678 310170 471250 310226
rect 471306 310170 471374 310226
rect 471430 310170 471498 310226
rect 471554 310170 471622 310226
rect 471678 310170 489250 310226
rect 489306 310170 489374 310226
rect 489430 310170 489498 310226
rect 489554 310170 489622 310226
rect 489678 310170 507250 310226
rect 507306 310170 507374 310226
rect 507430 310170 507498 310226
rect 507554 310170 507622 310226
rect 507678 310170 543250 310226
rect 543306 310170 543374 310226
rect 543430 310170 543498 310226
rect 543554 310170 543622 310226
rect 543678 310170 561250 310226
rect 561306 310170 561374 310226
rect 561430 310170 561498 310226
rect 561554 310170 561622 310226
rect 561678 310170 579250 310226
rect 579306 310170 579374 310226
rect 579430 310170 579498 310226
rect 579554 310170 579622 310226
rect 579678 310170 596496 310226
rect 596552 310170 596620 310226
rect 596676 310170 596744 310226
rect 596800 310170 596868 310226
rect 596924 310170 597980 310226
rect -1916 310102 597980 310170
rect -1916 310046 -860 310102
rect -804 310046 -736 310102
rect -680 310046 -612 310102
rect -556 310046 -488 310102
rect -432 310046 3250 310102
rect 3306 310046 3374 310102
rect 3430 310046 3498 310102
rect 3554 310046 3622 310102
rect 3678 310046 21250 310102
rect 21306 310046 21374 310102
rect 21430 310046 21498 310102
rect 21554 310046 21622 310102
rect 21678 310046 39250 310102
rect 39306 310046 39374 310102
rect 39430 310046 39498 310102
rect 39554 310046 39622 310102
rect 39678 310046 57250 310102
rect 57306 310046 57374 310102
rect 57430 310046 57498 310102
rect 57554 310046 57622 310102
rect 57678 310046 93250 310102
rect 93306 310046 93374 310102
rect 93430 310046 93498 310102
rect 93554 310046 93622 310102
rect 93678 310046 111250 310102
rect 111306 310046 111374 310102
rect 111430 310046 111498 310102
rect 111554 310046 111622 310102
rect 111678 310046 129250 310102
rect 129306 310046 129374 310102
rect 129430 310046 129498 310102
rect 129554 310046 129622 310102
rect 129678 310046 147250 310102
rect 147306 310046 147374 310102
rect 147430 310046 147498 310102
rect 147554 310046 147622 310102
rect 147678 310046 183250 310102
rect 183306 310046 183374 310102
rect 183430 310046 183498 310102
rect 183554 310046 183622 310102
rect 183678 310046 201250 310102
rect 201306 310046 201374 310102
rect 201430 310046 201498 310102
rect 201554 310046 201622 310102
rect 201678 310046 219250 310102
rect 219306 310046 219374 310102
rect 219430 310046 219498 310102
rect 219554 310046 219622 310102
rect 219678 310046 237250 310102
rect 237306 310046 237374 310102
rect 237430 310046 237498 310102
rect 237554 310046 237622 310102
rect 237678 310046 273250 310102
rect 273306 310046 273374 310102
rect 273430 310046 273498 310102
rect 273554 310046 273622 310102
rect 273678 310046 291250 310102
rect 291306 310046 291374 310102
rect 291430 310046 291498 310102
rect 291554 310046 291622 310102
rect 291678 310046 309250 310102
rect 309306 310046 309374 310102
rect 309430 310046 309498 310102
rect 309554 310046 309622 310102
rect 309678 310046 327250 310102
rect 327306 310046 327374 310102
rect 327430 310046 327498 310102
rect 327554 310046 327622 310102
rect 327678 310046 363250 310102
rect 363306 310046 363374 310102
rect 363430 310046 363498 310102
rect 363554 310046 363622 310102
rect 363678 310046 381250 310102
rect 381306 310046 381374 310102
rect 381430 310046 381498 310102
rect 381554 310046 381622 310102
rect 381678 310046 399250 310102
rect 399306 310046 399374 310102
rect 399430 310046 399498 310102
rect 399554 310046 399622 310102
rect 399678 310046 417250 310102
rect 417306 310046 417374 310102
rect 417430 310046 417498 310102
rect 417554 310046 417622 310102
rect 417678 310046 453250 310102
rect 453306 310046 453374 310102
rect 453430 310046 453498 310102
rect 453554 310046 453622 310102
rect 453678 310046 471250 310102
rect 471306 310046 471374 310102
rect 471430 310046 471498 310102
rect 471554 310046 471622 310102
rect 471678 310046 489250 310102
rect 489306 310046 489374 310102
rect 489430 310046 489498 310102
rect 489554 310046 489622 310102
rect 489678 310046 507250 310102
rect 507306 310046 507374 310102
rect 507430 310046 507498 310102
rect 507554 310046 507622 310102
rect 507678 310046 543250 310102
rect 543306 310046 543374 310102
rect 543430 310046 543498 310102
rect 543554 310046 543622 310102
rect 543678 310046 561250 310102
rect 561306 310046 561374 310102
rect 561430 310046 561498 310102
rect 561554 310046 561622 310102
rect 561678 310046 579250 310102
rect 579306 310046 579374 310102
rect 579430 310046 579498 310102
rect 579554 310046 579622 310102
rect 579678 310046 596496 310102
rect 596552 310046 596620 310102
rect 596676 310046 596744 310102
rect 596800 310046 596868 310102
rect 596924 310046 597980 310102
rect -1916 309978 597980 310046
rect -1916 309922 -860 309978
rect -804 309922 -736 309978
rect -680 309922 -612 309978
rect -556 309922 -488 309978
rect -432 309922 3250 309978
rect 3306 309922 3374 309978
rect 3430 309922 3498 309978
rect 3554 309922 3622 309978
rect 3678 309922 21250 309978
rect 21306 309922 21374 309978
rect 21430 309922 21498 309978
rect 21554 309922 21622 309978
rect 21678 309922 39250 309978
rect 39306 309922 39374 309978
rect 39430 309922 39498 309978
rect 39554 309922 39622 309978
rect 39678 309922 57250 309978
rect 57306 309922 57374 309978
rect 57430 309922 57498 309978
rect 57554 309922 57622 309978
rect 57678 309922 93250 309978
rect 93306 309922 93374 309978
rect 93430 309922 93498 309978
rect 93554 309922 93622 309978
rect 93678 309922 111250 309978
rect 111306 309922 111374 309978
rect 111430 309922 111498 309978
rect 111554 309922 111622 309978
rect 111678 309922 129250 309978
rect 129306 309922 129374 309978
rect 129430 309922 129498 309978
rect 129554 309922 129622 309978
rect 129678 309922 147250 309978
rect 147306 309922 147374 309978
rect 147430 309922 147498 309978
rect 147554 309922 147622 309978
rect 147678 309922 183250 309978
rect 183306 309922 183374 309978
rect 183430 309922 183498 309978
rect 183554 309922 183622 309978
rect 183678 309922 201250 309978
rect 201306 309922 201374 309978
rect 201430 309922 201498 309978
rect 201554 309922 201622 309978
rect 201678 309922 219250 309978
rect 219306 309922 219374 309978
rect 219430 309922 219498 309978
rect 219554 309922 219622 309978
rect 219678 309922 237250 309978
rect 237306 309922 237374 309978
rect 237430 309922 237498 309978
rect 237554 309922 237622 309978
rect 237678 309922 273250 309978
rect 273306 309922 273374 309978
rect 273430 309922 273498 309978
rect 273554 309922 273622 309978
rect 273678 309922 291250 309978
rect 291306 309922 291374 309978
rect 291430 309922 291498 309978
rect 291554 309922 291622 309978
rect 291678 309922 309250 309978
rect 309306 309922 309374 309978
rect 309430 309922 309498 309978
rect 309554 309922 309622 309978
rect 309678 309922 327250 309978
rect 327306 309922 327374 309978
rect 327430 309922 327498 309978
rect 327554 309922 327622 309978
rect 327678 309922 363250 309978
rect 363306 309922 363374 309978
rect 363430 309922 363498 309978
rect 363554 309922 363622 309978
rect 363678 309922 381250 309978
rect 381306 309922 381374 309978
rect 381430 309922 381498 309978
rect 381554 309922 381622 309978
rect 381678 309922 399250 309978
rect 399306 309922 399374 309978
rect 399430 309922 399498 309978
rect 399554 309922 399622 309978
rect 399678 309922 417250 309978
rect 417306 309922 417374 309978
rect 417430 309922 417498 309978
rect 417554 309922 417622 309978
rect 417678 309922 453250 309978
rect 453306 309922 453374 309978
rect 453430 309922 453498 309978
rect 453554 309922 453622 309978
rect 453678 309922 471250 309978
rect 471306 309922 471374 309978
rect 471430 309922 471498 309978
rect 471554 309922 471622 309978
rect 471678 309922 489250 309978
rect 489306 309922 489374 309978
rect 489430 309922 489498 309978
rect 489554 309922 489622 309978
rect 489678 309922 507250 309978
rect 507306 309922 507374 309978
rect 507430 309922 507498 309978
rect 507554 309922 507622 309978
rect 507678 309922 543250 309978
rect 543306 309922 543374 309978
rect 543430 309922 543498 309978
rect 543554 309922 543622 309978
rect 543678 309922 561250 309978
rect 561306 309922 561374 309978
rect 561430 309922 561498 309978
rect 561554 309922 561622 309978
rect 561678 309922 579250 309978
rect 579306 309922 579374 309978
rect 579430 309922 579498 309978
rect 579554 309922 579622 309978
rect 579678 309922 596496 309978
rect 596552 309922 596620 309978
rect 596676 309922 596744 309978
rect 596800 309922 596868 309978
rect 596924 309922 597980 309978
rect -1916 309826 597980 309922
rect -1916 298350 597980 298446
rect -1916 298294 -1820 298350
rect -1764 298294 -1696 298350
rect -1640 298294 -1572 298350
rect -1516 298294 -1448 298350
rect -1392 298294 6970 298350
rect 7026 298294 7094 298350
rect 7150 298294 7218 298350
rect 7274 298294 7342 298350
rect 7398 298294 24970 298350
rect 25026 298294 25094 298350
rect 25150 298294 25218 298350
rect 25274 298294 25342 298350
rect 25398 298294 42970 298350
rect 43026 298294 43094 298350
rect 43150 298294 43218 298350
rect 43274 298294 43342 298350
rect 43398 298294 60970 298350
rect 61026 298294 61094 298350
rect 61150 298294 61218 298350
rect 61274 298294 61342 298350
rect 61398 298294 78970 298350
rect 79026 298294 79094 298350
rect 79150 298294 79218 298350
rect 79274 298294 79342 298350
rect 79398 298294 96970 298350
rect 97026 298294 97094 298350
rect 97150 298294 97218 298350
rect 97274 298294 97342 298350
rect 97398 298294 132970 298350
rect 133026 298294 133094 298350
rect 133150 298294 133218 298350
rect 133274 298294 133342 298350
rect 133398 298294 150970 298350
rect 151026 298294 151094 298350
rect 151150 298294 151218 298350
rect 151274 298294 151342 298350
rect 151398 298294 168970 298350
rect 169026 298294 169094 298350
rect 169150 298294 169218 298350
rect 169274 298294 169342 298350
rect 169398 298294 186970 298350
rect 187026 298294 187094 298350
rect 187150 298294 187218 298350
rect 187274 298294 187342 298350
rect 187398 298294 222970 298350
rect 223026 298294 223094 298350
rect 223150 298294 223218 298350
rect 223274 298294 223342 298350
rect 223398 298294 240970 298350
rect 241026 298294 241094 298350
rect 241150 298294 241218 298350
rect 241274 298294 241342 298350
rect 241398 298294 258970 298350
rect 259026 298294 259094 298350
rect 259150 298294 259218 298350
rect 259274 298294 259342 298350
rect 259398 298294 276970 298350
rect 277026 298294 277094 298350
rect 277150 298294 277218 298350
rect 277274 298294 277342 298350
rect 277398 298294 312970 298350
rect 313026 298294 313094 298350
rect 313150 298294 313218 298350
rect 313274 298294 313342 298350
rect 313398 298294 330970 298350
rect 331026 298294 331094 298350
rect 331150 298294 331218 298350
rect 331274 298294 331342 298350
rect 331398 298294 348970 298350
rect 349026 298294 349094 298350
rect 349150 298294 349218 298350
rect 349274 298294 349342 298350
rect 349398 298294 366970 298350
rect 367026 298294 367094 298350
rect 367150 298294 367218 298350
rect 367274 298294 367342 298350
rect 367398 298294 402970 298350
rect 403026 298294 403094 298350
rect 403150 298294 403218 298350
rect 403274 298294 403342 298350
rect 403398 298294 420970 298350
rect 421026 298294 421094 298350
rect 421150 298294 421218 298350
rect 421274 298294 421342 298350
rect 421398 298294 438970 298350
rect 439026 298294 439094 298350
rect 439150 298294 439218 298350
rect 439274 298294 439342 298350
rect 439398 298294 456970 298350
rect 457026 298294 457094 298350
rect 457150 298294 457218 298350
rect 457274 298294 457342 298350
rect 457398 298294 492970 298350
rect 493026 298294 493094 298350
rect 493150 298294 493218 298350
rect 493274 298294 493342 298350
rect 493398 298294 510970 298350
rect 511026 298294 511094 298350
rect 511150 298294 511218 298350
rect 511274 298294 511342 298350
rect 511398 298294 528970 298350
rect 529026 298294 529094 298350
rect 529150 298294 529218 298350
rect 529274 298294 529342 298350
rect 529398 298294 546970 298350
rect 547026 298294 547094 298350
rect 547150 298294 547218 298350
rect 547274 298294 547342 298350
rect 547398 298294 564970 298350
rect 565026 298294 565094 298350
rect 565150 298294 565218 298350
rect 565274 298294 565342 298350
rect 565398 298294 582970 298350
rect 583026 298294 583094 298350
rect 583150 298294 583218 298350
rect 583274 298294 583342 298350
rect 583398 298294 597456 298350
rect 597512 298294 597580 298350
rect 597636 298294 597704 298350
rect 597760 298294 597828 298350
rect 597884 298294 597980 298350
rect -1916 298226 597980 298294
rect -1916 298170 -1820 298226
rect -1764 298170 -1696 298226
rect -1640 298170 -1572 298226
rect -1516 298170 -1448 298226
rect -1392 298170 6970 298226
rect 7026 298170 7094 298226
rect 7150 298170 7218 298226
rect 7274 298170 7342 298226
rect 7398 298170 24970 298226
rect 25026 298170 25094 298226
rect 25150 298170 25218 298226
rect 25274 298170 25342 298226
rect 25398 298170 42970 298226
rect 43026 298170 43094 298226
rect 43150 298170 43218 298226
rect 43274 298170 43342 298226
rect 43398 298170 60970 298226
rect 61026 298170 61094 298226
rect 61150 298170 61218 298226
rect 61274 298170 61342 298226
rect 61398 298170 78970 298226
rect 79026 298170 79094 298226
rect 79150 298170 79218 298226
rect 79274 298170 79342 298226
rect 79398 298170 96970 298226
rect 97026 298170 97094 298226
rect 97150 298170 97218 298226
rect 97274 298170 97342 298226
rect 97398 298170 132970 298226
rect 133026 298170 133094 298226
rect 133150 298170 133218 298226
rect 133274 298170 133342 298226
rect 133398 298170 150970 298226
rect 151026 298170 151094 298226
rect 151150 298170 151218 298226
rect 151274 298170 151342 298226
rect 151398 298170 168970 298226
rect 169026 298170 169094 298226
rect 169150 298170 169218 298226
rect 169274 298170 169342 298226
rect 169398 298170 186970 298226
rect 187026 298170 187094 298226
rect 187150 298170 187218 298226
rect 187274 298170 187342 298226
rect 187398 298170 222970 298226
rect 223026 298170 223094 298226
rect 223150 298170 223218 298226
rect 223274 298170 223342 298226
rect 223398 298170 240970 298226
rect 241026 298170 241094 298226
rect 241150 298170 241218 298226
rect 241274 298170 241342 298226
rect 241398 298170 258970 298226
rect 259026 298170 259094 298226
rect 259150 298170 259218 298226
rect 259274 298170 259342 298226
rect 259398 298170 276970 298226
rect 277026 298170 277094 298226
rect 277150 298170 277218 298226
rect 277274 298170 277342 298226
rect 277398 298170 312970 298226
rect 313026 298170 313094 298226
rect 313150 298170 313218 298226
rect 313274 298170 313342 298226
rect 313398 298170 330970 298226
rect 331026 298170 331094 298226
rect 331150 298170 331218 298226
rect 331274 298170 331342 298226
rect 331398 298170 348970 298226
rect 349026 298170 349094 298226
rect 349150 298170 349218 298226
rect 349274 298170 349342 298226
rect 349398 298170 366970 298226
rect 367026 298170 367094 298226
rect 367150 298170 367218 298226
rect 367274 298170 367342 298226
rect 367398 298170 402970 298226
rect 403026 298170 403094 298226
rect 403150 298170 403218 298226
rect 403274 298170 403342 298226
rect 403398 298170 420970 298226
rect 421026 298170 421094 298226
rect 421150 298170 421218 298226
rect 421274 298170 421342 298226
rect 421398 298170 438970 298226
rect 439026 298170 439094 298226
rect 439150 298170 439218 298226
rect 439274 298170 439342 298226
rect 439398 298170 456970 298226
rect 457026 298170 457094 298226
rect 457150 298170 457218 298226
rect 457274 298170 457342 298226
rect 457398 298170 492970 298226
rect 493026 298170 493094 298226
rect 493150 298170 493218 298226
rect 493274 298170 493342 298226
rect 493398 298170 510970 298226
rect 511026 298170 511094 298226
rect 511150 298170 511218 298226
rect 511274 298170 511342 298226
rect 511398 298170 528970 298226
rect 529026 298170 529094 298226
rect 529150 298170 529218 298226
rect 529274 298170 529342 298226
rect 529398 298170 546970 298226
rect 547026 298170 547094 298226
rect 547150 298170 547218 298226
rect 547274 298170 547342 298226
rect 547398 298170 564970 298226
rect 565026 298170 565094 298226
rect 565150 298170 565218 298226
rect 565274 298170 565342 298226
rect 565398 298170 582970 298226
rect 583026 298170 583094 298226
rect 583150 298170 583218 298226
rect 583274 298170 583342 298226
rect 583398 298170 597456 298226
rect 597512 298170 597580 298226
rect 597636 298170 597704 298226
rect 597760 298170 597828 298226
rect 597884 298170 597980 298226
rect -1916 298102 597980 298170
rect -1916 298046 -1820 298102
rect -1764 298046 -1696 298102
rect -1640 298046 -1572 298102
rect -1516 298046 -1448 298102
rect -1392 298046 6970 298102
rect 7026 298046 7094 298102
rect 7150 298046 7218 298102
rect 7274 298046 7342 298102
rect 7398 298046 24970 298102
rect 25026 298046 25094 298102
rect 25150 298046 25218 298102
rect 25274 298046 25342 298102
rect 25398 298046 42970 298102
rect 43026 298046 43094 298102
rect 43150 298046 43218 298102
rect 43274 298046 43342 298102
rect 43398 298046 60970 298102
rect 61026 298046 61094 298102
rect 61150 298046 61218 298102
rect 61274 298046 61342 298102
rect 61398 298046 78970 298102
rect 79026 298046 79094 298102
rect 79150 298046 79218 298102
rect 79274 298046 79342 298102
rect 79398 298046 96970 298102
rect 97026 298046 97094 298102
rect 97150 298046 97218 298102
rect 97274 298046 97342 298102
rect 97398 298046 132970 298102
rect 133026 298046 133094 298102
rect 133150 298046 133218 298102
rect 133274 298046 133342 298102
rect 133398 298046 150970 298102
rect 151026 298046 151094 298102
rect 151150 298046 151218 298102
rect 151274 298046 151342 298102
rect 151398 298046 168970 298102
rect 169026 298046 169094 298102
rect 169150 298046 169218 298102
rect 169274 298046 169342 298102
rect 169398 298046 186970 298102
rect 187026 298046 187094 298102
rect 187150 298046 187218 298102
rect 187274 298046 187342 298102
rect 187398 298046 222970 298102
rect 223026 298046 223094 298102
rect 223150 298046 223218 298102
rect 223274 298046 223342 298102
rect 223398 298046 240970 298102
rect 241026 298046 241094 298102
rect 241150 298046 241218 298102
rect 241274 298046 241342 298102
rect 241398 298046 258970 298102
rect 259026 298046 259094 298102
rect 259150 298046 259218 298102
rect 259274 298046 259342 298102
rect 259398 298046 276970 298102
rect 277026 298046 277094 298102
rect 277150 298046 277218 298102
rect 277274 298046 277342 298102
rect 277398 298046 312970 298102
rect 313026 298046 313094 298102
rect 313150 298046 313218 298102
rect 313274 298046 313342 298102
rect 313398 298046 330970 298102
rect 331026 298046 331094 298102
rect 331150 298046 331218 298102
rect 331274 298046 331342 298102
rect 331398 298046 348970 298102
rect 349026 298046 349094 298102
rect 349150 298046 349218 298102
rect 349274 298046 349342 298102
rect 349398 298046 366970 298102
rect 367026 298046 367094 298102
rect 367150 298046 367218 298102
rect 367274 298046 367342 298102
rect 367398 298046 402970 298102
rect 403026 298046 403094 298102
rect 403150 298046 403218 298102
rect 403274 298046 403342 298102
rect 403398 298046 420970 298102
rect 421026 298046 421094 298102
rect 421150 298046 421218 298102
rect 421274 298046 421342 298102
rect 421398 298046 438970 298102
rect 439026 298046 439094 298102
rect 439150 298046 439218 298102
rect 439274 298046 439342 298102
rect 439398 298046 456970 298102
rect 457026 298046 457094 298102
rect 457150 298046 457218 298102
rect 457274 298046 457342 298102
rect 457398 298046 492970 298102
rect 493026 298046 493094 298102
rect 493150 298046 493218 298102
rect 493274 298046 493342 298102
rect 493398 298046 510970 298102
rect 511026 298046 511094 298102
rect 511150 298046 511218 298102
rect 511274 298046 511342 298102
rect 511398 298046 528970 298102
rect 529026 298046 529094 298102
rect 529150 298046 529218 298102
rect 529274 298046 529342 298102
rect 529398 298046 546970 298102
rect 547026 298046 547094 298102
rect 547150 298046 547218 298102
rect 547274 298046 547342 298102
rect 547398 298046 564970 298102
rect 565026 298046 565094 298102
rect 565150 298046 565218 298102
rect 565274 298046 565342 298102
rect 565398 298046 582970 298102
rect 583026 298046 583094 298102
rect 583150 298046 583218 298102
rect 583274 298046 583342 298102
rect 583398 298046 597456 298102
rect 597512 298046 597580 298102
rect 597636 298046 597704 298102
rect 597760 298046 597828 298102
rect 597884 298046 597980 298102
rect -1916 297978 597980 298046
rect -1916 297922 -1820 297978
rect -1764 297922 -1696 297978
rect -1640 297922 -1572 297978
rect -1516 297922 -1448 297978
rect -1392 297922 6970 297978
rect 7026 297922 7094 297978
rect 7150 297922 7218 297978
rect 7274 297922 7342 297978
rect 7398 297922 24970 297978
rect 25026 297922 25094 297978
rect 25150 297922 25218 297978
rect 25274 297922 25342 297978
rect 25398 297922 42970 297978
rect 43026 297922 43094 297978
rect 43150 297922 43218 297978
rect 43274 297922 43342 297978
rect 43398 297922 60970 297978
rect 61026 297922 61094 297978
rect 61150 297922 61218 297978
rect 61274 297922 61342 297978
rect 61398 297922 78970 297978
rect 79026 297922 79094 297978
rect 79150 297922 79218 297978
rect 79274 297922 79342 297978
rect 79398 297922 96970 297978
rect 97026 297922 97094 297978
rect 97150 297922 97218 297978
rect 97274 297922 97342 297978
rect 97398 297922 132970 297978
rect 133026 297922 133094 297978
rect 133150 297922 133218 297978
rect 133274 297922 133342 297978
rect 133398 297922 150970 297978
rect 151026 297922 151094 297978
rect 151150 297922 151218 297978
rect 151274 297922 151342 297978
rect 151398 297922 168970 297978
rect 169026 297922 169094 297978
rect 169150 297922 169218 297978
rect 169274 297922 169342 297978
rect 169398 297922 186970 297978
rect 187026 297922 187094 297978
rect 187150 297922 187218 297978
rect 187274 297922 187342 297978
rect 187398 297922 222970 297978
rect 223026 297922 223094 297978
rect 223150 297922 223218 297978
rect 223274 297922 223342 297978
rect 223398 297922 240970 297978
rect 241026 297922 241094 297978
rect 241150 297922 241218 297978
rect 241274 297922 241342 297978
rect 241398 297922 258970 297978
rect 259026 297922 259094 297978
rect 259150 297922 259218 297978
rect 259274 297922 259342 297978
rect 259398 297922 276970 297978
rect 277026 297922 277094 297978
rect 277150 297922 277218 297978
rect 277274 297922 277342 297978
rect 277398 297922 312970 297978
rect 313026 297922 313094 297978
rect 313150 297922 313218 297978
rect 313274 297922 313342 297978
rect 313398 297922 330970 297978
rect 331026 297922 331094 297978
rect 331150 297922 331218 297978
rect 331274 297922 331342 297978
rect 331398 297922 348970 297978
rect 349026 297922 349094 297978
rect 349150 297922 349218 297978
rect 349274 297922 349342 297978
rect 349398 297922 366970 297978
rect 367026 297922 367094 297978
rect 367150 297922 367218 297978
rect 367274 297922 367342 297978
rect 367398 297922 402970 297978
rect 403026 297922 403094 297978
rect 403150 297922 403218 297978
rect 403274 297922 403342 297978
rect 403398 297922 420970 297978
rect 421026 297922 421094 297978
rect 421150 297922 421218 297978
rect 421274 297922 421342 297978
rect 421398 297922 438970 297978
rect 439026 297922 439094 297978
rect 439150 297922 439218 297978
rect 439274 297922 439342 297978
rect 439398 297922 456970 297978
rect 457026 297922 457094 297978
rect 457150 297922 457218 297978
rect 457274 297922 457342 297978
rect 457398 297922 492970 297978
rect 493026 297922 493094 297978
rect 493150 297922 493218 297978
rect 493274 297922 493342 297978
rect 493398 297922 510970 297978
rect 511026 297922 511094 297978
rect 511150 297922 511218 297978
rect 511274 297922 511342 297978
rect 511398 297922 528970 297978
rect 529026 297922 529094 297978
rect 529150 297922 529218 297978
rect 529274 297922 529342 297978
rect 529398 297922 546970 297978
rect 547026 297922 547094 297978
rect 547150 297922 547218 297978
rect 547274 297922 547342 297978
rect 547398 297922 564970 297978
rect 565026 297922 565094 297978
rect 565150 297922 565218 297978
rect 565274 297922 565342 297978
rect 565398 297922 582970 297978
rect 583026 297922 583094 297978
rect 583150 297922 583218 297978
rect 583274 297922 583342 297978
rect 583398 297922 597456 297978
rect 597512 297922 597580 297978
rect 597636 297922 597704 297978
rect 597760 297922 597828 297978
rect 597884 297922 597980 297978
rect -1916 297826 597980 297922
rect -1916 292350 597980 292446
rect -1916 292294 -860 292350
rect -804 292294 -736 292350
rect -680 292294 -612 292350
rect -556 292294 -488 292350
rect -432 292294 3250 292350
rect 3306 292294 3374 292350
rect 3430 292294 3498 292350
rect 3554 292294 3622 292350
rect 3678 292294 21250 292350
rect 21306 292294 21374 292350
rect 21430 292294 21498 292350
rect 21554 292294 21622 292350
rect 21678 292294 39250 292350
rect 39306 292294 39374 292350
rect 39430 292294 39498 292350
rect 39554 292294 39622 292350
rect 39678 292294 57250 292350
rect 57306 292294 57374 292350
rect 57430 292294 57498 292350
rect 57554 292294 57622 292350
rect 57678 292294 93250 292350
rect 93306 292294 93374 292350
rect 93430 292294 93498 292350
rect 93554 292294 93622 292350
rect 93678 292294 111250 292350
rect 111306 292294 111374 292350
rect 111430 292294 111498 292350
rect 111554 292294 111622 292350
rect 111678 292294 129250 292350
rect 129306 292294 129374 292350
rect 129430 292294 129498 292350
rect 129554 292294 129622 292350
rect 129678 292294 147250 292350
rect 147306 292294 147374 292350
rect 147430 292294 147498 292350
rect 147554 292294 147622 292350
rect 147678 292294 183250 292350
rect 183306 292294 183374 292350
rect 183430 292294 183498 292350
rect 183554 292294 183622 292350
rect 183678 292294 201250 292350
rect 201306 292294 201374 292350
rect 201430 292294 201498 292350
rect 201554 292294 201622 292350
rect 201678 292294 219250 292350
rect 219306 292294 219374 292350
rect 219430 292294 219498 292350
rect 219554 292294 219622 292350
rect 219678 292294 237250 292350
rect 237306 292294 237374 292350
rect 237430 292294 237498 292350
rect 237554 292294 237622 292350
rect 237678 292294 273250 292350
rect 273306 292294 273374 292350
rect 273430 292294 273498 292350
rect 273554 292294 273622 292350
rect 273678 292294 291250 292350
rect 291306 292294 291374 292350
rect 291430 292294 291498 292350
rect 291554 292294 291622 292350
rect 291678 292294 309250 292350
rect 309306 292294 309374 292350
rect 309430 292294 309498 292350
rect 309554 292294 309622 292350
rect 309678 292294 327250 292350
rect 327306 292294 327374 292350
rect 327430 292294 327498 292350
rect 327554 292294 327622 292350
rect 327678 292294 363250 292350
rect 363306 292294 363374 292350
rect 363430 292294 363498 292350
rect 363554 292294 363622 292350
rect 363678 292294 381250 292350
rect 381306 292294 381374 292350
rect 381430 292294 381498 292350
rect 381554 292294 381622 292350
rect 381678 292294 399250 292350
rect 399306 292294 399374 292350
rect 399430 292294 399498 292350
rect 399554 292294 399622 292350
rect 399678 292294 417250 292350
rect 417306 292294 417374 292350
rect 417430 292294 417498 292350
rect 417554 292294 417622 292350
rect 417678 292294 453250 292350
rect 453306 292294 453374 292350
rect 453430 292294 453498 292350
rect 453554 292294 453622 292350
rect 453678 292294 471250 292350
rect 471306 292294 471374 292350
rect 471430 292294 471498 292350
rect 471554 292294 471622 292350
rect 471678 292294 489250 292350
rect 489306 292294 489374 292350
rect 489430 292294 489498 292350
rect 489554 292294 489622 292350
rect 489678 292294 507250 292350
rect 507306 292294 507374 292350
rect 507430 292294 507498 292350
rect 507554 292294 507622 292350
rect 507678 292294 543250 292350
rect 543306 292294 543374 292350
rect 543430 292294 543498 292350
rect 543554 292294 543622 292350
rect 543678 292294 561250 292350
rect 561306 292294 561374 292350
rect 561430 292294 561498 292350
rect 561554 292294 561622 292350
rect 561678 292294 579250 292350
rect 579306 292294 579374 292350
rect 579430 292294 579498 292350
rect 579554 292294 579622 292350
rect 579678 292294 596496 292350
rect 596552 292294 596620 292350
rect 596676 292294 596744 292350
rect 596800 292294 596868 292350
rect 596924 292294 597980 292350
rect -1916 292226 597980 292294
rect -1916 292170 -860 292226
rect -804 292170 -736 292226
rect -680 292170 -612 292226
rect -556 292170 -488 292226
rect -432 292170 3250 292226
rect 3306 292170 3374 292226
rect 3430 292170 3498 292226
rect 3554 292170 3622 292226
rect 3678 292170 21250 292226
rect 21306 292170 21374 292226
rect 21430 292170 21498 292226
rect 21554 292170 21622 292226
rect 21678 292170 39250 292226
rect 39306 292170 39374 292226
rect 39430 292170 39498 292226
rect 39554 292170 39622 292226
rect 39678 292170 57250 292226
rect 57306 292170 57374 292226
rect 57430 292170 57498 292226
rect 57554 292170 57622 292226
rect 57678 292170 93250 292226
rect 93306 292170 93374 292226
rect 93430 292170 93498 292226
rect 93554 292170 93622 292226
rect 93678 292170 111250 292226
rect 111306 292170 111374 292226
rect 111430 292170 111498 292226
rect 111554 292170 111622 292226
rect 111678 292170 129250 292226
rect 129306 292170 129374 292226
rect 129430 292170 129498 292226
rect 129554 292170 129622 292226
rect 129678 292170 147250 292226
rect 147306 292170 147374 292226
rect 147430 292170 147498 292226
rect 147554 292170 147622 292226
rect 147678 292170 183250 292226
rect 183306 292170 183374 292226
rect 183430 292170 183498 292226
rect 183554 292170 183622 292226
rect 183678 292170 201250 292226
rect 201306 292170 201374 292226
rect 201430 292170 201498 292226
rect 201554 292170 201622 292226
rect 201678 292170 219250 292226
rect 219306 292170 219374 292226
rect 219430 292170 219498 292226
rect 219554 292170 219622 292226
rect 219678 292170 237250 292226
rect 237306 292170 237374 292226
rect 237430 292170 237498 292226
rect 237554 292170 237622 292226
rect 237678 292170 273250 292226
rect 273306 292170 273374 292226
rect 273430 292170 273498 292226
rect 273554 292170 273622 292226
rect 273678 292170 291250 292226
rect 291306 292170 291374 292226
rect 291430 292170 291498 292226
rect 291554 292170 291622 292226
rect 291678 292170 309250 292226
rect 309306 292170 309374 292226
rect 309430 292170 309498 292226
rect 309554 292170 309622 292226
rect 309678 292170 327250 292226
rect 327306 292170 327374 292226
rect 327430 292170 327498 292226
rect 327554 292170 327622 292226
rect 327678 292170 363250 292226
rect 363306 292170 363374 292226
rect 363430 292170 363498 292226
rect 363554 292170 363622 292226
rect 363678 292170 381250 292226
rect 381306 292170 381374 292226
rect 381430 292170 381498 292226
rect 381554 292170 381622 292226
rect 381678 292170 399250 292226
rect 399306 292170 399374 292226
rect 399430 292170 399498 292226
rect 399554 292170 399622 292226
rect 399678 292170 417250 292226
rect 417306 292170 417374 292226
rect 417430 292170 417498 292226
rect 417554 292170 417622 292226
rect 417678 292170 453250 292226
rect 453306 292170 453374 292226
rect 453430 292170 453498 292226
rect 453554 292170 453622 292226
rect 453678 292170 471250 292226
rect 471306 292170 471374 292226
rect 471430 292170 471498 292226
rect 471554 292170 471622 292226
rect 471678 292170 489250 292226
rect 489306 292170 489374 292226
rect 489430 292170 489498 292226
rect 489554 292170 489622 292226
rect 489678 292170 507250 292226
rect 507306 292170 507374 292226
rect 507430 292170 507498 292226
rect 507554 292170 507622 292226
rect 507678 292170 543250 292226
rect 543306 292170 543374 292226
rect 543430 292170 543498 292226
rect 543554 292170 543622 292226
rect 543678 292170 561250 292226
rect 561306 292170 561374 292226
rect 561430 292170 561498 292226
rect 561554 292170 561622 292226
rect 561678 292170 579250 292226
rect 579306 292170 579374 292226
rect 579430 292170 579498 292226
rect 579554 292170 579622 292226
rect 579678 292170 596496 292226
rect 596552 292170 596620 292226
rect 596676 292170 596744 292226
rect 596800 292170 596868 292226
rect 596924 292170 597980 292226
rect -1916 292102 597980 292170
rect -1916 292046 -860 292102
rect -804 292046 -736 292102
rect -680 292046 -612 292102
rect -556 292046 -488 292102
rect -432 292046 3250 292102
rect 3306 292046 3374 292102
rect 3430 292046 3498 292102
rect 3554 292046 3622 292102
rect 3678 292046 21250 292102
rect 21306 292046 21374 292102
rect 21430 292046 21498 292102
rect 21554 292046 21622 292102
rect 21678 292046 39250 292102
rect 39306 292046 39374 292102
rect 39430 292046 39498 292102
rect 39554 292046 39622 292102
rect 39678 292046 57250 292102
rect 57306 292046 57374 292102
rect 57430 292046 57498 292102
rect 57554 292046 57622 292102
rect 57678 292046 93250 292102
rect 93306 292046 93374 292102
rect 93430 292046 93498 292102
rect 93554 292046 93622 292102
rect 93678 292046 111250 292102
rect 111306 292046 111374 292102
rect 111430 292046 111498 292102
rect 111554 292046 111622 292102
rect 111678 292046 129250 292102
rect 129306 292046 129374 292102
rect 129430 292046 129498 292102
rect 129554 292046 129622 292102
rect 129678 292046 147250 292102
rect 147306 292046 147374 292102
rect 147430 292046 147498 292102
rect 147554 292046 147622 292102
rect 147678 292046 183250 292102
rect 183306 292046 183374 292102
rect 183430 292046 183498 292102
rect 183554 292046 183622 292102
rect 183678 292046 201250 292102
rect 201306 292046 201374 292102
rect 201430 292046 201498 292102
rect 201554 292046 201622 292102
rect 201678 292046 219250 292102
rect 219306 292046 219374 292102
rect 219430 292046 219498 292102
rect 219554 292046 219622 292102
rect 219678 292046 237250 292102
rect 237306 292046 237374 292102
rect 237430 292046 237498 292102
rect 237554 292046 237622 292102
rect 237678 292046 273250 292102
rect 273306 292046 273374 292102
rect 273430 292046 273498 292102
rect 273554 292046 273622 292102
rect 273678 292046 291250 292102
rect 291306 292046 291374 292102
rect 291430 292046 291498 292102
rect 291554 292046 291622 292102
rect 291678 292046 309250 292102
rect 309306 292046 309374 292102
rect 309430 292046 309498 292102
rect 309554 292046 309622 292102
rect 309678 292046 327250 292102
rect 327306 292046 327374 292102
rect 327430 292046 327498 292102
rect 327554 292046 327622 292102
rect 327678 292046 363250 292102
rect 363306 292046 363374 292102
rect 363430 292046 363498 292102
rect 363554 292046 363622 292102
rect 363678 292046 381250 292102
rect 381306 292046 381374 292102
rect 381430 292046 381498 292102
rect 381554 292046 381622 292102
rect 381678 292046 399250 292102
rect 399306 292046 399374 292102
rect 399430 292046 399498 292102
rect 399554 292046 399622 292102
rect 399678 292046 417250 292102
rect 417306 292046 417374 292102
rect 417430 292046 417498 292102
rect 417554 292046 417622 292102
rect 417678 292046 453250 292102
rect 453306 292046 453374 292102
rect 453430 292046 453498 292102
rect 453554 292046 453622 292102
rect 453678 292046 471250 292102
rect 471306 292046 471374 292102
rect 471430 292046 471498 292102
rect 471554 292046 471622 292102
rect 471678 292046 489250 292102
rect 489306 292046 489374 292102
rect 489430 292046 489498 292102
rect 489554 292046 489622 292102
rect 489678 292046 507250 292102
rect 507306 292046 507374 292102
rect 507430 292046 507498 292102
rect 507554 292046 507622 292102
rect 507678 292046 543250 292102
rect 543306 292046 543374 292102
rect 543430 292046 543498 292102
rect 543554 292046 543622 292102
rect 543678 292046 561250 292102
rect 561306 292046 561374 292102
rect 561430 292046 561498 292102
rect 561554 292046 561622 292102
rect 561678 292046 579250 292102
rect 579306 292046 579374 292102
rect 579430 292046 579498 292102
rect 579554 292046 579622 292102
rect 579678 292046 596496 292102
rect 596552 292046 596620 292102
rect 596676 292046 596744 292102
rect 596800 292046 596868 292102
rect 596924 292046 597980 292102
rect -1916 291978 597980 292046
rect -1916 291922 -860 291978
rect -804 291922 -736 291978
rect -680 291922 -612 291978
rect -556 291922 -488 291978
rect -432 291922 3250 291978
rect 3306 291922 3374 291978
rect 3430 291922 3498 291978
rect 3554 291922 3622 291978
rect 3678 291922 21250 291978
rect 21306 291922 21374 291978
rect 21430 291922 21498 291978
rect 21554 291922 21622 291978
rect 21678 291922 39250 291978
rect 39306 291922 39374 291978
rect 39430 291922 39498 291978
rect 39554 291922 39622 291978
rect 39678 291922 57250 291978
rect 57306 291922 57374 291978
rect 57430 291922 57498 291978
rect 57554 291922 57622 291978
rect 57678 291922 93250 291978
rect 93306 291922 93374 291978
rect 93430 291922 93498 291978
rect 93554 291922 93622 291978
rect 93678 291922 111250 291978
rect 111306 291922 111374 291978
rect 111430 291922 111498 291978
rect 111554 291922 111622 291978
rect 111678 291922 129250 291978
rect 129306 291922 129374 291978
rect 129430 291922 129498 291978
rect 129554 291922 129622 291978
rect 129678 291922 147250 291978
rect 147306 291922 147374 291978
rect 147430 291922 147498 291978
rect 147554 291922 147622 291978
rect 147678 291922 183250 291978
rect 183306 291922 183374 291978
rect 183430 291922 183498 291978
rect 183554 291922 183622 291978
rect 183678 291922 201250 291978
rect 201306 291922 201374 291978
rect 201430 291922 201498 291978
rect 201554 291922 201622 291978
rect 201678 291922 219250 291978
rect 219306 291922 219374 291978
rect 219430 291922 219498 291978
rect 219554 291922 219622 291978
rect 219678 291922 237250 291978
rect 237306 291922 237374 291978
rect 237430 291922 237498 291978
rect 237554 291922 237622 291978
rect 237678 291922 273250 291978
rect 273306 291922 273374 291978
rect 273430 291922 273498 291978
rect 273554 291922 273622 291978
rect 273678 291922 291250 291978
rect 291306 291922 291374 291978
rect 291430 291922 291498 291978
rect 291554 291922 291622 291978
rect 291678 291922 309250 291978
rect 309306 291922 309374 291978
rect 309430 291922 309498 291978
rect 309554 291922 309622 291978
rect 309678 291922 327250 291978
rect 327306 291922 327374 291978
rect 327430 291922 327498 291978
rect 327554 291922 327622 291978
rect 327678 291922 363250 291978
rect 363306 291922 363374 291978
rect 363430 291922 363498 291978
rect 363554 291922 363622 291978
rect 363678 291922 381250 291978
rect 381306 291922 381374 291978
rect 381430 291922 381498 291978
rect 381554 291922 381622 291978
rect 381678 291922 399250 291978
rect 399306 291922 399374 291978
rect 399430 291922 399498 291978
rect 399554 291922 399622 291978
rect 399678 291922 417250 291978
rect 417306 291922 417374 291978
rect 417430 291922 417498 291978
rect 417554 291922 417622 291978
rect 417678 291922 453250 291978
rect 453306 291922 453374 291978
rect 453430 291922 453498 291978
rect 453554 291922 453622 291978
rect 453678 291922 471250 291978
rect 471306 291922 471374 291978
rect 471430 291922 471498 291978
rect 471554 291922 471622 291978
rect 471678 291922 489250 291978
rect 489306 291922 489374 291978
rect 489430 291922 489498 291978
rect 489554 291922 489622 291978
rect 489678 291922 507250 291978
rect 507306 291922 507374 291978
rect 507430 291922 507498 291978
rect 507554 291922 507622 291978
rect 507678 291922 543250 291978
rect 543306 291922 543374 291978
rect 543430 291922 543498 291978
rect 543554 291922 543622 291978
rect 543678 291922 561250 291978
rect 561306 291922 561374 291978
rect 561430 291922 561498 291978
rect 561554 291922 561622 291978
rect 561678 291922 579250 291978
rect 579306 291922 579374 291978
rect 579430 291922 579498 291978
rect 579554 291922 579622 291978
rect 579678 291922 596496 291978
rect 596552 291922 596620 291978
rect 596676 291922 596744 291978
rect 596800 291922 596868 291978
rect 596924 291922 597980 291978
rect -1916 291826 597980 291922
rect -1916 280350 597980 280446
rect -1916 280294 -1820 280350
rect -1764 280294 -1696 280350
rect -1640 280294 -1572 280350
rect -1516 280294 -1448 280350
rect -1392 280294 6970 280350
rect 7026 280294 7094 280350
rect 7150 280294 7218 280350
rect 7274 280294 7342 280350
rect 7398 280294 24970 280350
rect 25026 280294 25094 280350
rect 25150 280294 25218 280350
rect 25274 280294 25342 280350
rect 25398 280294 42970 280350
rect 43026 280294 43094 280350
rect 43150 280294 43218 280350
rect 43274 280294 43342 280350
rect 43398 280294 60970 280350
rect 61026 280294 61094 280350
rect 61150 280294 61218 280350
rect 61274 280294 61342 280350
rect 61398 280294 78970 280350
rect 79026 280294 79094 280350
rect 79150 280294 79218 280350
rect 79274 280294 79342 280350
rect 79398 280294 96970 280350
rect 97026 280294 97094 280350
rect 97150 280294 97218 280350
rect 97274 280294 97342 280350
rect 97398 280294 132970 280350
rect 133026 280294 133094 280350
rect 133150 280294 133218 280350
rect 133274 280294 133342 280350
rect 133398 280294 150970 280350
rect 151026 280294 151094 280350
rect 151150 280294 151218 280350
rect 151274 280294 151342 280350
rect 151398 280294 168970 280350
rect 169026 280294 169094 280350
rect 169150 280294 169218 280350
rect 169274 280294 169342 280350
rect 169398 280294 186970 280350
rect 187026 280294 187094 280350
rect 187150 280294 187218 280350
rect 187274 280294 187342 280350
rect 187398 280294 222970 280350
rect 223026 280294 223094 280350
rect 223150 280294 223218 280350
rect 223274 280294 223342 280350
rect 223398 280294 240970 280350
rect 241026 280294 241094 280350
rect 241150 280294 241218 280350
rect 241274 280294 241342 280350
rect 241398 280294 258970 280350
rect 259026 280294 259094 280350
rect 259150 280294 259218 280350
rect 259274 280294 259342 280350
rect 259398 280294 276970 280350
rect 277026 280294 277094 280350
rect 277150 280294 277218 280350
rect 277274 280294 277342 280350
rect 277398 280294 312970 280350
rect 313026 280294 313094 280350
rect 313150 280294 313218 280350
rect 313274 280294 313342 280350
rect 313398 280294 330970 280350
rect 331026 280294 331094 280350
rect 331150 280294 331218 280350
rect 331274 280294 331342 280350
rect 331398 280294 348970 280350
rect 349026 280294 349094 280350
rect 349150 280294 349218 280350
rect 349274 280294 349342 280350
rect 349398 280294 366970 280350
rect 367026 280294 367094 280350
rect 367150 280294 367218 280350
rect 367274 280294 367342 280350
rect 367398 280294 402970 280350
rect 403026 280294 403094 280350
rect 403150 280294 403218 280350
rect 403274 280294 403342 280350
rect 403398 280294 420970 280350
rect 421026 280294 421094 280350
rect 421150 280294 421218 280350
rect 421274 280294 421342 280350
rect 421398 280294 438970 280350
rect 439026 280294 439094 280350
rect 439150 280294 439218 280350
rect 439274 280294 439342 280350
rect 439398 280294 456970 280350
rect 457026 280294 457094 280350
rect 457150 280294 457218 280350
rect 457274 280294 457342 280350
rect 457398 280294 492970 280350
rect 493026 280294 493094 280350
rect 493150 280294 493218 280350
rect 493274 280294 493342 280350
rect 493398 280294 510970 280350
rect 511026 280294 511094 280350
rect 511150 280294 511218 280350
rect 511274 280294 511342 280350
rect 511398 280294 528970 280350
rect 529026 280294 529094 280350
rect 529150 280294 529218 280350
rect 529274 280294 529342 280350
rect 529398 280294 546970 280350
rect 547026 280294 547094 280350
rect 547150 280294 547218 280350
rect 547274 280294 547342 280350
rect 547398 280294 564970 280350
rect 565026 280294 565094 280350
rect 565150 280294 565218 280350
rect 565274 280294 565342 280350
rect 565398 280294 582970 280350
rect 583026 280294 583094 280350
rect 583150 280294 583218 280350
rect 583274 280294 583342 280350
rect 583398 280294 597456 280350
rect 597512 280294 597580 280350
rect 597636 280294 597704 280350
rect 597760 280294 597828 280350
rect 597884 280294 597980 280350
rect -1916 280226 597980 280294
rect -1916 280170 -1820 280226
rect -1764 280170 -1696 280226
rect -1640 280170 -1572 280226
rect -1516 280170 -1448 280226
rect -1392 280170 6970 280226
rect 7026 280170 7094 280226
rect 7150 280170 7218 280226
rect 7274 280170 7342 280226
rect 7398 280170 24970 280226
rect 25026 280170 25094 280226
rect 25150 280170 25218 280226
rect 25274 280170 25342 280226
rect 25398 280170 42970 280226
rect 43026 280170 43094 280226
rect 43150 280170 43218 280226
rect 43274 280170 43342 280226
rect 43398 280170 60970 280226
rect 61026 280170 61094 280226
rect 61150 280170 61218 280226
rect 61274 280170 61342 280226
rect 61398 280170 78970 280226
rect 79026 280170 79094 280226
rect 79150 280170 79218 280226
rect 79274 280170 79342 280226
rect 79398 280170 96970 280226
rect 97026 280170 97094 280226
rect 97150 280170 97218 280226
rect 97274 280170 97342 280226
rect 97398 280170 132970 280226
rect 133026 280170 133094 280226
rect 133150 280170 133218 280226
rect 133274 280170 133342 280226
rect 133398 280170 150970 280226
rect 151026 280170 151094 280226
rect 151150 280170 151218 280226
rect 151274 280170 151342 280226
rect 151398 280170 168970 280226
rect 169026 280170 169094 280226
rect 169150 280170 169218 280226
rect 169274 280170 169342 280226
rect 169398 280170 186970 280226
rect 187026 280170 187094 280226
rect 187150 280170 187218 280226
rect 187274 280170 187342 280226
rect 187398 280170 222970 280226
rect 223026 280170 223094 280226
rect 223150 280170 223218 280226
rect 223274 280170 223342 280226
rect 223398 280170 240970 280226
rect 241026 280170 241094 280226
rect 241150 280170 241218 280226
rect 241274 280170 241342 280226
rect 241398 280170 258970 280226
rect 259026 280170 259094 280226
rect 259150 280170 259218 280226
rect 259274 280170 259342 280226
rect 259398 280170 276970 280226
rect 277026 280170 277094 280226
rect 277150 280170 277218 280226
rect 277274 280170 277342 280226
rect 277398 280170 312970 280226
rect 313026 280170 313094 280226
rect 313150 280170 313218 280226
rect 313274 280170 313342 280226
rect 313398 280170 330970 280226
rect 331026 280170 331094 280226
rect 331150 280170 331218 280226
rect 331274 280170 331342 280226
rect 331398 280170 348970 280226
rect 349026 280170 349094 280226
rect 349150 280170 349218 280226
rect 349274 280170 349342 280226
rect 349398 280170 366970 280226
rect 367026 280170 367094 280226
rect 367150 280170 367218 280226
rect 367274 280170 367342 280226
rect 367398 280170 402970 280226
rect 403026 280170 403094 280226
rect 403150 280170 403218 280226
rect 403274 280170 403342 280226
rect 403398 280170 420970 280226
rect 421026 280170 421094 280226
rect 421150 280170 421218 280226
rect 421274 280170 421342 280226
rect 421398 280170 438970 280226
rect 439026 280170 439094 280226
rect 439150 280170 439218 280226
rect 439274 280170 439342 280226
rect 439398 280170 456970 280226
rect 457026 280170 457094 280226
rect 457150 280170 457218 280226
rect 457274 280170 457342 280226
rect 457398 280170 492970 280226
rect 493026 280170 493094 280226
rect 493150 280170 493218 280226
rect 493274 280170 493342 280226
rect 493398 280170 510970 280226
rect 511026 280170 511094 280226
rect 511150 280170 511218 280226
rect 511274 280170 511342 280226
rect 511398 280170 528970 280226
rect 529026 280170 529094 280226
rect 529150 280170 529218 280226
rect 529274 280170 529342 280226
rect 529398 280170 546970 280226
rect 547026 280170 547094 280226
rect 547150 280170 547218 280226
rect 547274 280170 547342 280226
rect 547398 280170 564970 280226
rect 565026 280170 565094 280226
rect 565150 280170 565218 280226
rect 565274 280170 565342 280226
rect 565398 280170 582970 280226
rect 583026 280170 583094 280226
rect 583150 280170 583218 280226
rect 583274 280170 583342 280226
rect 583398 280170 597456 280226
rect 597512 280170 597580 280226
rect 597636 280170 597704 280226
rect 597760 280170 597828 280226
rect 597884 280170 597980 280226
rect -1916 280102 597980 280170
rect -1916 280046 -1820 280102
rect -1764 280046 -1696 280102
rect -1640 280046 -1572 280102
rect -1516 280046 -1448 280102
rect -1392 280046 6970 280102
rect 7026 280046 7094 280102
rect 7150 280046 7218 280102
rect 7274 280046 7342 280102
rect 7398 280046 24970 280102
rect 25026 280046 25094 280102
rect 25150 280046 25218 280102
rect 25274 280046 25342 280102
rect 25398 280046 42970 280102
rect 43026 280046 43094 280102
rect 43150 280046 43218 280102
rect 43274 280046 43342 280102
rect 43398 280046 60970 280102
rect 61026 280046 61094 280102
rect 61150 280046 61218 280102
rect 61274 280046 61342 280102
rect 61398 280046 78970 280102
rect 79026 280046 79094 280102
rect 79150 280046 79218 280102
rect 79274 280046 79342 280102
rect 79398 280046 96970 280102
rect 97026 280046 97094 280102
rect 97150 280046 97218 280102
rect 97274 280046 97342 280102
rect 97398 280046 132970 280102
rect 133026 280046 133094 280102
rect 133150 280046 133218 280102
rect 133274 280046 133342 280102
rect 133398 280046 150970 280102
rect 151026 280046 151094 280102
rect 151150 280046 151218 280102
rect 151274 280046 151342 280102
rect 151398 280046 168970 280102
rect 169026 280046 169094 280102
rect 169150 280046 169218 280102
rect 169274 280046 169342 280102
rect 169398 280046 186970 280102
rect 187026 280046 187094 280102
rect 187150 280046 187218 280102
rect 187274 280046 187342 280102
rect 187398 280046 222970 280102
rect 223026 280046 223094 280102
rect 223150 280046 223218 280102
rect 223274 280046 223342 280102
rect 223398 280046 240970 280102
rect 241026 280046 241094 280102
rect 241150 280046 241218 280102
rect 241274 280046 241342 280102
rect 241398 280046 258970 280102
rect 259026 280046 259094 280102
rect 259150 280046 259218 280102
rect 259274 280046 259342 280102
rect 259398 280046 276970 280102
rect 277026 280046 277094 280102
rect 277150 280046 277218 280102
rect 277274 280046 277342 280102
rect 277398 280046 312970 280102
rect 313026 280046 313094 280102
rect 313150 280046 313218 280102
rect 313274 280046 313342 280102
rect 313398 280046 330970 280102
rect 331026 280046 331094 280102
rect 331150 280046 331218 280102
rect 331274 280046 331342 280102
rect 331398 280046 348970 280102
rect 349026 280046 349094 280102
rect 349150 280046 349218 280102
rect 349274 280046 349342 280102
rect 349398 280046 366970 280102
rect 367026 280046 367094 280102
rect 367150 280046 367218 280102
rect 367274 280046 367342 280102
rect 367398 280046 402970 280102
rect 403026 280046 403094 280102
rect 403150 280046 403218 280102
rect 403274 280046 403342 280102
rect 403398 280046 420970 280102
rect 421026 280046 421094 280102
rect 421150 280046 421218 280102
rect 421274 280046 421342 280102
rect 421398 280046 438970 280102
rect 439026 280046 439094 280102
rect 439150 280046 439218 280102
rect 439274 280046 439342 280102
rect 439398 280046 456970 280102
rect 457026 280046 457094 280102
rect 457150 280046 457218 280102
rect 457274 280046 457342 280102
rect 457398 280046 492970 280102
rect 493026 280046 493094 280102
rect 493150 280046 493218 280102
rect 493274 280046 493342 280102
rect 493398 280046 510970 280102
rect 511026 280046 511094 280102
rect 511150 280046 511218 280102
rect 511274 280046 511342 280102
rect 511398 280046 528970 280102
rect 529026 280046 529094 280102
rect 529150 280046 529218 280102
rect 529274 280046 529342 280102
rect 529398 280046 546970 280102
rect 547026 280046 547094 280102
rect 547150 280046 547218 280102
rect 547274 280046 547342 280102
rect 547398 280046 564970 280102
rect 565026 280046 565094 280102
rect 565150 280046 565218 280102
rect 565274 280046 565342 280102
rect 565398 280046 582970 280102
rect 583026 280046 583094 280102
rect 583150 280046 583218 280102
rect 583274 280046 583342 280102
rect 583398 280046 597456 280102
rect 597512 280046 597580 280102
rect 597636 280046 597704 280102
rect 597760 280046 597828 280102
rect 597884 280046 597980 280102
rect -1916 279978 597980 280046
rect -1916 279922 -1820 279978
rect -1764 279922 -1696 279978
rect -1640 279922 -1572 279978
rect -1516 279922 -1448 279978
rect -1392 279922 6970 279978
rect 7026 279922 7094 279978
rect 7150 279922 7218 279978
rect 7274 279922 7342 279978
rect 7398 279922 24970 279978
rect 25026 279922 25094 279978
rect 25150 279922 25218 279978
rect 25274 279922 25342 279978
rect 25398 279922 42970 279978
rect 43026 279922 43094 279978
rect 43150 279922 43218 279978
rect 43274 279922 43342 279978
rect 43398 279922 60970 279978
rect 61026 279922 61094 279978
rect 61150 279922 61218 279978
rect 61274 279922 61342 279978
rect 61398 279922 78970 279978
rect 79026 279922 79094 279978
rect 79150 279922 79218 279978
rect 79274 279922 79342 279978
rect 79398 279922 96970 279978
rect 97026 279922 97094 279978
rect 97150 279922 97218 279978
rect 97274 279922 97342 279978
rect 97398 279922 132970 279978
rect 133026 279922 133094 279978
rect 133150 279922 133218 279978
rect 133274 279922 133342 279978
rect 133398 279922 150970 279978
rect 151026 279922 151094 279978
rect 151150 279922 151218 279978
rect 151274 279922 151342 279978
rect 151398 279922 168970 279978
rect 169026 279922 169094 279978
rect 169150 279922 169218 279978
rect 169274 279922 169342 279978
rect 169398 279922 186970 279978
rect 187026 279922 187094 279978
rect 187150 279922 187218 279978
rect 187274 279922 187342 279978
rect 187398 279922 222970 279978
rect 223026 279922 223094 279978
rect 223150 279922 223218 279978
rect 223274 279922 223342 279978
rect 223398 279922 240970 279978
rect 241026 279922 241094 279978
rect 241150 279922 241218 279978
rect 241274 279922 241342 279978
rect 241398 279922 258970 279978
rect 259026 279922 259094 279978
rect 259150 279922 259218 279978
rect 259274 279922 259342 279978
rect 259398 279922 276970 279978
rect 277026 279922 277094 279978
rect 277150 279922 277218 279978
rect 277274 279922 277342 279978
rect 277398 279922 312970 279978
rect 313026 279922 313094 279978
rect 313150 279922 313218 279978
rect 313274 279922 313342 279978
rect 313398 279922 330970 279978
rect 331026 279922 331094 279978
rect 331150 279922 331218 279978
rect 331274 279922 331342 279978
rect 331398 279922 348970 279978
rect 349026 279922 349094 279978
rect 349150 279922 349218 279978
rect 349274 279922 349342 279978
rect 349398 279922 366970 279978
rect 367026 279922 367094 279978
rect 367150 279922 367218 279978
rect 367274 279922 367342 279978
rect 367398 279922 402970 279978
rect 403026 279922 403094 279978
rect 403150 279922 403218 279978
rect 403274 279922 403342 279978
rect 403398 279922 420970 279978
rect 421026 279922 421094 279978
rect 421150 279922 421218 279978
rect 421274 279922 421342 279978
rect 421398 279922 438970 279978
rect 439026 279922 439094 279978
rect 439150 279922 439218 279978
rect 439274 279922 439342 279978
rect 439398 279922 456970 279978
rect 457026 279922 457094 279978
rect 457150 279922 457218 279978
rect 457274 279922 457342 279978
rect 457398 279922 492970 279978
rect 493026 279922 493094 279978
rect 493150 279922 493218 279978
rect 493274 279922 493342 279978
rect 493398 279922 510970 279978
rect 511026 279922 511094 279978
rect 511150 279922 511218 279978
rect 511274 279922 511342 279978
rect 511398 279922 528970 279978
rect 529026 279922 529094 279978
rect 529150 279922 529218 279978
rect 529274 279922 529342 279978
rect 529398 279922 546970 279978
rect 547026 279922 547094 279978
rect 547150 279922 547218 279978
rect 547274 279922 547342 279978
rect 547398 279922 564970 279978
rect 565026 279922 565094 279978
rect 565150 279922 565218 279978
rect 565274 279922 565342 279978
rect 565398 279922 582970 279978
rect 583026 279922 583094 279978
rect 583150 279922 583218 279978
rect 583274 279922 583342 279978
rect 583398 279922 597456 279978
rect 597512 279922 597580 279978
rect 597636 279922 597704 279978
rect 597760 279922 597828 279978
rect 597884 279922 597980 279978
rect -1916 279826 597980 279922
rect -1916 274350 597980 274446
rect -1916 274294 -860 274350
rect -804 274294 -736 274350
rect -680 274294 -612 274350
rect -556 274294 -488 274350
rect -432 274294 3250 274350
rect 3306 274294 3374 274350
rect 3430 274294 3498 274350
rect 3554 274294 3622 274350
rect 3678 274294 21250 274350
rect 21306 274294 21374 274350
rect 21430 274294 21498 274350
rect 21554 274294 21622 274350
rect 21678 274294 39250 274350
rect 39306 274294 39374 274350
rect 39430 274294 39498 274350
rect 39554 274294 39622 274350
rect 39678 274294 57250 274350
rect 57306 274294 57374 274350
rect 57430 274294 57498 274350
rect 57554 274294 57622 274350
rect 57678 274294 93250 274350
rect 93306 274294 93374 274350
rect 93430 274294 93498 274350
rect 93554 274294 93622 274350
rect 93678 274294 111250 274350
rect 111306 274294 111374 274350
rect 111430 274294 111498 274350
rect 111554 274294 111622 274350
rect 111678 274294 129250 274350
rect 129306 274294 129374 274350
rect 129430 274294 129498 274350
rect 129554 274294 129622 274350
rect 129678 274294 147250 274350
rect 147306 274294 147374 274350
rect 147430 274294 147498 274350
rect 147554 274294 147622 274350
rect 147678 274294 183250 274350
rect 183306 274294 183374 274350
rect 183430 274294 183498 274350
rect 183554 274294 183622 274350
rect 183678 274294 201250 274350
rect 201306 274294 201374 274350
rect 201430 274294 201498 274350
rect 201554 274294 201622 274350
rect 201678 274294 219250 274350
rect 219306 274294 219374 274350
rect 219430 274294 219498 274350
rect 219554 274294 219622 274350
rect 219678 274294 237250 274350
rect 237306 274294 237374 274350
rect 237430 274294 237498 274350
rect 237554 274294 237622 274350
rect 237678 274294 273250 274350
rect 273306 274294 273374 274350
rect 273430 274294 273498 274350
rect 273554 274294 273622 274350
rect 273678 274294 291250 274350
rect 291306 274294 291374 274350
rect 291430 274294 291498 274350
rect 291554 274294 291622 274350
rect 291678 274294 309250 274350
rect 309306 274294 309374 274350
rect 309430 274294 309498 274350
rect 309554 274294 309622 274350
rect 309678 274294 327250 274350
rect 327306 274294 327374 274350
rect 327430 274294 327498 274350
rect 327554 274294 327622 274350
rect 327678 274294 363250 274350
rect 363306 274294 363374 274350
rect 363430 274294 363498 274350
rect 363554 274294 363622 274350
rect 363678 274294 381250 274350
rect 381306 274294 381374 274350
rect 381430 274294 381498 274350
rect 381554 274294 381622 274350
rect 381678 274294 399250 274350
rect 399306 274294 399374 274350
rect 399430 274294 399498 274350
rect 399554 274294 399622 274350
rect 399678 274294 417250 274350
rect 417306 274294 417374 274350
rect 417430 274294 417498 274350
rect 417554 274294 417622 274350
rect 417678 274294 453250 274350
rect 453306 274294 453374 274350
rect 453430 274294 453498 274350
rect 453554 274294 453622 274350
rect 453678 274294 471250 274350
rect 471306 274294 471374 274350
rect 471430 274294 471498 274350
rect 471554 274294 471622 274350
rect 471678 274294 489250 274350
rect 489306 274294 489374 274350
rect 489430 274294 489498 274350
rect 489554 274294 489622 274350
rect 489678 274294 507250 274350
rect 507306 274294 507374 274350
rect 507430 274294 507498 274350
rect 507554 274294 507622 274350
rect 507678 274294 543250 274350
rect 543306 274294 543374 274350
rect 543430 274294 543498 274350
rect 543554 274294 543622 274350
rect 543678 274294 561250 274350
rect 561306 274294 561374 274350
rect 561430 274294 561498 274350
rect 561554 274294 561622 274350
rect 561678 274294 579250 274350
rect 579306 274294 579374 274350
rect 579430 274294 579498 274350
rect 579554 274294 579622 274350
rect 579678 274294 596496 274350
rect 596552 274294 596620 274350
rect 596676 274294 596744 274350
rect 596800 274294 596868 274350
rect 596924 274294 597980 274350
rect -1916 274226 597980 274294
rect -1916 274170 -860 274226
rect -804 274170 -736 274226
rect -680 274170 -612 274226
rect -556 274170 -488 274226
rect -432 274170 3250 274226
rect 3306 274170 3374 274226
rect 3430 274170 3498 274226
rect 3554 274170 3622 274226
rect 3678 274170 21250 274226
rect 21306 274170 21374 274226
rect 21430 274170 21498 274226
rect 21554 274170 21622 274226
rect 21678 274170 39250 274226
rect 39306 274170 39374 274226
rect 39430 274170 39498 274226
rect 39554 274170 39622 274226
rect 39678 274170 57250 274226
rect 57306 274170 57374 274226
rect 57430 274170 57498 274226
rect 57554 274170 57622 274226
rect 57678 274170 93250 274226
rect 93306 274170 93374 274226
rect 93430 274170 93498 274226
rect 93554 274170 93622 274226
rect 93678 274170 111250 274226
rect 111306 274170 111374 274226
rect 111430 274170 111498 274226
rect 111554 274170 111622 274226
rect 111678 274170 129250 274226
rect 129306 274170 129374 274226
rect 129430 274170 129498 274226
rect 129554 274170 129622 274226
rect 129678 274170 147250 274226
rect 147306 274170 147374 274226
rect 147430 274170 147498 274226
rect 147554 274170 147622 274226
rect 147678 274170 183250 274226
rect 183306 274170 183374 274226
rect 183430 274170 183498 274226
rect 183554 274170 183622 274226
rect 183678 274170 201250 274226
rect 201306 274170 201374 274226
rect 201430 274170 201498 274226
rect 201554 274170 201622 274226
rect 201678 274170 219250 274226
rect 219306 274170 219374 274226
rect 219430 274170 219498 274226
rect 219554 274170 219622 274226
rect 219678 274170 237250 274226
rect 237306 274170 237374 274226
rect 237430 274170 237498 274226
rect 237554 274170 237622 274226
rect 237678 274170 273250 274226
rect 273306 274170 273374 274226
rect 273430 274170 273498 274226
rect 273554 274170 273622 274226
rect 273678 274170 291250 274226
rect 291306 274170 291374 274226
rect 291430 274170 291498 274226
rect 291554 274170 291622 274226
rect 291678 274170 309250 274226
rect 309306 274170 309374 274226
rect 309430 274170 309498 274226
rect 309554 274170 309622 274226
rect 309678 274170 327250 274226
rect 327306 274170 327374 274226
rect 327430 274170 327498 274226
rect 327554 274170 327622 274226
rect 327678 274170 363250 274226
rect 363306 274170 363374 274226
rect 363430 274170 363498 274226
rect 363554 274170 363622 274226
rect 363678 274170 381250 274226
rect 381306 274170 381374 274226
rect 381430 274170 381498 274226
rect 381554 274170 381622 274226
rect 381678 274170 399250 274226
rect 399306 274170 399374 274226
rect 399430 274170 399498 274226
rect 399554 274170 399622 274226
rect 399678 274170 417250 274226
rect 417306 274170 417374 274226
rect 417430 274170 417498 274226
rect 417554 274170 417622 274226
rect 417678 274170 453250 274226
rect 453306 274170 453374 274226
rect 453430 274170 453498 274226
rect 453554 274170 453622 274226
rect 453678 274170 471250 274226
rect 471306 274170 471374 274226
rect 471430 274170 471498 274226
rect 471554 274170 471622 274226
rect 471678 274170 489250 274226
rect 489306 274170 489374 274226
rect 489430 274170 489498 274226
rect 489554 274170 489622 274226
rect 489678 274170 507250 274226
rect 507306 274170 507374 274226
rect 507430 274170 507498 274226
rect 507554 274170 507622 274226
rect 507678 274170 543250 274226
rect 543306 274170 543374 274226
rect 543430 274170 543498 274226
rect 543554 274170 543622 274226
rect 543678 274170 561250 274226
rect 561306 274170 561374 274226
rect 561430 274170 561498 274226
rect 561554 274170 561622 274226
rect 561678 274170 579250 274226
rect 579306 274170 579374 274226
rect 579430 274170 579498 274226
rect 579554 274170 579622 274226
rect 579678 274170 596496 274226
rect 596552 274170 596620 274226
rect 596676 274170 596744 274226
rect 596800 274170 596868 274226
rect 596924 274170 597980 274226
rect -1916 274102 597980 274170
rect -1916 274046 -860 274102
rect -804 274046 -736 274102
rect -680 274046 -612 274102
rect -556 274046 -488 274102
rect -432 274046 3250 274102
rect 3306 274046 3374 274102
rect 3430 274046 3498 274102
rect 3554 274046 3622 274102
rect 3678 274046 21250 274102
rect 21306 274046 21374 274102
rect 21430 274046 21498 274102
rect 21554 274046 21622 274102
rect 21678 274046 39250 274102
rect 39306 274046 39374 274102
rect 39430 274046 39498 274102
rect 39554 274046 39622 274102
rect 39678 274046 57250 274102
rect 57306 274046 57374 274102
rect 57430 274046 57498 274102
rect 57554 274046 57622 274102
rect 57678 274046 93250 274102
rect 93306 274046 93374 274102
rect 93430 274046 93498 274102
rect 93554 274046 93622 274102
rect 93678 274046 111250 274102
rect 111306 274046 111374 274102
rect 111430 274046 111498 274102
rect 111554 274046 111622 274102
rect 111678 274046 129250 274102
rect 129306 274046 129374 274102
rect 129430 274046 129498 274102
rect 129554 274046 129622 274102
rect 129678 274046 147250 274102
rect 147306 274046 147374 274102
rect 147430 274046 147498 274102
rect 147554 274046 147622 274102
rect 147678 274046 183250 274102
rect 183306 274046 183374 274102
rect 183430 274046 183498 274102
rect 183554 274046 183622 274102
rect 183678 274046 201250 274102
rect 201306 274046 201374 274102
rect 201430 274046 201498 274102
rect 201554 274046 201622 274102
rect 201678 274046 219250 274102
rect 219306 274046 219374 274102
rect 219430 274046 219498 274102
rect 219554 274046 219622 274102
rect 219678 274046 237250 274102
rect 237306 274046 237374 274102
rect 237430 274046 237498 274102
rect 237554 274046 237622 274102
rect 237678 274046 273250 274102
rect 273306 274046 273374 274102
rect 273430 274046 273498 274102
rect 273554 274046 273622 274102
rect 273678 274046 291250 274102
rect 291306 274046 291374 274102
rect 291430 274046 291498 274102
rect 291554 274046 291622 274102
rect 291678 274046 309250 274102
rect 309306 274046 309374 274102
rect 309430 274046 309498 274102
rect 309554 274046 309622 274102
rect 309678 274046 327250 274102
rect 327306 274046 327374 274102
rect 327430 274046 327498 274102
rect 327554 274046 327622 274102
rect 327678 274046 363250 274102
rect 363306 274046 363374 274102
rect 363430 274046 363498 274102
rect 363554 274046 363622 274102
rect 363678 274046 381250 274102
rect 381306 274046 381374 274102
rect 381430 274046 381498 274102
rect 381554 274046 381622 274102
rect 381678 274046 399250 274102
rect 399306 274046 399374 274102
rect 399430 274046 399498 274102
rect 399554 274046 399622 274102
rect 399678 274046 417250 274102
rect 417306 274046 417374 274102
rect 417430 274046 417498 274102
rect 417554 274046 417622 274102
rect 417678 274046 453250 274102
rect 453306 274046 453374 274102
rect 453430 274046 453498 274102
rect 453554 274046 453622 274102
rect 453678 274046 471250 274102
rect 471306 274046 471374 274102
rect 471430 274046 471498 274102
rect 471554 274046 471622 274102
rect 471678 274046 489250 274102
rect 489306 274046 489374 274102
rect 489430 274046 489498 274102
rect 489554 274046 489622 274102
rect 489678 274046 507250 274102
rect 507306 274046 507374 274102
rect 507430 274046 507498 274102
rect 507554 274046 507622 274102
rect 507678 274046 543250 274102
rect 543306 274046 543374 274102
rect 543430 274046 543498 274102
rect 543554 274046 543622 274102
rect 543678 274046 561250 274102
rect 561306 274046 561374 274102
rect 561430 274046 561498 274102
rect 561554 274046 561622 274102
rect 561678 274046 579250 274102
rect 579306 274046 579374 274102
rect 579430 274046 579498 274102
rect 579554 274046 579622 274102
rect 579678 274046 596496 274102
rect 596552 274046 596620 274102
rect 596676 274046 596744 274102
rect 596800 274046 596868 274102
rect 596924 274046 597980 274102
rect -1916 273978 597980 274046
rect -1916 273922 -860 273978
rect -804 273922 -736 273978
rect -680 273922 -612 273978
rect -556 273922 -488 273978
rect -432 273922 3250 273978
rect 3306 273922 3374 273978
rect 3430 273922 3498 273978
rect 3554 273922 3622 273978
rect 3678 273922 21250 273978
rect 21306 273922 21374 273978
rect 21430 273922 21498 273978
rect 21554 273922 21622 273978
rect 21678 273922 39250 273978
rect 39306 273922 39374 273978
rect 39430 273922 39498 273978
rect 39554 273922 39622 273978
rect 39678 273922 57250 273978
rect 57306 273922 57374 273978
rect 57430 273922 57498 273978
rect 57554 273922 57622 273978
rect 57678 273922 93250 273978
rect 93306 273922 93374 273978
rect 93430 273922 93498 273978
rect 93554 273922 93622 273978
rect 93678 273922 111250 273978
rect 111306 273922 111374 273978
rect 111430 273922 111498 273978
rect 111554 273922 111622 273978
rect 111678 273922 129250 273978
rect 129306 273922 129374 273978
rect 129430 273922 129498 273978
rect 129554 273922 129622 273978
rect 129678 273922 147250 273978
rect 147306 273922 147374 273978
rect 147430 273922 147498 273978
rect 147554 273922 147622 273978
rect 147678 273922 183250 273978
rect 183306 273922 183374 273978
rect 183430 273922 183498 273978
rect 183554 273922 183622 273978
rect 183678 273922 201250 273978
rect 201306 273922 201374 273978
rect 201430 273922 201498 273978
rect 201554 273922 201622 273978
rect 201678 273922 219250 273978
rect 219306 273922 219374 273978
rect 219430 273922 219498 273978
rect 219554 273922 219622 273978
rect 219678 273922 237250 273978
rect 237306 273922 237374 273978
rect 237430 273922 237498 273978
rect 237554 273922 237622 273978
rect 237678 273922 273250 273978
rect 273306 273922 273374 273978
rect 273430 273922 273498 273978
rect 273554 273922 273622 273978
rect 273678 273922 291250 273978
rect 291306 273922 291374 273978
rect 291430 273922 291498 273978
rect 291554 273922 291622 273978
rect 291678 273922 309250 273978
rect 309306 273922 309374 273978
rect 309430 273922 309498 273978
rect 309554 273922 309622 273978
rect 309678 273922 327250 273978
rect 327306 273922 327374 273978
rect 327430 273922 327498 273978
rect 327554 273922 327622 273978
rect 327678 273922 363250 273978
rect 363306 273922 363374 273978
rect 363430 273922 363498 273978
rect 363554 273922 363622 273978
rect 363678 273922 381250 273978
rect 381306 273922 381374 273978
rect 381430 273922 381498 273978
rect 381554 273922 381622 273978
rect 381678 273922 399250 273978
rect 399306 273922 399374 273978
rect 399430 273922 399498 273978
rect 399554 273922 399622 273978
rect 399678 273922 417250 273978
rect 417306 273922 417374 273978
rect 417430 273922 417498 273978
rect 417554 273922 417622 273978
rect 417678 273922 453250 273978
rect 453306 273922 453374 273978
rect 453430 273922 453498 273978
rect 453554 273922 453622 273978
rect 453678 273922 471250 273978
rect 471306 273922 471374 273978
rect 471430 273922 471498 273978
rect 471554 273922 471622 273978
rect 471678 273922 489250 273978
rect 489306 273922 489374 273978
rect 489430 273922 489498 273978
rect 489554 273922 489622 273978
rect 489678 273922 507250 273978
rect 507306 273922 507374 273978
rect 507430 273922 507498 273978
rect 507554 273922 507622 273978
rect 507678 273922 543250 273978
rect 543306 273922 543374 273978
rect 543430 273922 543498 273978
rect 543554 273922 543622 273978
rect 543678 273922 561250 273978
rect 561306 273922 561374 273978
rect 561430 273922 561498 273978
rect 561554 273922 561622 273978
rect 561678 273922 579250 273978
rect 579306 273922 579374 273978
rect 579430 273922 579498 273978
rect 579554 273922 579622 273978
rect 579678 273922 596496 273978
rect 596552 273922 596620 273978
rect 596676 273922 596744 273978
rect 596800 273922 596868 273978
rect 596924 273922 597980 273978
rect -1916 273826 597980 273922
rect -1916 262350 597980 262446
rect -1916 262294 -1820 262350
rect -1764 262294 -1696 262350
rect -1640 262294 -1572 262350
rect -1516 262294 -1448 262350
rect -1392 262294 6970 262350
rect 7026 262294 7094 262350
rect 7150 262294 7218 262350
rect 7274 262294 7342 262350
rect 7398 262294 24970 262350
rect 25026 262294 25094 262350
rect 25150 262294 25218 262350
rect 25274 262294 25342 262350
rect 25398 262294 42970 262350
rect 43026 262294 43094 262350
rect 43150 262294 43218 262350
rect 43274 262294 43342 262350
rect 43398 262294 60970 262350
rect 61026 262294 61094 262350
rect 61150 262294 61218 262350
rect 61274 262294 61342 262350
rect 61398 262294 78970 262350
rect 79026 262294 79094 262350
rect 79150 262294 79218 262350
rect 79274 262294 79342 262350
rect 79398 262294 96970 262350
rect 97026 262294 97094 262350
rect 97150 262294 97218 262350
rect 97274 262294 97342 262350
rect 97398 262294 132970 262350
rect 133026 262294 133094 262350
rect 133150 262294 133218 262350
rect 133274 262294 133342 262350
rect 133398 262294 150970 262350
rect 151026 262294 151094 262350
rect 151150 262294 151218 262350
rect 151274 262294 151342 262350
rect 151398 262294 168970 262350
rect 169026 262294 169094 262350
rect 169150 262294 169218 262350
rect 169274 262294 169342 262350
rect 169398 262294 186970 262350
rect 187026 262294 187094 262350
rect 187150 262294 187218 262350
rect 187274 262294 187342 262350
rect 187398 262294 222970 262350
rect 223026 262294 223094 262350
rect 223150 262294 223218 262350
rect 223274 262294 223342 262350
rect 223398 262294 240970 262350
rect 241026 262294 241094 262350
rect 241150 262294 241218 262350
rect 241274 262294 241342 262350
rect 241398 262294 258970 262350
rect 259026 262294 259094 262350
rect 259150 262294 259218 262350
rect 259274 262294 259342 262350
rect 259398 262294 276970 262350
rect 277026 262294 277094 262350
rect 277150 262294 277218 262350
rect 277274 262294 277342 262350
rect 277398 262294 312970 262350
rect 313026 262294 313094 262350
rect 313150 262294 313218 262350
rect 313274 262294 313342 262350
rect 313398 262294 330970 262350
rect 331026 262294 331094 262350
rect 331150 262294 331218 262350
rect 331274 262294 331342 262350
rect 331398 262294 348970 262350
rect 349026 262294 349094 262350
rect 349150 262294 349218 262350
rect 349274 262294 349342 262350
rect 349398 262294 366970 262350
rect 367026 262294 367094 262350
rect 367150 262294 367218 262350
rect 367274 262294 367342 262350
rect 367398 262294 402970 262350
rect 403026 262294 403094 262350
rect 403150 262294 403218 262350
rect 403274 262294 403342 262350
rect 403398 262294 420970 262350
rect 421026 262294 421094 262350
rect 421150 262294 421218 262350
rect 421274 262294 421342 262350
rect 421398 262294 438970 262350
rect 439026 262294 439094 262350
rect 439150 262294 439218 262350
rect 439274 262294 439342 262350
rect 439398 262294 456970 262350
rect 457026 262294 457094 262350
rect 457150 262294 457218 262350
rect 457274 262294 457342 262350
rect 457398 262294 492970 262350
rect 493026 262294 493094 262350
rect 493150 262294 493218 262350
rect 493274 262294 493342 262350
rect 493398 262294 510970 262350
rect 511026 262294 511094 262350
rect 511150 262294 511218 262350
rect 511274 262294 511342 262350
rect 511398 262294 528970 262350
rect 529026 262294 529094 262350
rect 529150 262294 529218 262350
rect 529274 262294 529342 262350
rect 529398 262294 546970 262350
rect 547026 262294 547094 262350
rect 547150 262294 547218 262350
rect 547274 262294 547342 262350
rect 547398 262294 564970 262350
rect 565026 262294 565094 262350
rect 565150 262294 565218 262350
rect 565274 262294 565342 262350
rect 565398 262294 582970 262350
rect 583026 262294 583094 262350
rect 583150 262294 583218 262350
rect 583274 262294 583342 262350
rect 583398 262294 597456 262350
rect 597512 262294 597580 262350
rect 597636 262294 597704 262350
rect 597760 262294 597828 262350
rect 597884 262294 597980 262350
rect -1916 262226 597980 262294
rect -1916 262170 -1820 262226
rect -1764 262170 -1696 262226
rect -1640 262170 -1572 262226
rect -1516 262170 -1448 262226
rect -1392 262170 6970 262226
rect 7026 262170 7094 262226
rect 7150 262170 7218 262226
rect 7274 262170 7342 262226
rect 7398 262170 24970 262226
rect 25026 262170 25094 262226
rect 25150 262170 25218 262226
rect 25274 262170 25342 262226
rect 25398 262170 42970 262226
rect 43026 262170 43094 262226
rect 43150 262170 43218 262226
rect 43274 262170 43342 262226
rect 43398 262170 60970 262226
rect 61026 262170 61094 262226
rect 61150 262170 61218 262226
rect 61274 262170 61342 262226
rect 61398 262170 78970 262226
rect 79026 262170 79094 262226
rect 79150 262170 79218 262226
rect 79274 262170 79342 262226
rect 79398 262170 96970 262226
rect 97026 262170 97094 262226
rect 97150 262170 97218 262226
rect 97274 262170 97342 262226
rect 97398 262170 132970 262226
rect 133026 262170 133094 262226
rect 133150 262170 133218 262226
rect 133274 262170 133342 262226
rect 133398 262170 150970 262226
rect 151026 262170 151094 262226
rect 151150 262170 151218 262226
rect 151274 262170 151342 262226
rect 151398 262170 168970 262226
rect 169026 262170 169094 262226
rect 169150 262170 169218 262226
rect 169274 262170 169342 262226
rect 169398 262170 186970 262226
rect 187026 262170 187094 262226
rect 187150 262170 187218 262226
rect 187274 262170 187342 262226
rect 187398 262170 222970 262226
rect 223026 262170 223094 262226
rect 223150 262170 223218 262226
rect 223274 262170 223342 262226
rect 223398 262170 240970 262226
rect 241026 262170 241094 262226
rect 241150 262170 241218 262226
rect 241274 262170 241342 262226
rect 241398 262170 258970 262226
rect 259026 262170 259094 262226
rect 259150 262170 259218 262226
rect 259274 262170 259342 262226
rect 259398 262170 276970 262226
rect 277026 262170 277094 262226
rect 277150 262170 277218 262226
rect 277274 262170 277342 262226
rect 277398 262170 312970 262226
rect 313026 262170 313094 262226
rect 313150 262170 313218 262226
rect 313274 262170 313342 262226
rect 313398 262170 330970 262226
rect 331026 262170 331094 262226
rect 331150 262170 331218 262226
rect 331274 262170 331342 262226
rect 331398 262170 348970 262226
rect 349026 262170 349094 262226
rect 349150 262170 349218 262226
rect 349274 262170 349342 262226
rect 349398 262170 366970 262226
rect 367026 262170 367094 262226
rect 367150 262170 367218 262226
rect 367274 262170 367342 262226
rect 367398 262170 402970 262226
rect 403026 262170 403094 262226
rect 403150 262170 403218 262226
rect 403274 262170 403342 262226
rect 403398 262170 420970 262226
rect 421026 262170 421094 262226
rect 421150 262170 421218 262226
rect 421274 262170 421342 262226
rect 421398 262170 438970 262226
rect 439026 262170 439094 262226
rect 439150 262170 439218 262226
rect 439274 262170 439342 262226
rect 439398 262170 456970 262226
rect 457026 262170 457094 262226
rect 457150 262170 457218 262226
rect 457274 262170 457342 262226
rect 457398 262170 492970 262226
rect 493026 262170 493094 262226
rect 493150 262170 493218 262226
rect 493274 262170 493342 262226
rect 493398 262170 510970 262226
rect 511026 262170 511094 262226
rect 511150 262170 511218 262226
rect 511274 262170 511342 262226
rect 511398 262170 528970 262226
rect 529026 262170 529094 262226
rect 529150 262170 529218 262226
rect 529274 262170 529342 262226
rect 529398 262170 546970 262226
rect 547026 262170 547094 262226
rect 547150 262170 547218 262226
rect 547274 262170 547342 262226
rect 547398 262170 564970 262226
rect 565026 262170 565094 262226
rect 565150 262170 565218 262226
rect 565274 262170 565342 262226
rect 565398 262170 582970 262226
rect 583026 262170 583094 262226
rect 583150 262170 583218 262226
rect 583274 262170 583342 262226
rect 583398 262170 597456 262226
rect 597512 262170 597580 262226
rect 597636 262170 597704 262226
rect 597760 262170 597828 262226
rect 597884 262170 597980 262226
rect -1916 262102 597980 262170
rect -1916 262046 -1820 262102
rect -1764 262046 -1696 262102
rect -1640 262046 -1572 262102
rect -1516 262046 -1448 262102
rect -1392 262046 6970 262102
rect 7026 262046 7094 262102
rect 7150 262046 7218 262102
rect 7274 262046 7342 262102
rect 7398 262046 24970 262102
rect 25026 262046 25094 262102
rect 25150 262046 25218 262102
rect 25274 262046 25342 262102
rect 25398 262046 42970 262102
rect 43026 262046 43094 262102
rect 43150 262046 43218 262102
rect 43274 262046 43342 262102
rect 43398 262046 60970 262102
rect 61026 262046 61094 262102
rect 61150 262046 61218 262102
rect 61274 262046 61342 262102
rect 61398 262046 78970 262102
rect 79026 262046 79094 262102
rect 79150 262046 79218 262102
rect 79274 262046 79342 262102
rect 79398 262046 96970 262102
rect 97026 262046 97094 262102
rect 97150 262046 97218 262102
rect 97274 262046 97342 262102
rect 97398 262046 132970 262102
rect 133026 262046 133094 262102
rect 133150 262046 133218 262102
rect 133274 262046 133342 262102
rect 133398 262046 150970 262102
rect 151026 262046 151094 262102
rect 151150 262046 151218 262102
rect 151274 262046 151342 262102
rect 151398 262046 168970 262102
rect 169026 262046 169094 262102
rect 169150 262046 169218 262102
rect 169274 262046 169342 262102
rect 169398 262046 186970 262102
rect 187026 262046 187094 262102
rect 187150 262046 187218 262102
rect 187274 262046 187342 262102
rect 187398 262046 222970 262102
rect 223026 262046 223094 262102
rect 223150 262046 223218 262102
rect 223274 262046 223342 262102
rect 223398 262046 240970 262102
rect 241026 262046 241094 262102
rect 241150 262046 241218 262102
rect 241274 262046 241342 262102
rect 241398 262046 258970 262102
rect 259026 262046 259094 262102
rect 259150 262046 259218 262102
rect 259274 262046 259342 262102
rect 259398 262046 276970 262102
rect 277026 262046 277094 262102
rect 277150 262046 277218 262102
rect 277274 262046 277342 262102
rect 277398 262046 312970 262102
rect 313026 262046 313094 262102
rect 313150 262046 313218 262102
rect 313274 262046 313342 262102
rect 313398 262046 330970 262102
rect 331026 262046 331094 262102
rect 331150 262046 331218 262102
rect 331274 262046 331342 262102
rect 331398 262046 348970 262102
rect 349026 262046 349094 262102
rect 349150 262046 349218 262102
rect 349274 262046 349342 262102
rect 349398 262046 366970 262102
rect 367026 262046 367094 262102
rect 367150 262046 367218 262102
rect 367274 262046 367342 262102
rect 367398 262046 402970 262102
rect 403026 262046 403094 262102
rect 403150 262046 403218 262102
rect 403274 262046 403342 262102
rect 403398 262046 420970 262102
rect 421026 262046 421094 262102
rect 421150 262046 421218 262102
rect 421274 262046 421342 262102
rect 421398 262046 438970 262102
rect 439026 262046 439094 262102
rect 439150 262046 439218 262102
rect 439274 262046 439342 262102
rect 439398 262046 456970 262102
rect 457026 262046 457094 262102
rect 457150 262046 457218 262102
rect 457274 262046 457342 262102
rect 457398 262046 492970 262102
rect 493026 262046 493094 262102
rect 493150 262046 493218 262102
rect 493274 262046 493342 262102
rect 493398 262046 510970 262102
rect 511026 262046 511094 262102
rect 511150 262046 511218 262102
rect 511274 262046 511342 262102
rect 511398 262046 528970 262102
rect 529026 262046 529094 262102
rect 529150 262046 529218 262102
rect 529274 262046 529342 262102
rect 529398 262046 546970 262102
rect 547026 262046 547094 262102
rect 547150 262046 547218 262102
rect 547274 262046 547342 262102
rect 547398 262046 564970 262102
rect 565026 262046 565094 262102
rect 565150 262046 565218 262102
rect 565274 262046 565342 262102
rect 565398 262046 582970 262102
rect 583026 262046 583094 262102
rect 583150 262046 583218 262102
rect 583274 262046 583342 262102
rect 583398 262046 597456 262102
rect 597512 262046 597580 262102
rect 597636 262046 597704 262102
rect 597760 262046 597828 262102
rect 597884 262046 597980 262102
rect -1916 261978 597980 262046
rect -1916 261922 -1820 261978
rect -1764 261922 -1696 261978
rect -1640 261922 -1572 261978
rect -1516 261922 -1448 261978
rect -1392 261922 6970 261978
rect 7026 261922 7094 261978
rect 7150 261922 7218 261978
rect 7274 261922 7342 261978
rect 7398 261922 24970 261978
rect 25026 261922 25094 261978
rect 25150 261922 25218 261978
rect 25274 261922 25342 261978
rect 25398 261922 42970 261978
rect 43026 261922 43094 261978
rect 43150 261922 43218 261978
rect 43274 261922 43342 261978
rect 43398 261922 60970 261978
rect 61026 261922 61094 261978
rect 61150 261922 61218 261978
rect 61274 261922 61342 261978
rect 61398 261922 78970 261978
rect 79026 261922 79094 261978
rect 79150 261922 79218 261978
rect 79274 261922 79342 261978
rect 79398 261922 96970 261978
rect 97026 261922 97094 261978
rect 97150 261922 97218 261978
rect 97274 261922 97342 261978
rect 97398 261922 132970 261978
rect 133026 261922 133094 261978
rect 133150 261922 133218 261978
rect 133274 261922 133342 261978
rect 133398 261922 150970 261978
rect 151026 261922 151094 261978
rect 151150 261922 151218 261978
rect 151274 261922 151342 261978
rect 151398 261922 168970 261978
rect 169026 261922 169094 261978
rect 169150 261922 169218 261978
rect 169274 261922 169342 261978
rect 169398 261922 186970 261978
rect 187026 261922 187094 261978
rect 187150 261922 187218 261978
rect 187274 261922 187342 261978
rect 187398 261922 222970 261978
rect 223026 261922 223094 261978
rect 223150 261922 223218 261978
rect 223274 261922 223342 261978
rect 223398 261922 240970 261978
rect 241026 261922 241094 261978
rect 241150 261922 241218 261978
rect 241274 261922 241342 261978
rect 241398 261922 258970 261978
rect 259026 261922 259094 261978
rect 259150 261922 259218 261978
rect 259274 261922 259342 261978
rect 259398 261922 276970 261978
rect 277026 261922 277094 261978
rect 277150 261922 277218 261978
rect 277274 261922 277342 261978
rect 277398 261922 312970 261978
rect 313026 261922 313094 261978
rect 313150 261922 313218 261978
rect 313274 261922 313342 261978
rect 313398 261922 330970 261978
rect 331026 261922 331094 261978
rect 331150 261922 331218 261978
rect 331274 261922 331342 261978
rect 331398 261922 348970 261978
rect 349026 261922 349094 261978
rect 349150 261922 349218 261978
rect 349274 261922 349342 261978
rect 349398 261922 366970 261978
rect 367026 261922 367094 261978
rect 367150 261922 367218 261978
rect 367274 261922 367342 261978
rect 367398 261922 402970 261978
rect 403026 261922 403094 261978
rect 403150 261922 403218 261978
rect 403274 261922 403342 261978
rect 403398 261922 420970 261978
rect 421026 261922 421094 261978
rect 421150 261922 421218 261978
rect 421274 261922 421342 261978
rect 421398 261922 438970 261978
rect 439026 261922 439094 261978
rect 439150 261922 439218 261978
rect 439274 261922 439342 261978
rect 439398 261922 456970 261978
rect 457026 261922 457094 261978
rect 457150 261922 457218 261978
rect 457274 261922 457342 261978
rect 457398 261922 492970 261978
rect 493026 261922 493094 261978
rect 493150 261922 493218 261978
rect 493274 261922 493342 261978
rect 493398 261922 510970 261978
rect 511026 261922 511094 261978
rect 511150 261922 511218 261978
rect 511274 261922 511342 261978
rect 511398 261922 528970 261978
rect 529026 261922 529094 261978
rect 529150 261922 529218 261978
rect 529274 261922 529342 261978
rect 529398 261922 546970 261978
rect 547026 261922 547094 261978
rect 547150 261922 547218 261978
rect 547274 261922 547342 261978
rect 547398 261922 564970 261978
rect 565026 261922 565094 261978
rect 565150 261922 565218 261978
rect 565274 261922 565342 261978
rect 565398 261922 582970 261978
rect 583026 261922 583094 261978
rect 583150 261922 583218 261978
rect 583274 261922 583342 261978
rect 583398 261922 597456 261978
rect 597512 261922 597580 261978
rect 597636 261922 597704 261978
rect 597760 261922 597828 261978
rect 597884 261922 597980 261978
rect -1916 261826 597980 261922
rect -1916 256350 597980 256446
rect -1916 256294 -860 256350
rect -804 256294 -736 256350
rect -680 256294 -612 256350
rect -556 256294 -488 256350
rect -432 256294 3250 256350
rect 3306 256294 3374 256350
rect 3430 256294 3498 256350
rect 3554 256294 3622 256350
rect 3678 256294 21250 256350
rect 21306 256294 21374 256350
rect 21430 256294 21498 256350
rect 21554 256294 21622 256350
rect 21678 256294 39250 256350
rect 39306 256294 39374 256350
rect 39430 256294 39498 256350
rect 39554 256294 39622 256350
rect 39678 256294 57250 256350
rect 57306 256294 57374 256350
rect 57430 256294 57498 256350
rect 57554 256294 57622 256350
rect 57678 256294 93250 256350
rect 93306 256294 93374 256350
rect 93430 256294 93498 256350
rect 93554 256294 93622 256350
rect 93678 256294 111250 256350
rect 111306 256294 111374 256350
rect 111430 256294 111498 256350
rect 111554 256294 111622 256350
rect 111678 256294 129250 256350
rect 129306 256294 129374 256350
rect 129430 256294 129498 256350
rect 129554 256294 129622 256350
rect 129678 256294 147250 256350
rect 147306 256294 147374 256350
rect 147430 256294 147498 256350
rect 147554 256294 147622 256350
rect 147678 256294 183250 256350
rect 183306 256294 183374 256350
rect 183430 256294 183498 256350
rect 183554 256294 183622 256350
rect 183678 256294 201250 256350
rect 201306 256294 201374 256350
rect 201430 256294 201498 256350
rect 201554 256294 201622 256350
rect 201678 256294 219250 256350
rect 219306 256294 219374 256350
rect 219430 256294 219498 256350
rect 219554 256294 219622 256350
rect 219678 256294 237250 256350
rect 237306 256294 237374 256350
rect 237430 256294 237498 256350
rect 237554 256294 237622 256350
rect 237678 256294 273250 256350
rect 273306 256294 273374 256350
rect 273430 256294 273498 256350
rect 273554 256294 273622 256350
rect 273678 256294 291250 256350
rect 291306 256294 291374 256350
rect 291430 256294 291498 256350
rect 291554 256294 291622 256350
rect 291678 256294 309250 256350
rect 309306 256294 309374 256350
rect 309430 256294 309498 256350
rect 309554 256294 309622 256350
rect 309678 256294 327250 256350
rect 327306 256294 327374 256350
rect 327430 256294 327498 256350
rect 327554 256294 327622 256350
rect 327678 256294 363250 256350
rect 363306 256294 363374 256350
rect 363430 256294 363498 256350
rect 363554 256294 363622 256350
rect 363678 256294 381250 256350
rect 381306 256294 381374 256350
rect 381430 256294 381498 256350
rect 381554 256294 381622 256350
rect 381678 256294 399250 256350
rect 399306 256294 399374 256350
rect 399430 256294 399498 256350
rect 399554 256294 399622 256350
rect 399678 256294 417250 256350
rect 417306 256294 417374 256350
rect 417430 256294 417498 256350
rect 417554 256294 417622 256350
rect 417678 256294 453250 256350
rect 453306 256294 453374 256350
rect 453430 256294 453498 256350
rect 453554 256294 453622 256350
rect 453678 256294 471250 256350
rect 471306 256294 471374 256350
rect 471430 256294 471498 256350
rect 471554 256294 471622 256350
rect 471678 256294 489250 256350
rect 489306 256294 489374 256350
rect 489430 256294 489498 256350
rect 489554 256294 489622 256350
rect 489678 256294 507250 256350
rect 507306 256294 507374 256350
rect 507430 256294 507498 256350
rect 507554 256294 507622 256350
rect 507678 256294 543250 256350
rect 543306 256294 543374 256350
rect 543430 256294 543498 256350
rect 543554 256294 543622 256350
rect 543678 256294 561250 256350
rect 561306 256294 561374 256350
rect 561430 256294 561498 256350
rect 561554 256294 561622 256350
rect 561678 256294 579250 256350
rect 579306 256294 579374 256350
rect 579430 256294 579498 256350
rect 579554 256294 579622 256350
rect 579678 256294 596496 256350
rect 596552 256294 596620 256350
rect 596676 256294 596744 256350
rect 596800 256294 596868 256350
rect 596924 256294 597980 256350
rect -1916 256226 597980 256294
rect -1916 256170 -860 256226
rect -804 256170 -736 256226
rect -680 256170 -612 256226
rect -556 256170 -488 256226
rect -432 256170 3250 256226
rect 3306 256170 3374 256226
rect 3430 256170 3498 256226
rect 3554 256170 3622 256226
rect 3678 256170 21250 256226
rect 21306 256170 21374 256226
rect 21430 256170 21498 256226
rect 21554 256170 21622 256226
rect 21678 256170 39250 256226
rect 39306 256170 39374 256226
rect 39430 256170 39498 256226
rect 39554 256170 39622 256226
rect 39678 256170 57250 256226
rect 57306 256170 57374 256226
rect 57430 256170 57498 256226
rect 57554 256170 57622 256226
rect 57678 256170 93250 256226
rect 93306 256170 93374 256226
rect 93430 256170 93498 256226
rect 93554 256170 93622 256226
rect 93678 256170 111250 256226
rect 111306 256170 111374 256226
rect 111430 256170 111498 256226
rect 111554 256170 111622 256226
rect 111678 256170 129250 256226
rect 129306 256170 129374 256226
rect 129430 256170 129498 256226
rect 129554 256170 129622 256226
rect 129678 256170 147250 256226
rect 147306 256170 147374 256226
rect 147430 256170 147498 256226
rect 147554 256170 147622 256226
rect 147678 256170 183250 256226
rect 183306 256170 183374 256226
rect 183430 256170 183498 256226
rect 183554 256170 183622 256226
rect 183678 256170 201250 256226
rect 201306 256170 201374 256226
rect 201430 256170 201498 256226
rect 201554 256170 201622 256226
rect 201678 256170 219250 256226
rect 219306 256170 219374 256226
rect 219430 256170 219498 256226
rect 219554 256170 219622 256226
rect 219678 256170 237250 256226
rect 237306 256170 237374 256226
rect 237430 256170 237498 256226
rect 237554 256170 237622 256226
rect 237678 256170 273250 256226
rect 273306 256170 273374 256226
rect 273430 256170 273498 256226
rect 273554 256170 273622 256226
rect 273678 256170 291250 256226
rect 291306 256170 291374 256226
rect 291430 256170 291498 256226
rect 291554 256170 291622 256226
rect 291678 256170 309250 256226
rect 309306 256170 309374 256226
rect 309430 256170 309498 256226
rect 309554 256170 309622 256226
rect 309678 256170 327250 256226
rect 327306 256170 327374 256226
rect 327430 256170 327498 256226
rect 327554 256170 327622 256226
rect 327678 256170 363250 256226
rect 363306 256170 363374 256226
rect 363430 256170 363498 256226
rect 363554 256170 363622 256226
rect 363678 256170 381250 256226
rect 381306 256170 381374 256226
rect 381430 256170 381498 256226
rect 381554 256170 381622 256226
rect 381678 256170 399250 256226
rect 399306 256170 399374 256226
rect 399430 256170 399498 256226
rect 399554 256170 399622 256226
rect 399678 256170 417250 256226
rect 417306 256170 417374 256226
rect 417430 256170 417498 256226
rect 417554 256170 417622 256226
rect 417678 256170 453250 256226
rect 453306 256170 453374 256226
rect 453430 256170 453498 256226
rect 453554 256170 453622 256226
rect 453678 256170 471250 256226
rect 471306 256170 471374 256226
rect 471430 256170 471498 256226
rect 471554 256170 471622 256226
rect 471678 256170 489250 256226
rect 489306 256170 489374 256226
rect 489430 256170 489498 256226
rect 489554 256170 489622 256226
rect 489678 256170 507250 256226
rect 507306 256170 507374 256226
rect 507430 256170 507498 256226
rect 507554 256170 507622 256226
rect 507678 256170 543250 256226
rect 543306 256170 543374 256226
rect 543430 256170 543498 256226
rect 543554 256170 543622 256226
rect 543678 256170 561250 256226
rect 561306 256170 561374 256226
rect 561430 256170 561498 256226
rect 561554 256170 561622 256226
rect 561678 256170 579250 256226
rect 579306 256170 579374 256226
rect 579430 256170 579498 256226
rect 579554 256170 579622 256226
rect 579678 256170 596496 256226
rect 596552 256170 596620 256226
rect 596676 256170 596744 256226
rect 596800 256170 596868 256226
rect 596924 256170 597980 256226
rect -1916 256102 597980 256170
rect -1916 256046 -860 256102
rect -804 256046 -736 256102
rect -680 256046 -612 256102
rect -556 256046 -488 256102
rect -432 256046 3250 256102
rect 3306 256046 3374 256102
rect 3430 256046 3498 256102
rect 3554 256046 3622 256102
rect 3678 256046 21250 256102
rect 21306 256046 21374 256102
rect 21430 256046 21498 256102
rect 21554 256046 21622 256102
rect 21678 256046 39250 256102
rect 39306 256046 39374 256102
rect 39430 256046 39498 256102
rect 39554 256046 39622 256102
rect 39678 256046 57250 256102
rect 57306 256046 57374 256102
rect 57430 256046 57498 256102
rect 57554 256046 57622 256102
rect 57678 256046 93250 256102
rect 93306 256046 93374 256102
rect 93430 256046 93498 256102
rect 93554 256046 93622 256102
rect 93678 256046 111250 256102
rect 111306 256046 111374 256102
rect 111430 256046 111498 256102
rect 111554 256046 111622 256102
rect 111678 256046 129250 256102
rect 129306 256046 129374 256102
rect 129430 256046 129498 256102
rect 129554 256046 129622 256102
rect 129678 256046 147250 256102
rect 147306 256046 147374 256102
rect 147430 256046 147498 256102
rect 147554 256046 147622 256102
rect 147678 256046 183250 256102
rect 183306 256046 183374 256102
rect 183430 256046 183498 256102
rect 183554 256046 183622 256102
rect 183678 256046 201250 256102
rect 201306 256046 201374 256102
rect 201430 256046 201498 256102
rect 201554 256046 201622 256102
rect 201678 256046 219250 256102
rect 219306 256046 219374 256102
rect 219430 256046 219498 256102
rect 219554 256046 219622 256102
rect 219678 256046 237250 256102
rect 237306 256046 237374 256102
rect 237430 256046 237498 256102
rect 237554 256046 237622 256102
rect 237678 256046 273250 256102
rect 273306 256046 273374 256102
rect 273430 256046 273498 256102
rect 273554 256046 273622 256102
rect 273678 256046 291250 256102
rect 291306 256046 291374 256102
rect 291430 256046 291498 256102
rect 291554 256046 291622 256102
rect 291678 256046 309250 256102
rect 309306 256046 309374 256102
rect 309430 256046 309498 256102
rect 309554 256046 309622 256102
rect 309678 256046 327250 256102
rect 327306 256046 327374 256102
rect 327430 256046 327498 256102
rect 327554 256046 327622 256102
rect 327678 256046 363250 256102
rect 363306 256046 363374 256102
rect 363430 256046 363498 256102
rect 363554 256046 363622 256102
rect 363678 256046 381250 256102
rect 381306 256046 381374 256102
rect 381430 256046 381498 256102
rect 381554 256046 381622 256102
rect 381678 256046 399250 256102
rect 399306 256046 399374 256102
rect 399430 256046 399498 256102
rect 399554 256046 399622 256102
rect 399678 256046 417250 256102
rect 417306 256046 417374 256102
rect 417430 256046 417498 256102
rect 417554 256046 417622 256102
rect 417678 256046 453250 256102
rect 453306 256046 453374 256102
rect 453430 256046 453498 256102
rect 453554 256046 453622 256102
rect 453678 256046 471250 256102
rect 471306 256046 471374 256102
rect 471430 256046 471498 256102
rect 471554 256046 471622 256102
rect 471678 256046 489250 256102
rect 489306 256046 489374 256102
rect 489430 256046 489498 256102
rect 489554 256046 489622 256102
rect 489678 256046 507250 256102
rect 507306 256046 507374 256102
rect 507430 256046 507498 256102
rect 507554 256046 507622 256102
rect 507678 256046 543250 256102
rect 543306 256046 543374 256102
rect 543430 256046 543498 256102
rect 543554 256046 543622 256102
rect 543678 256046 561250 256102
rect 561306 256046 561374 256102
rect 561430 256046 561498 256102
rect 561554 256046 561622 256102
rect 561678 256046 579250 256102
rect 579306 256046 579374 256102
rect 579430 256046 579498 256102
rect 579554 256046 579622 256102
rect 579678 256046 596496 256102
rect 596552 256046 596620 256102
rect 596676 256046 596744 256102
rect 596800 256046 596868 256102
rect 596924 256046 597980 256102
rect -1916 255978 597980 256046
rect -1916 255922 -860 255978
rect -804 255922 -736 255978
rect -680 255922 -612 255978
rect -556 255922 -488 255978
rect -432 255922 3250 255978
rect 3306 255922 3374 255978
rect 3430 255922 3498 255978
rect 3554 255922 3622 255978
rect 3678 255922 21250 255978
rect 21306 255922 21374 255978
rect 21430 255922 21498 255978
rect 21554 255922 21622 255978
rect 21678 255922 39250 255978
rect 39306 255922 39374 255978
rect 39430 255922 39498 255978
rect 39554 255922 39622 255978
rect 39678 255922 57250 255978
rect 57306 255922 57374 255978
rect 57430 255922 57498 255978
rect 57554 255922 57622 255978
rect 57678 255922 93250 255978
rect 93306 255922 93374 255978
rect 93430 255922 93498 255978
rect 93554 255922 93622 255978
rect 93678 255922 111250 255978
rect 111306 255922 111374 255978
rect 111430 255922 111498 255978
rect 111554 255922 111622 255978
rect 111678 255922 129250 255978
rect 129306 255922 129374 255978
rect 129430 255922 129498 255978
rect 129554 255922 129622 255978
rect 129678 255922 147250 255978
rect 147306 255922 147374 255978
rect 147430 255922 147498 255978
rect 147554 255922 147622 255978
rect 147678 255922 183250 255978
rect 183306 255922 183374 255978
rect 183430 255922 183498 255978
rect 183554 255922 183622 255978
rect 183678 255922 201250 255978
rect 201306 255922 201374 255978
rect 201430 255922 201498 255978
rect 201554 255922 201622 255978
rect 201678 255922 219250 255978
rect 219306 255922 219374 255978
rect 219430 255922 219498 255978
rect 219554 255922 219622 255978
rect 219678 255922 237250 255978
rect 237306 255922 237374 255978
rect 237430 255922 237498 255978
rect 237554 255922 237622 255978
rect 237678 255922 273250 255978
rect 273306 255922 273374 255978
rect 273430 255922 273498 255978
rect 273554 255922 273622 255978
rect 273678 255922 291250 255978
rect 291306 255922 291374 255978
rect 291430 255922 291498 255978
rect 291554 255922 291622 255978
rect 291678 255922 309250 255978
rect 309306 255922 309374 255978
rect 309430 255922 309498 255978
rect 309554 255922 309622 255978
rect 309678 255922 327250 255978
rect 327306 255922 327374 255978
rect 327430 255922 327498 255978
rect 327554 255922 327622 255978
rect 327678 255922 363250 255978
rect 363306 255922 363374 255978
rect 363430 255922 363498 255978
rect 363554 255922 363622 255978
rect 363678 255922 381250 255978
rect 381306 255922 381374 255978
rect 381430 255922 381498 255978
rect 381554 255922 381622 255978
rect 381678 255922 399250 255978
rect 399306 255922 399374 255978
rect 399430 255922 399498 255978
rect 399554 255922 399622 255978
rect 399678 255922 417250 255978
rect 417306 255922 417374 255978
rect 417430 255922 417498 255978
rect 417554 255922 417622 255978
rect 417678 255922 453250 255978
rect 453306 255922 453374 255978
rect 453430 255922 453498 255978
rect 453554 255922 453622 255978
rect 453678 255922 471250 255978
rect 471306 255922 471374 255978
rect 471430 255922 471498 255978
rect 471554 255922 471622 255978
rect 471678 255922 489250 255978
rect 489306 255922 489374 255978
rect 489430 255922 489498 255978
rect 489554 255922 489622 255978
rect 489678 255922 507250 255978
rect 507306 255922 507374 255978
rect 507430 255922 507498 255978
rect 507554 255922 507622 255978
rect 507678 255922 543250 255978
rect 543306 255922 543374 255978
rect 543430 255922 543498 255978
rect 543554 255922 543622 255978
rect 543678 255922 561250 255978
rect 561306 255922 561374 255978
rect 561430 255922 561498 255978
rect 561554 255922 561622 255978
rect 561678 255922 579250 255978
rect 579306 255922 579374 255978
rect 579430 255922 579498 255978
rect 579554 255922 579622 255978
rect 579678 255922 596496 255978
rect 596552 255922 596620 255978
rect 596676 255922 596744 255978
rect 596800 255922 596868 255978
rect 596924 255922 597980 255978
rect -1916 255826 597980 255922
rect -1916 244350 597980 244446
rect -1916 244294 -1820 244350
rect -1764 244294 -1696 244350
rect -1640 244294 -1572 244350
rect -1516 244294 -1448 244350
rect -1392 244294 6970 244350
rect 7026 244294 7094 244350
rect 7150 244294 7218 244350
rect 7274 244294 7342 244350
rect 7398 244294 24970 244350
rect 25026 244294 25094 244350
rect 25150 244294 25218 244350
rect 25274 244294 25342 244350
rect 25398 244294 42970 244350
rect 43026 244294 43094 244350
rect 43150 244294 43218 244350
rect 43274 244294 43342 244350
rect 43398 244294 60970 244350
rect 61026 244294 61094 244350
rect 61150 244294 61218 244350
rect 61274 244294 61342 244350
rect 61398 244294 78970 244350
rect 79026 244294 79094 244350
rect 79150 244294 79218 244350
rect 79274 244294 79342 244350
rect 79398 244294 96970 244350
rect 97026 244294 97094 244350
rect 97150 244294 97218 244350
rect 97274 244294 97342 244350
rect 97398 244294 132970 244350
rect 133026 244294 133094 244350
rect 133150 244294 133218 244350
rect 133274 244294 133342 244350
rect 133398 244294 150970 244350
rect 151026 244294 151094 244350
rect 151150 244294 151218 244350
rect 151274 244294 151342 244350
rect 151398 244294 168970 244350
rect 169026 244294 169094 244350
rect 169150 244294 169218 244350
rect 169274 244294 169342 244350
rect 169398 244294 186970 244350
rect 187026 244294 187094 244350
rect 187150 244294 187218 244350
rect 187274 244294 187342 244350
rect 187398 244294 222970 244350
rect 223026 244294 223094 244350
rect 223150 244294 223218 244350
rect 223274 244294 223342 244350
rect 223398 244294 240970 244350
rect 241026 244294 241094 244350
rect 241150 244294 241218 244350
rect 241274 244294 241342 244350
rect 241398 244294 258970 244350
rect 259026 244294 259094 244350
rect 259150 244294 259218 244350
rect 259274 244294 259342 244350
rect 259398 244294 276970 244350
rect 277026 244294 277094 244350
rect 277150 244294 277218 244350
rect 277274 244294 277342 244350
rect 277398 244294 312970 244350
rect 313026 244294 313094 244350
rect 313150 244294 313218 244350
rect 313274 244294 313342 244350
rect 313398 244294 330970 244350
rect 331026 244294 331094 244350
rect 331150 244294 331218 244350
rect 331274 244294 331342 244350
rect 331398 244294 348970 244350
rect 349026 244294 349094 244350
rect 349150 244294 349218 244350
rect 349274 244294 349342 244350
rect 349398 244294 366970 244350
rect 367026 244294 367094 244350
rect 367150 244294 367218 244350
rect 367274 244294 367342 244350
rect 367398 244294 402970 244350
rect 403026 244294 403094 244350
rect 403150 244294 403218 244350
rect 403274 244294 403342 244350
rect 403398 244294 420970 244350
rect 421026 244294 421094 244350
rect 421150 244294 421218 244350
rect 421274 244294 421342 244350
rect 421398 244294 438970 244350
rect 439026 244294 439094 244350
rect 439150 244294 439218 244350
rect 439274 244294 439342 244350
rect 439398 244294 456970 244350
rect 457026 244294 457094 244350
rect 457150 244294 457218 244350
rect 457274 244294 457342 244350
rect 457398 244294 492970 244350
rect 493026 244294 493094 244350
rect 493150 244294 493218 244350
rect 493274 244294 493342 244350
rect 493398 244294 510970 244350
rect 511026 244294 511094 244350
rect 511150 244294 511218 244350
rect 511274 244294 511342 244350
rect 511398 244294 528970 244350
rect 529026 244294 529094 244350
rect 529150 244294 529218 244350
rect 529274 244294 529342 244350
rect 529398 244294 546970 244350
rect 547026 244294 547094 244350
rect 547150 244294 547218 244350
rect 547274 244294 547342 244350
rect 547398 244294 564970 244350
rect 565026 244294 565094 244350
rect 565150 244294 565218 244350
rect 565274 244294 565342 244350
rect 565398 244294 582970 244350
rect 583026 244294 583094 244350
rect 583150 244294 583218 244350
rect 583274 244294 583342 244350
rect 583398 244294 597456 244350
rect 597512 244294 597580 244350
rect 597636 244294 597704 244350
rect 597760 244294 597828 244350
rect 597884 244294 597980 244350
rect -1916 244226 597980 244294
rect -1916 244170 -1820 244226
rect -1764 244170 -1696 244226
rect -1640 244170 -1572 244226
rect -1516 244170 -1448 244226
rect -1392 244170 6970 244226
rect 7026 244170 7094 244226
rect 7150 244170 7218 244226
rect 7274 244170 7342 244226
rect 7398 244170 24970 244226
rect 25026 244170 25094 244226
rect 25150 244170 25218 244226
rect 25274 244170 25342 244226
rect 25398 244170 42970 244226
rect 43026 244170 43094 244226
rect 43150 244170 43218 244226
rect 43274 244170 43342 244226
rect 43398 244170 60970 244226
rect 61026 244170 61094 244226
rect 61150 244170 61218 244226
rect 61274 244170 61342 244226
rect 61398 244170 78970 244226
rect 79026 244170 79094 244226
rect 79150 244170 79218 244226
rect 79274 244170 79342 244226
rect 79398 244170 96970 244226
rect 97026 244170 97094 244226
rect 97150 244170 97218 244226
rect 97274 244170 97342 244226
rect 97398 244170 132970 244226
rect 133026 244170 133094 244226
rect 133150 244170 133218 244226
rect 133274 244170 133342 244226
rect 133398 244170 150970 244226
rect 151026 244170 151094 244226
rect 151150 244170 151218 244226
rect 151274 244170 151342 244226
rect 151398 244170 168970 244226
rect 169026 244170 169094 244226
rect 169150 244170 169218 244226
rect 169274 244170 169342 244226
rect 169398 244170 186970 244226
rect 187026 244170 187094 244226
rect 187150 244170 187218 244226
rect 187274 244170 187342 244226
rect 187398 244170 222970 244226
rect 223026 244170 223094 244226
rect 223150 244170 223218 244226
rect 223274 244170 223342 244226
rect 223398 244170 240970 244226
rect 241026 244170 241094 244226
rect 241150 244170 241218 244226
rect 241274 244170 241342 244226
rect 241398 244170 258970 244226
rect 259026 244170 259094 244226
rect 259150 244170 259218 244226
rect 259274 244170 259342 244226
rect 259398 244170 276970 244226
rect 277026 244170 277094 244226
rect 277150 244170 277218 244226
rect 277274 244170 277342 244226
rect 277398 244170 312970 244226
rect 313026 244170 313094 244226
rect 313150 244170 313218 244226
rect 313274 244170 313342 244226
rect 313398 244170 330970 244226
rect 331026 244170 331094 244226
rect 331150 244170 331218 244226
rect 331274 244170 331342 244226
rect 331398 244170 348970 244226
rect 349026 244170 349094 244226
rect 349150 244170 349218 244226
rect 349274 244170 349342 244226
rect 349398 244170 366970 244226
rect 367026 244170 367094 244226
rect 367150 244170 367218 244226
rect 367274 244170 367342 244226
rect 367398 244170 402970 244226
rect 403026 244170 403094 244226
rect 403150 244170 403218 244226
rect 403274 244170 403342 244226
rect 403398 244170 420970 244226
rect 421026 244170 421094 244226
rect 421150 244170 421218 244226
rect 421274 244170 421342 244226
rect 421398 244170 438970 244226
rect 439026 244170 439094 244226
rect 439150 244170 439218 244226
rect 439274 244170 439342 244226
rect 439398 244170 456970 244226
rect 457026 244170 457094 244226
rect 457150 244170 457218 244226
rect 457274 244170 457342 244226
rect 457398 244170 492970 244226
rect 493026 244170 493094 244226
rect 493150 244170 493218 244226
rect 493274 244170 493342 244226
rect 493398 244170 510970 244226
rect 511026 244170 511094 244226
rect 511150 244170 511218 244226
rect 511274 244170 511342 244226
rect 511398 244170 528970 244226
rect 529026 244170 529094 244226
rect 529150 244170 529218 244226
rect 529274 244170 529342 244226
rect 529398 244170 546970 244226
rect 547026 244170 547094 244226
rect 547150 244170 547218 244226
rect 547274 244170 547342 244226
rect 547398 244170 564970 244226
rect 565026 244170 565094 244226
rect 565150 244170 565218 244226
rect 565274 244170 565342 244226
rect 565398 244170 582970 244226
rect 583026 244170 583094 244226
rect 583150 244170 583218 244226
rect 583274 244170 583342 244226
rect 583398 244170 597456 244226
rect 597512 244170 597580 244226
rect 597636 244170 597704 244226
rect 597760 244170 597828 244226
rect 597884 244170 597980 244226
rect -1916 244102 597980 244170
rect -1916 244046 -1820 244102
rect -1764 244046 -1696 244102
rect -1640 244046 -1572 244102
rect -1516 244046 -1448 244102
rect -1392 244046 6970 244102
rect 7026 244046 7094 244102
rect 7150 244046 7218 244102
rect 7274 244046 7342 244102
rect 7398 244046 24970 244102
rect 25026 244046 25094 244102
rect 25150 244046 25218 244102
rect 25274 244046 25342 244102
rect 25398 244046 42970 244102
rect 43026 244046 43094 244102
rect 43150 244046 43218 244102
rect 43274 244046 43342 244102
rect 43398 244046 60970 244102
rect 61026 244046 61094 244102
rect 61150 244046 61218 244102
rect 61274 244046 61342 244102
rect 61398 244046 78970 244102
rect 79026 244046 79094 244102
rect 79150 244046 79218 244102
rect 79274 244046 79342 244102
rect 79398 244046 96970 244102
rect 97026 244046 97094 244102
rect 97150 244046 97218 244102
rect 97274 244046 97342 244102
rect 97398 244046 132970 244102
rect 133026 244046 133094 244102
rect 133150 244046 133218 244102
rect 133274 244046 133342 244102
rect 133398 244046 150970 244102
rect 151026 244046 151094 244102
rect 151150 244046 151218 244102
rect 151274 244046 151342 244102
rect 151398 244046 168970 244102
rect 169026 244046 169094 244102
rect 169150 244046 169218 244102
rect 169274 244046 169342 244102
rect 169398 244046 186970 244102
rect 187026 244046 187094 244102
rect 187150 244046 187218 244102
rect 187274 244046 187342 244102
rect 187398 244046 222970 244102
rect 223026 244046 223094 244102
rect 223150 244046 223218 244102
rect 223274 244046 223342 244102
rect 223398 244046 240970 244102
rect 241026 244046 241094 244102
rect 241150 244046 241218 244102
rect 241274 244046 241342 244102
rect 241398 244046 258970 244102
rect 259026 244046 259094 244102
rect 259150 244046 259218 244102
rect 259274 244046 259342 244102
rect 259398 244046 276970 244102
rect 277026 244046 277094 244102
rect 277150 244046 277218 244102
rect 277274 244046 277342 244102
rect 277398 244046 312970 244102
rect 313026 244046 313094 244102
rect 313150 244046 313218 244102
rect 313274 244046 313342 244102
rect 313398 244046 330970 244102
rect 331026 244046 331094 244102
rect 331150 244046 331218 244102
rect 331274 244046 331342 244102
rect 331398 244046 348970 244102
rect 349026 244046 349094 244102
rect 349150 244046 349218 244102
rect 349274 244046 349342 244102
rect 349398 244046 366970 244102
rect 367026 244046 367094 244102
rect 367150 244046 367218 244102
rect 367274 244046 367342 244102
rect 367398 244046 402970 244102
rect 403026 244046 403094 244102
rect 403150 244046 403218 244102
rect 403274 244046 403342 244102
rect 403398 244046 420970 244102
rect 421026 244046 421094 244102
rect 421150 244046 421218 244102
rect 421274 244046 421342 244102
rect 421398 244046 438970 244102
rect 439026 244046 439094 244102
rect 439150 244046 439218 244102
rect 439274 244046 439342 244102
rect 439398 244046 456970 244102
rect 457026 244046 457094 244102
rect 457150 244046 457218 244102
rect 457274 244046 457342 244102
rect 457398 244046 492970 244102
rect 493026 244046 493094 244102
rect 493150 244046 493218 244102
rect 493274 244046 493342 244102
rect 493398 244046 510970 244102
rect 511026 244046 511094 244102
rect 511150 244046 511218 244102
rect 511274 244046 511342 244102
rect 511398 244046 528970 244102
rect 529026 244046 529094 244102
rect 529150 244046 529218 244102
rect 529274 244046 529342 244102
rect 529398 244046 546970 244102
rect 547026 244046 547094 244102
rect 547150 244046 547218 244102
rect 547274 244046 547342 244102
rect 547398 244046 564970 244102
rect 565026 244046 565094 244102
rect 565150 244046 565218 244102
rect 565274 244046 565342 244102
rect 565398 244046 582970 244102
rect 583026 244046 583094 244102
rect 583150 244046 583218 244102
rect 583274 244046 583342 244102
rect 583398 244046 597456 244102
rect 597512 244046 597580 244102
rect 597636 244046 597704 244102
rect 597760 244046 597828 244102
rect 597884 244046 597980 244102
rect -1916 243978 597980 244046
rect -1916 243922 -1820 243978
rect -1764 243922 -1696 243978
rect -1640 243922 -1572 243978
rect -1516 243922 -1448 243978
rect -1392 243922 6970 243978
rect 7026 243922 7094 243978
rect 7150 243922 7218 243978
rect 7274 243922 7342 243978
rect 7398 243922 24970 243978
rect 25026 243922 25094 243978
rect 25150 243922 25218 243978
rect 25274 243922 25342 243978
rect 25398 243922 42970 243978
rect 43026 243922 43094 243978
rect 43150 243922 43218 243978
rect 43274 243922 43342 243978
rect 43398 243922 60970 243978
rect 61026 243922 61094 243978
rect 61150 243922 61218 243978
rect 61274 243922 61342 243978
rect 61398 243922 78970 243978
rect 79026 243922 79094 243978
rect 79150 243922 79218 243978
rect 79274 243922 79342 243978
rect 79398 243922 96970 243978
rect 97026 243922 97094 243978
rect 97150 243922 97218 243978
rect 97274 243922 97342 243978
rect 97398 243922 132970 243978
rect 133026 243922 133094 243978
rect 133150 243922 133218 243978
rect 133274 243922 133342 243978
rect 133398 243922 150970 243978
rect 151026 243922 151094 243978
rect 151150 243922 151218 243978
rect 151274 243922 151342 243978
rect 151398 243922 168970 243978
rect 169026 243922 169094 243978
rect 169150 243922 169218 243978
rect 169274 243922 169342 243978
rect 169398 243922 186970 243978
rect 187026 243922 187094 243978
rect 187150 243922 187218 243978
rect 187274 243922 187342 243978
rect 187398 243922 222970 243978
rect 223026 243922 223094 243978
rect 223150 243922 223218 243978
rect 223274 243922 223342 243978
rect 223398 243922 240970 243978
rect 241026 243922 241094 243978
rect 241150 243922 241218 243978
rect 241274 243922 241342 243978
rect 241398 243922 258970 243978
rect 259026 243922 259094 243978
rect 259150 243922 259218 243978
rect 259274 243922 259342 243978
rect 259398 243922 276970 243978
rect 277026 243922 277094 243978
rect 277150 243922 277218 243978
rect 277274 243922 277342 243978
rect 277398 243922 312970 243978
rect 313026 243922 313094 243978
rect 313150 243922 313218 243978
rect 313274 243922 313342 243978
rect 313398 243922 330970 243978
rect 331026 243922 331094 243978
rect 331150 243922 331218 243978
rect 331274 243922 331342 243978
rect 331398 243922 348970 243978
rect 349026 243922 349094 243978
rect 349150 243922 349218 243978
rect 349274 243922 349342 243978
rect 349398 243922 366970 243978
rect 367026 243922 367094 243978
rect 367150 243922 367218 243978
rect 367274 243922 367342 243978
rect 367398 243922 402970 243978
rect 403026 243922 403094 243978
rect 403150 243922 403218 243978
rect 403274 243922 403342 243978
rect 403398 243922 420970 243978
rect 421026 243922 421094 243978
rect 421150 243922 421218 243978
rect 421274 243922 421342 243978
rect 421398 243922 438970 243978
rect 439026 243922 439094 243978
rect 439150 243922 439218 243978
rect 439274 243922 439342 243978
rect 439398 243922 456970 243978
rect 457026 243922 457094 243978
rect 457150 243922 457218 243978
rect 457274 243922 457342 243978
rect 457398 243922 492970 243978
rect 493026 243922 493094 243978
rect 493150 243922 493218 243978
rect 493274 243922 493342 243978
rect 493398 243922 510970 243978
rect 511026 243922 511094 243978
rect 511150 243922 511218 243978
rect 511274 243922 511342 243978
rect 511398 243922 528970 243978
rect 529026 243922 529094 243978
rect 529150 243922 529218 243978
rect 529274 243922 529342 243978
rect 529398 243922 546970 243978
rect 547026 243922 547094 243978
rect 547150 243922 547218 243978
rect 547274 243922 547342 243978
rect 547398 243922 564970 243978
rect 565026 243922 565094 243978
rect 565150 243922 565218 243978
rect 565274 243922 565342 243978
rect 565398 243922 582970 243978
rect 583026 243922 583094 243978
rect 583150 243922 583218 243978
rect 583274 243922 583342 243978
rect 583398 243922 597456 243978
rect 597512 243922 597580 243978
rect 597636 243922 597704 243978
rect 597760 243922 597828 243978
rect 597884 243922 597980 243978
rect -1916 243826 597980 243922
rect -1916 238350 597980 238446
rect -1916 238294 -860 238350
rect -804 238294 -736 238350
rect -680 238294 -612 238350
rect -556 238294 -488 238350
rect -432 238294 3250 238350
rect 3306 238294 3374 238350
rect 3430 238294 3498 238350
rect 3554 238294 3622 238350
rect 3678 238294 21250 238350
rect 21306 238294 21374 238350
rect 21430 238294 21498 238350
rect 21554 238294 21622 238350
rect 21678 238294 39250 238350
rect 39306 238294 39374 238350
rect 39430 238294 39498 238350
rect 39554 238294 39622 238350
rect 39678 238294 57250 238350
rect 57306 238294 57374 238350
rect 57430 238294 57498 238350
rect 57554 238294 57622 238350
rect 57678 238294 75250 238350
rect 75306 238294 75374 238350
rect 75430 238294 75498 238350
rect 75554 238294 75622 238350
rect 75678 238294 93250 238350
rect 93306 238294 93374 238350
rect 93430 238294 93498 238350
rect 93554 238294 93622 238350
rect 93678 238294 111250 238350
rect 111306 238294 111374 238350
rect 111430 238294 111498 238350
rect 111554 238294 111622 238350
rect 111678 238294 129250 238350
rect 129306 238294 129374 238350
rect 129430 238294 129498 238350
rect 129554 238294 129622 238350
rect 129678 238294 147250 238350
rect 147306 238294 147374 238350
rect 147430 238294 147498 238350
rect 147554 238294 147622 238350
rect 147678 238294 165250 238350
rect 165306 238294 165374 238350
rect 165430 238294 165498 238350
rect 165554 238294 165622 238350
rect 165678 238294 183250 238350
rect 183306 238294 183374 238350
rect 183430 238294 183498 238350
rect 183554 238294 183622 238350
rect 183678 238294 201250 238350
rect 201306 238294 201374 238350
rect 201430 238294 201498 238350
rect 201554 238294 201622 238350
rect 201678 238294 219250 238350
rect 219306 238294 219374 238350
rect 219430 238294 219498 238350
rect 219554 238294 219622 238350
rect 219678 238294 237250 238350
rect 237306 238294 237374 238350
rect 237430 238294 237498 238350
rect 237554 238294 237622 238350
rect 237678 238294 255250 238350
rect 255306 238294 255374 238350
rect 255430 238294 255498 238350
rect 255554 238294 255622 238350
rect 255678 238294 273250 238350
rect 273306 238294 273374 238350
rect 273430 238294 273498 238350
rect 273554 238294 273622 238350
rect 273678 238294 291250 238350
rect 291306 238294 291374 238350
rect 291430 238294 291498 238350
rect 291554 238294 291622 238350
rect 291678 238294 309250 238350
rect 309306 238294 309374 238350
rect 309430 238294 309498 238350
rect 309554 238294 309622 238350
rect 309678 238294 327250 238350
rect 327306 238294 327374 238350
rect 327430 238294 327498 238350
rect 327554 238294 327622 238350
rect 327678 238294 345250 238350
rect 345306 238294 345374 238350
rect 345430 238294 345498 238350
rect 345554 238294 345622 238350
rect 345678 238294 363250 238350
rect 363306 238294 363374 238350
rect 363430 238294 363498 238350
rect 363554 238294 363622 238350
rect 363678 238294 381250 238350
rect 381306 238294 381374 238350
rect 381430 238294 381498 238350
rect 381554 238294 381622 238350
rect 381678 238294 399250 238350
rect 399306 238294 399374 238350
rect 399430 238294 399498 238350
rect 399554 238294 399622 238350
rect 399678 238294 417250 238350
rect 417306 238294 417374 238350
rect 417430 238294 417498 238350
rect 417554 238294 417622 238350
rect 417678 238294 435250 238350
rect 435306 238294 435374 238350
rect 435430 238294 435498 238350
rect 435554 238294 435622 238350
rect 435678 238294 453250 238350
rect 453306 238294 453374 238350
rect 453430 238294 453498 238350
rect 453554 238294 453622 238350
rect 453678 238294 471250 238350
rect 471306 238294 471374 238350
rect 471430 238294 471498 238350
rect 471554 238294 471622 238350
rect 471678 238294 489250 238350
rect 489306 238294 489374 238350
rect 489430 238294 489498 238350
rect 489554 238294 489622 238350
rect 489678 238294 507250 238350
rect 507306 238294 507374 238350
rect 507430 238294 507498 238350
rect 507554 238294 507622 238350
rect 507678 238294 525250 238350
rect 525306 238294 525374 238350
rect 525430 238294 525498 238350
rect 525554 238294 525622 238350
rect 525678 238294 543250 238350
rect 543306 238294 543374 238350
rect 543430 238294 543498 238350
rect 543554 238294 543622 238350
rect 543678 238294 561250 238350
rect 561306 238294 561374 238350
rect 561430 238294 561498 238350
rect 561554 238294 561622 238350
rect 561678 238294 579250 238350
rect 579306 238294 579374 238350
rect 579430 238294 579498 238350
rect 579554 238294 579622 238350
rect 579678 238294 596496 238350
rect 596552 238294 596620 238350
rect 596676 238294 596744 238350
rect 596800 238294 596868 238350
rect 596924 238294 597980 238350
rect -1916 238226 597980 238294
rect -1916 238170 -860 238226
rect -804 238170 -736 238226
rect -680 238170 -612 238226
rect -556 238170 -488 238226
rect -432 238170 3250 238226
rect 3306 238170 3374 238226
rect 3430 238170 3498 238226
rect 3554 238170 3622 238226
rect 3678 238170 21250 238226
rect 21306 238170 21374 238226
rect 21430 238170 21498 238226
rect 21554 238170 21622 238226
rect 21678 238170 39250 238226
rect 39306 238170 39374 238226
rect 39430 238170 39498 238226
rect 39554 238170 39622 238226
rect 39678 238170 57250 238226
rect 57306 238170 57374 238226
rect 57430 238170 57498 238226
rect 57554 238170 57622 238226
rect 57678 238170 75250 238226
rect 75306 238170 75374 238226
rect 75430 238170 75498 238226
rect 75554 238170 75622 238226
rect 75678 238170 93250 238226
rect 93306 238170 93374 238226
rect 93430 238170 93498 238226
rect 93554 238170 93622 238226
rect 93678 238170 111250 238226
rect 111306 238170 111374 238226
rect 111430 238170 111498 238226
rect 111554 238170 111622 238226
rect 111678 238170 129250 238226
rect 129306 238170 129374 238226
rect 129430 238170 129498 238226
rect 129554 238170 129622 238226
rect 129678 238170 147250 238226
rect 147306 238170 147374 238226
rect 147430 238170 147498 238226
rect 147554 238170 147622 238226
rect 147678 238170 165250 238226
rect 165306 238170 165374 238226
rect 165430 238170 165498 238226
rect 165554 238170 165622 238226
rect 165678 238170 183250 238226
rect 183306 238170 183374 238226
rect 183430 238170 183498 238226
rect 183554 238170 183622 238226
rect 183678 238170 201250 238226
rect 201306 238170 201374 238226
rect 201430 238170 201498 238226
rect 201554 238170 201622 238226
rect 201678 238170 219250 238226
rect 219306 238170 219374 238226
rect 219430 238170 219498 238226
rect 219554 238170 219622 238226
rect 219678 238170 237250 238226
rect 237306 238170 237374 238226
rect 237430 238170 237498 238226
rect 237554 238170 237622 238226
rect 237678 238170 255250 238226
rect 255306 238170 255374 238226
rect 255430 238170 255498 238226
rect 255554 238170 255622 238226
rect 255678 238170 273250 238226
rect 273306 238170 273374 238226
rect 273430 238170 273498 238226
rect 273554 238170 273622 238226
rect 273678 238170 291250 238226
rect 291306 238170 291374 238226
rect 291430 238170 291498 238226
rect 291554 238170 291622 238226
rect 291678 238170 309250 238226
rect 309306 238170 309374 238226
rect 309430 238170 309498 238226
rect 309554 238170 309622 238226
rect 309678 238170 327250 238226
rect 327306 238170 327374 238226
rect 327430 238170 327498 238226
rect 327554 238170 327622 238226
rect 327678 238170 345250 238226
rect 345306 238170 345374 238226
rect 345430 238170 345498 238226
rect 345554 238170 345622 238226
rect 345678 238170 363250 238226
rect 363306 238170 363374 238226
rect 363430 238170 363498 238226
rect 363554 238170 363622 238226
rect 363678 238170 381250 238226
rect 381306 238170 381374 238226
rect 381430 238170 381498 238226
rect 381554 238170 381622 238226
rect 381678 238170 399250 238226
rect 399306 238170 399374 238226
rect 399430 238170 399498 238226
rect 399554 238170 399622 238226
rect 399678 238170 417250 238226
rect 417306 238170 417374 238226
rect 417430 238170 417498 238226
rect 417554 238170 417622 238226
rect 417678 238170 435250 238226
rect 435306 238170 435374 238226
rect 435430 238170 435498 238226
rect 435554 238170 435622 238226
rect 435678 238170 453250 238226
rect 453306 238170 453374 238226
rect 453430 238170 453498 238226
rect 453554 238170 453622 238226
rect 453678 238170 471250 238226
rect 471306 238170 471374 238226
rect 471430 238170 471498 238226
rect 471554 238170 471622 238226
rect 471678 238170 489250 238226
rect 489306 238170 489374 238226
rect 489430 238170 489498 238226
rect 489554 238170 489622 238226
rect 489678 238170 507250 238226
rect 507306 238170 507374 238226
rect 507430 238170 507498 238226
rect 507554 238170 507622 238226
rect 507678 238170 525250 238226
rect 525306 238170 525374 238226
rect 525430 238170 525498 238226
rect 525554 238170 525622 238226
rect 525678 238170 543250 238226
rect 543306 238170 543374 238226
rect 543430 238170 543498 238226
rect 543554 238170 543622 238226
rect 543678 238170 561250 238226
rect 561306 238170 561374 238226
rect 561430 238170 561498 238226
rect 561554 238170 561622 238226
rect 561678 238170 579250 238226
rect 579306 238170 579374 238226
rect 579430 238170 579498 238226
rect 579554 238170 579622 238226
rect 579678 238170 596496 238226
rect 596552 238170 596620 238226
rect 596676 238170 596744 238226
rect 596800 238170 596868 238226
rect 596924 238170 597980 238226
rect -1916 238102 597980 238170
rect -1916 238046 -860 238102
rect -804 238046 -736 238102
rect -680 238046 -612 238102
rect -556 238046 -488 238102
rect -432 238046 3250 238102
rect 3306 238046 3374 238102
rect 3430 238046 3498 238102
rect 3554 238046 3622 238102
rect 3678 238046 21250 238102
rect 21306 238046 21374 238102
rect 21430 238046 21498 238102
rect 21554 238046 21622 238102
rect 21678 238046 39250 238102
rect 39306 238046 39374 238102
rect 39430 238046 39498 238102
rect 39554 238046 39622 238102
rect 39678 238046 57250 238102
rect 57306 238046 57374 238102
rect 57430 238046 57498 238102
rect 57554 238046 57622 238102
rect 57678 238046 75250 238102
rect 75306 238046 75374 238102
rect 75430 238046 75498 238102
rect 75554 238046 75622 238102
rect 75678 238046 93250 238102
rect 93306 238046 93374 238102
rect 93430 238046 93498 238102
rect 93554 238046 93622 238102
rect 93678 238046 111250 238102
rect 111306 238046 111374 238102
rect 111430 238046 111498 238102
rect 111554 238046 111622 238102
rect 111678 238046 129250 238102
rect 129306 238046 129374 238102
rect 129430 238046 129498 238102
rect 129554 238046 129622 238102
rect 129678 238046 147250 238102
rect 147306 238046 147374 238102
rect 147430 238046 147498 238102
rect 147554 238046 147622 238102
rect 147678 238046 165250 238102
rect 165306 238046 165374 238102
rect 165430 238046 165498 238102
rect 165554 238046 165622 238102
rect 165678 238046 183250 238102
rect 183306 238046 183374 238102
rect 183430 238046 183498 238102
rect 183554 238046 183622 238102
rect 183678 238046 201250 238102
rect 201306 238046 201374 238102
rect 201430 238046 201498 238102
rect 201554 238046 201622 238102
rect 201678 238046 219250 238102
rect 219306 238046 219374 238102
rect 219430 238046 219498 238102
rect 219554 238046 219622 238102
rect 219678 238046 237250 238102
rect 237306 238046 237374 238102
rect 237430 238046 237498 238102
rect 237554 238046 237622 238102
rect 237678 238046 255250 238102
rect 255306 238046 255374 238102
rect 255430 238046 255498 238102
rect 255554 238046 255622 238102
rect 255678 238046 273250 238102
rect 273306 238046 273374 238102
rect 273430 238046 273498 238102
rect 273554 238046 273622 238102
rect 273678 238046 291250 238102
rect 291306 238046 291374 238102
rect 291430 238046 291498 238102
rect 291554 238046 291622 238102
rect 291678 238046 309250 238102
rect 309306 238046 309374 238102
rect 309430 238046 309498 238102
rect 309554 238046 309622 238102
rect 309678 238046 327250 238102
rect 327306 238046 327374 238102
rect 327430 238046 327498 238102
rect 327554 238046 327622 238102
rect 327678 238046 345250 238102
rect 345306 238046 345374 238102
rect 345430 238046 345498 238102
rect 345554 238046 345622 238102
rect 345678 238046 363250 238102
rect 363306 238046 363374 238102
rect 363430 238046 363498 238102
rect 363554 238046 363622 238102
rect 363678 238046 381250 238102
rect 381306 238046 381374 238102
rect 381430 238046 381498 238102
rect 381554 238046 381622 238102
rect 381678 238046 399250 238102
rect 399306 238046 399374 238102
rect 399430 238046 399498 238102
rect 399554 238046 399622 238102
rect 399678 238046 417250 238102
rect 417306 238046 417374 238102
rect 417430 238046 417498 238102
rect 417554 238046 417622 238102
rect 417678 238046 435250 238102
rect 435306 238046 435374 238102
rect 435430 238046 435498 238102
rect 435554 238046 435622 238102
rect 435678 238046 453250 238102
rect 453306 238046 453374 238102
rect 453430 238046 453498 238102
rect 453554 238046 453622 238102
rect 453678 238046 471250 238102
rect 471306 238046 471374 238102
rect 471430 238046 471498 238102
rect 471554 238046 471622 238102
rect 471678 238046 489250 238102
rect 489306 238046 489374 238102
rect 489430 238046 489498 238102
rect 489554 238046 489622 238102
rect 489678 238046 507250 238102
rect 507306 238046 507374 238102
rect 507430 238046 507498 238102
rect 507554 238046 507622 238102
rect 507678 238046 525250 238102
rect 525306 238046 525374 238102
rect 525430 238046 525498 238102
rect 525554 238046 525622 238102
rect 525678 238046 543250 238102
rect 543306 238046 543374 238102
rect 543430 238046 543498 238102
rect 543554 238046 543622 238102
rect 543678 238046 561250 238102
rect 561306 238046 561374 238102
rect 561430 238046 561498 238102
rect 561554 238046 561622 238102
rect 561678 238046 579250 238102
rect 579306 238046 579374 238102
rect 579430 238046 579498 238102
rect 579554 238046 579622 238102
rect 579678 238046 596496 238102
rect 596552 238046 596620 238102
rect 596676 238046 596744 238102
rect 596800 238046 596868 238102
rect 596924 238046 597980 238102
rect -1916 237978 597980 238046
rect -1916 237922 -860 237978
rect -804 237922 -736 237978
rect -680 237922 -612 237978
rect -556 237922 -488 237978
rect -432 237922 3250 237978
rect 3306 237922 3374 237978
rect 3430 237922 3498 237978
rect 3554 237922 3622 237978
rect 3678 237922 21250 237978
rect 21306 237922 21374 237978
rect 21430 237922 21498 237978
rect 21554 237922 21622 237978
rect 21678 237922 39250 237978
rect 39306 237922 39374 237978
rect 39430 237922 39498 237978
rect 39554 237922 39622 237978
rect 39678 237922 57250 237978
rect 57306 237922 57374 237978
rect 57430 237922 57498 237978
rect 57554 237922 57622 237978
rect 57678 237922 75250 237978
rect 75306 237922 75374 237978
rect 75430 237922 75498 237978
rect 75554 237922 75622 237978
rect 75678 237922 93250 237978
rect 93306 237922 93374 237978
rect 93430 237922 93498 237978
rect 93554 237922 93622 237978
rect 93678 237922 111250 237978
rect 111306 237922 111374 237978
rect 111430 237922 111498 237978
rect 111554 237922 111622 237978
rect 111678 237922 129250 237978
rect 129306 237922 129374 237978
rect 129430 237922 129498 237978
rect 129554 237922 129622 237978
rect 129678 237922 147250 237978
rect 147306 237922 147374 237978
rect 147430 237922 147498 237978
rect 147554 237922 147622 237978
rect 147678 237922 165250 237978
rect 165306 237922 165374 237978
rect 165430 237922 165498 237978
rect 165554 237922 165622 237978
rect 165678 237922 183250 237978
rect 183306 237922 183374 237978
rect 183430 237922 183498 237978
rect 183554 237922 183622 237978
rect 183678 237922 201250 237978
rect 201306 237922 201374 237978
rect 201430 237922 201498 237978
rect 201554 237922 201622 237978
rect 201678 237922 219250 237978
rect 219306 237922 219374 237978
rect 219430 237922 219498 237978
rect 219554 237922 219622 237978
rect 219678 237922 237250 237978
rect 237306 237922 237374 237978
rect 237430 237922 237498 237978
rect 237554 237922 237622 237978
rect 237678 237922 255250 237978
rect 255306 237922 255374 237978
rect 255430 237922 255498 237978
rect 255554 237922 255622 237978
rect 255678 237922 273250 237978
rect 273306 237922 273374 237978
rect 273430 237922 273498 237978
rect 273554 237922 273622 237978
rect 273678 237922 291250 237978
rect 291306 237922 291374 237978
rect 291430 237922 291498 237978
rect 291554 237922 291622 237978
rect 291678 237922 309250 237978
rect 309306 237922 309374 237978
rect 309430 237922 309498 237978
rect 309554 237922 309622 237978
rect 309678 237922 327250 237978
rect 327306 237922 327374 237978
rect 327430 237922 327498 237978
rect 327554 237922 327622 237978
rect 327678 237922 345250 237978
rect 345306 237922 345374 237978
rect 345430 237922 345498 237978
rect 345554 237922 345622 237978
rect 345678 237922 363250 237978
rect 363306 237922 363374 237978
rect 363430 237922 363498 237978
rect 363554 237922 363622 237978
rect 363678 237922 381250 237978
rect 381306 237922 381374 237978
rect 381430 237922 381498 237978
rect 381554 237922 381622 237978
rect 381678 237922 399250 237978
rect 399306 237922 399374 237978
rect 399430 237922 399498 237978
rect 399554 237922 399622 237978
rect 399678 237922 417250 237978
rect 417306 237922 417374 237978
rect 417430 237922 417498 237978
rect 417554 237922 417622 237978
rect 417678 237922 435250 237978
rect 435306 237922 435374 237978
rect 435430 237922 435498 237978
rect 435554 237922 435622 237978
rect 435678 237922 453250 237978
rect 453306 237922 453374 237978
rect 453430 237922 453498 237978
rect 453554 237922 453622 237978
rect 453678 237922 471250 237978
rect 471306 237922 471374 237978
rect 471430 237922 471498 237978
rect 471554 237922 471622 237978
rect 471678 237922 489250 237978
rect 489306 237922 489374 237978
rect 489430 237922 489498 237978
rect 489554 237922 489622 237978
rect 489678 237922 507250 237978
rect 507306 237922 507374 237978
rect 507430 237922 507498 237978
rect 507554 237922 507622 237978
rect 507678 237922 525250 237978
rect 525306 237922 525374 237978
rect 525430 237922 525498 237978
rect 525554 237922 525622 237978
rect 525678 237922 543250 237978
rect 543306 237922 543374 237978
rect 543430 237922 543498 237978
rect 543554 237922 543622 237978
rect 543678 237922 561250 237978
rect 561306 237922 561374 237978
rect 561430 237922 561498 237978
rect 561554 237922 561622 237978
rect 561678 237922 579250 237978
rect 579306 237922 579374 237978
rect 579430 237922 579498 237978
rect 579554 237922 579622 237978
rect 579678 237922 596496 237978
rect 596552 237922 596620 237978
rect 596676 237922 596744 237978
rect 596800 237922 596868 237978
rect 596924 237922 597980 237978
rect -1916 237826 597980 237922
rect -1916 226350 597980 226446
rect -1916 226294 -1820 226350
rect -1764 226294 -1696 226350
rect -1640 226294 -1572 226350
rect -1516 226294 -1448 226350
rect -1392 226294 6970 226350
rect 7026 226294 7094 226350
rect 7150 226294 7218 226350
rect 7274 226294 7342 226350
rect 7398 226294 24970 226350
rect 25026 226294 25094 226350
rect 25150 226294 25218 226350
rect 25274 226294 25342 226350
rect 25398 226294 42970 226350
rect 43026 226294 43094 226350
rect 43150 226294 43218 226350
rect 43274 226294 43342 226350
rect 43398 226294 60970 226350
rect 61026 226294 61094 226350
rect 61150 226294 61218 226350
rect 61274 226294 61342 226350
rect 61398 226294 78970 226350
rect 79026 226294 79094 226350
rect 79150 226294 79218 226350
rect 79274 226294 79342 226350
rect 79398 226294 79878 226350
rect 79934 226294 80002 226350
rect 80058 226294 96970 226350
rect 97026 226294 97094 226350
rect 97150 226294 97218 226350
rect 97274 226294 97342 226350
rect 97398 226294 110598 226350
rect 110654 226294 110722 226350
rect 110778 226294 114970 226350
rect 115026 226294 115094 226350
rect 115150 226294 115218 226350
rect 115274 226294 115342 226350
rect 115398 226294 132970 226350
rect 133026 226294 133094 226350
rect 133150 226294 133218 226350
rect 133274 226294 133342 226350
rect 133398 226294 141318 226350
rect 141374 226294 141442 226350
rect 141498 226294 150970 226350
rect 151026 226294 151094 226350
rect 151150 226294 151218 226350
rect 151274 226294 151342 226350
rect 151398 226294 168970 226350
rect 169026 226294 169094 226350
rect 169150 226294 169218 226350
rect 169274 226294 169342 226350
rect 169398 226294 172038 226350
rect 172094 226294 172162 226350
rect 172218 226294 202758 226350
rect 202814 226294 202882 226350
rect 202938 226294 204970 226350
rect 205026 226294 205094 226350
rect 205150 226294 205218 226350
rect 205274 226294 205342 226350
rect 205398 226294 222970 226350
rect 223026 226294 223094 226350
rect 223150 226294 223218 226350
rect 223274 226294 223342 226350
rect 223398 226294 233478 226350
rect 233534 226294 233602 226350
rect 233658 226294 240970 226350
rect 241026 226294 241094 226350
rect 241150 226294 241218 226350
rect 241274 226294 241342 226350
rect 241398 226294 258970 226350
rect 259026 226294 259094 226350
rect 259150 226294 259218 226350
rect 259274 226294 259342 226350
rect 259398 226294 276970 226350
rect 277026 226294 277094 226350
rect 277150 226294 277218 226350
rect 277274 226294 277342 226350
rect 277398 226294 294970 226350
rect 295026 226294 295094 226350
rect 295150 226294 295218 226350
rect 295274 226294 295342 226350
rect 295398 226294 312970 226350
rect 313026 226294 313094 226350
rect 313150 226294 313218 226350
rect 313274 226294 313342 226350
rect 313398 226294 330970 226350
rect 331026 226294 331094 226350
rect 331150 226294 331218 226350
rect 331274 226294 331342 226350
rect 331398 226294 348970 226350
rect 349026 226294 349094 226350
rect 349150 226294 349218 226350
rect 349274 226294 349342 226350
rect 349398 226294 366970 226350
rect 367026 226294 367094 226350
rect 367150 226294 367218 226350
rect 367274 226294 367342 226350
rect 367398 226294 402970 226350
rect 403026 226294 403094 226350
rect 403150 226294 403218 226350
rect 403274 226294 403342 226350
rect 403398 226294 420970 226350
rect 421026 226294 421094 226350
rect 421150 226294 421218 226350
rect 421274 226294 421342 226350
rect 421398 226294 438970 226350
rect 439026 226294 439094 226350
rect 439150 226294 439218 226350
rect 439274 226294 439342 226350
rect 439398 226294 456970 226350
rect 457026 226294 457094 226350
rect 457150 226294 457218 226350
rect 457274 226294 457342 226350
rect 457398 226294 492970 226350
rect 493026 226294 493094 226350
rect 493150 226294 493218 226350
rect 493274 226294 493342 226350
rect 493398 226294 510970 226350
rect 511026 226294 511094 226350
rect 511150 226294 511218 226350
rect 511274 226294 511342 226350
rect 511398 226294 528970 226350
rect 529026 226294 529094 226350
rect 529150 226294 529218 226350
rect 529274 226294 529342 226350
rect 529398 226294 546970 226350
rect 547026 226294 547094 226350
rect 547150 226294 547218 226350
rect 547274 226294 547342 226350
rect 547398 226294 564970 226350
rect 565026 226294 565094 226350
rect 565150 226294 565218 226350
rect 565274 226294 565342 226350
rect 565398 226294 582970 226350
rect 583026 226294 583094 226350
rect 583150 226294 583218 226350
rect 583274 226294 583342 226350
rect 583398 226294 597456 226350
rect 597512 226294 597580 226350
rect 597636 226294 597704 226350
rect 597760 226294 597828 226350
rect 597884 226294 597980 226350
rect -1916 226226 597980 226294
rect -1916 226170 -1820 226226
rect -1764 226170 -1696 226226
rect -1640 226170 -1572 226226
rect -1516 226170 -1448 226226
rect -1392 226170 6970 226226
rect 7026 226170 7094 226226
rect 7150 226170 7218 226226
rect 7274 226170 7342 226226
rect 7398 226170 24970 226226
rect 25026 226170 25094 226226
rect 25150 226170 25218 226226
rect 25274 226170 25342 226226
rect 25398 226170 42970 226226
rect 43026 226170 43094 226226
rect 43150 226170 43218 226226
rect 43274 226170 43342 226226
rect 43398 226170 60970 226226
rect 61026 226170 61094 226226
rect 61150 226170 61218 226226
rect 61274 226170 61342 226226
rect 61398 226170 78970 226226
rect 79026 226170 79094 226226
rect 79150 226170 79218 226226
rect 79274 226170 79342 226226
rect 79398 226170 79878 226226
rect 79934 226170 80002 226226
rect 80058 226170 96970 226226
rect 97026 226170 97094 226226
rect 97150 226170 97218 226226
rect 97274 226170 97342 226226
rect 97398 226170 110598 226226
rect 110654 226170 110722 226226
rect 110778 226170 114970 226226
rect 115026 226170 115094 226226
rect 115150 226170 115218 226226
rect 115274 226170 115342 226226
rect 115398 226170 132970 226226
rect 133026 226170 133094 226226
rect 133150 226170 133218 226226
rect 133274 226170 133342 226226
rect 133398 226170 141318 226226
rect 141374 226170 141442 226226
rect 141498 226170 150970 226226
rect 151026 226170 151094 226226
rect 151150 226170 151218 226226
rect 151274 226170 151342 226226
rect 151398 226170 168970 226226
rect 169026 226170 169094 226226
rect 169150 226170 169218 226226
rect 169274 226170 169342 226226
rect 169398 226170 172038 226226
rect 172094 226170 172162 226226
rect 172218 226170 202758 226226
rect 202814 226170 202882 226226
rect 202938 226170 204970 226226
rect 205026 226170 205094 226226
rect 205150 226170 205218 226226
rect 205274 226170 205342 226226
rect 205398 226170 222970 226226
rect 223026 226170 223094 226226
rect 223150 226170 223218 226226
rect 223274 226170 223342 226226
rect 223398 226170 233478 226226
rect 233534 226170 233602 226226
rect 233658 226170 240970 226226
rect 241026 226170 241094 226226
rect 241150 226170 241218 226226
rect 241274 226170 241342 226226
rect 241398 226170 258970 226226
rect 259026 226170 259094 226226
rect 259150 226170 259218 226226
rect 259274 226170 259342 226226
rect 259398 226170 276970 226226
rect 277026 226170 277094 226226
rect 277150 226170 277218 226226
rect 277274 226170 277342 226226
rect 277398 226170 294970 226226
rect 295026 226170 295094 226226
rect 295150 226170 295218 226226
rect 295274 226170 295342 226226
rect 295398 226170 312970 226226
rect 313026 226170 313094 226226
rect 313150 226170 313218 226226
rect 313274 226170 313342 226226
rect 313398 226170 330970 226226
rect 331026 226170 331094 226226
rect 331150 226170 331218 226226
rect 331274 226170 331342 226226
rect 331398 226170 348970 226226
rect 349026 226170 349094 226226
rect 349150 226170 349218 226226
rect 349274 226170 349342 226226
rect 349398 226170 366970 226226
rect 367026 226170 367094 226226
rect 367150 226170 367218 226226
rect 367274 226170 367342 226226
rect 367398 226170 402970 226226
rect 403026 226170 403094 226226
rect 403150 226170 403218 226226
rect 403274 226170 403342 226226
rect 403398 226170 420970 226226
rect 421026 226170 421094 226226
rect 421150 226170 421218 226226
rect 421274 226170 421342 226226
rect 421398 226170 438970 226226
rect 439026 226170 439094 226226
rect 439150 226170 439218 226226
rect 439274 226170 439342 226226
rect 439398 226170 456970 226226
rect 457026 226170 457094 226226
rect 457150 226170 457218 226226
rect 457274 226170 457342 226226
rect 457398 226170 492970 226226
rect 493026 226170 493094 226226
rect 493150 226170 493218 226226
rect 493274 226170 493342 226226
rect 493398 226170 510970 226226
rect 511026 226170 511094 226226
rect 511150 226170 511218 226226
rect 511274 226170 511342 226226
rect 511398 226170 528970 226226
rect 529026 226170 529094 226226
rect 529150 226170 529218 226226
rect 529274 226170 529342 226226
rect 529398 226170 546970 226226
rect 547026 226170 547094 226226
rect 547150 226170 547218 226226
rect 547274 226170 547342 226226
rect 547398 226170 564970 226226
rect 565026 226170 565094 226226
rect 565150 226170 565218 226226
rect 565274 226170 565342 226226
rect 565398 226170 582970 226226
rect 583026 226170 583094 226226
rect 583150 226170 583218 226226
rect 583274 226170 583342 226226
rect 583398 226170 597456 226226
rect 597512 226170 597580 226226
rect 597636 226170 597704 226226
rect 597760 226170 597828 226226
rect 597884 226170 597980 226226
rect -1916 226102 597980 226170
rect -1916 226046 -1820 226102
rect -1764 226046 -1696 226102
rect -1640 226046 -1572 226102
rect -1516 226046 -1448 226102
rect -1392 226046 6970 226102
rect 7026 226046 7094 226102
rect 7150 226046 7218 226102
rect 7274 226046 7342 226102
rect 7398 226046 24970 226102
rect 25026 226046 25094 226102
rect 25150 226046 25218 226102
rect 25274 226046 25342 226102
rect 25398 226046 42970 226102
rect 43026 226046 43094 226102
rect 43150 226046 43218 226102
rect 43274 226046 43342 226102
rect 43398 226046 60970 226102
rect 61026 226046 61094 226102
rect 61150 226046 61218 226102
rect 61274 226046 61342 226102
rect 61398 226046 78970 226102
rect 79026 226046 79094 226102
rect 79150 226046 79218 226102
rect 79274 226046 79342 226102
rect 79398 226046 79878 226102
rect 79934 226046 80002 226102
rect 80058 226046 96970 226102
rect 97026 226046 97094 226102
rect 97150 226046 97218 226102
rect 97274 226046 97342 226102
rect 97398 226046 110598 226102
rect 110654 226046 110722 226102
rect 110778 226046 114970 226102
rect 115026 226046 115094 226102
rect 115150 226046 115218 226102
rect 115274 226046 115342 226102
rect 115398 226046 132970 226102
rect 133026 226046 133094 226102
rect 133150 226046 133218 226102
rect 133274 226046 133342 226102
rect 133398 226046 141318 226102
rect 141374 226046 141442 226102
rect 141498 226046 150970 226102
rect 151026 226046 151094 226102
rect 151150 226046 151218 226102
rect 151274 226046 151342 226102
rect 151398 226046 168970 226102
rect 169026 226046 169094 226102
rect 169150 226046 169218 226102
rect 169274 226046 169342 226102
rect 169398 226046 172038 226102
rect 172094 226046 172162 226102
rect 172218 226046 202758 226102
rect 202814 226046 202882 226102
rect 202938 226046 204970 226102
rect 205026 226046 205094 226102
rect 205150 226046 205218 226102
rect 205274 226046 205342 226102
rect 205398 226046 222970 226102
rect 223026 226046 223094 226102
rect 223150 226046 223218 226102
rect 223274 226046 223342 226102
rect 223398 226046 233478 226102
rect 233534 226046 233602 226102
rect 233658 226046 240970 226102
rect 241026 226046 241094 226102
rect 241150 226046 241218 226102
rect 241274 226046 241342 226102
rect 241398 226046 258970 226102
rect 259026 226046 259094 226102
rect 259150 226046 259218 226102
rect 259274 226046 259342 226102
rect 259398 226046 276970 226102
rect 277026 226046 277094 226102
rect 277150 226046 277218 226102
rect 277274 226046 277342 226102
rect 277398 226046 294970 226102
rect 295026 226046 295094 226102
rect 295150 226046 295218 226102
rect 295274 226046 295342 226102
rect 295398 226046 312970 226102
rect 313026 226046 313094 226102
rect 313150 226046 313218 226102
rect 313274 226046 313342 226102
rect 313398 226046 330970 226102
rect 331026 226046 331094 226102
rect 331150 226046 331218 226102
rect 331274 226046 331342 226102
rect 331398 226046 348970 226102
rect 349026 226046 349094 226102
rect 349150 226046 349218 226102
rect 349274 226046 349342 226102
rect 349398 226046 366970 226102
rect 367026 226046 367094 226102
rect 367150 226046 367218 226102
rect 367274 226046 367342 226102
rect 367398 226046 402970 226102
rect 403026 226046 403094 226102
rect 403150 226046 403218 226102
rect 403274 226046 403342 226102
rect 403398 226046 420970 226102
rect 421026 226046 421094 226102
rect 421150 226046 421218 226102
rect 421274 226046 421342 226102
rect 421398 226046 438970 226102
rect 439026 226046 439094 226102
rect 439150 226046 439218 226102
rect 439274 226046 439342 226102
rect 439398 226046 456970 226102
rect 457026 226046 457094 226102
rect 457150 226046 457218 226102
rect 457274 226046 457342 226102
rect 457398 226046 492970 226102
rect 493026 226046 493094 226102
rect 493150 226046 493218 226102
rect 493274 226046 493342 226102
rect 493398 226046 510970 226102
rect 511026 226046 511094 226102
rect 511150 226046 511218 226102
rect 511274 226046 511342 226102
rect 511398 226046 528970 226102
rect 529026 226046 529094 226102
rect 529150 226046 529218 226102
rect 529274 226046 529342 226102
rect 529398 226046 546970 226102
rect 547026 226046 547094 226102
rect 547150 226046 547218 226102
rect 547274 226046 547342 226102
rect 547398 226046 564970 226102
rect 565026 226046 565094 226102
rect 565150 226046 565218 226102
rect 565274 226046 565342 226102
rect 565398 226046 582970 226102
rect 583026 226046 583094 226102
rect 583150 226046 583218 226102
rect 583274 226046 583342 226102
rect 583398 226046 597456 226102
rect 597512 226046 597580 226102
rect 597636 226046 597704 226102
rect 597760 226046 597828 226102
rect 597884 226046 597980 226102
rect -1916 225978 597980 226046
rect -1916 225922 -1820 225978
rect -1764 225922 -1696 225978
rect -1640 225922 -1572 225978
rect -1516 225922 -1448 225978
rect -1392 225922 6970 225978
rect 7026 225922 7094 225978
rect 7150 225922 7218 225978
rect 7274 225922 7342 225978
rect 7398 225922 24970 225978
rect 25026 225922 25094 225978
rect 25150 225922 25218 225978
rect 25274 225922 25342 225978
rect 25398 225922 42970 225978
rect 43026 225922 43094 225978
rect 43150 225922 43218 225978
rect 43274 225922 43342 225978
rect 43398 225922 60970 225978
rect 61026 225922 61094 225978
rect 61150 225922 61218 225978
rect 61274 225922 61342 225978
rect 61398 225922 78970 225978
rect 79026 225922 79094 225978
rect 79150 225922 79218 225978
rect 79274 225922 79342 225978
rect 79398 225922 79878 225978
rect 79934 225922 80002 225978
rect 80058 225922 96970 225978
rect 97026 225922 97094 225978
rect 97150 225922 97218 225978
rect 97274 225922 97342 225978
rect 97398 225922 110598 225978
rect 110654 225922 110722 225978
rect 110778 225922 114970 225978
rect 115026 225922 115094 225978
rect 115150 225922 115218 225978
rect 115274 225922 115342 225978
rect 115398 225922 132970 225978
rect 133026 225922 133094 225978
rect 133150 225922 133218 225978
rect 133274 225922 133342 225978
rect 133398 225922 141318 225978
rect 141374 225922 141442 225978
rect 141498 225922 150970 225978
rect 151026 225922 151094 225978
rect 151150 225922 151218 225978
rect 151274 225922 151342 225978
rect 151398 225922 168970 225978
rect 169026 225922 169094 225978
rect 169150 225922 169218 225978
rect 169274 225922 169342 225978
rect 169398 225922 172038 225978
rect 172094 225922 172162 225978
rect 172218 225922 202758 225978
rect 202814 225922 202882 225978
rect 202938 225922 204970 225978
rect 205026 225922 205094 225978
rect 205150 225922 205218 225978
rect 205274 225922 205342 225978
rect 205398 225922 222970 225978
rect 223026 225922 223094 225978
rect 223150 225922 223218 225978
rect 223274 225922 223342 225978
rect 223398 225922 233478 225978
rect 233534 225922 233602 225978
rect 233658 225922 240970 225978
rect 241026 225922 241094 225978
rect 241150 225922 241218 225978
rect 241274 225922 241342 225978
rect 241398 225922 258970 225978
rect 259026 225922 259094 225978
rect 259150 225922 259218 225978
rect 259274 225922 259342 225978
rect 259398 225922 276970 225978
rect 277026 225922 277094 225978
rect 277150 225922 277218 225978
rect 277274 225922 277342 225978
rect 277398 225922 294970 225978
rect 295026 225922 295094 225978
rect 295150 225922 295218 225978
rect 295274 225922 295342 225978
rect 295398 225922 312970 225978
rect 313026 225922 313094 225978
rect 313150 225922 313218 225978
rect 313274 225922 313342 225978
rect 313398 225922 330970 225978
rect 331026 225922 331094 225978
rect 331150 225922 331218 225978
rect 331274 225922 331342 225978
rect 331398 225922 348970 225978
rect 349026 225922 349094 225978
rect 349150 225922 349218 225978
rect 349274 225922 349342 225978
rect 349398 225922 366970 225978
rect 367026 225922 367094 225978
rect 367150 225922 367218 225978
rect 367274 225922 367342 225978
rect 367398 225922 402970 225978
rect 403026 225922 403094 225978
rect 403150 225922 403218 225978
rect 403274 225922 403342 225978
rect 403398 225922 420970 225978
rect 421026 225922 421094 225978
rect 421150 225922 421218 225978
rect 421274 225922 421342 225978
rect 421398 225922 438970 225978
rect 439026 225922 439094 225978
rect 439150 225922 439218 225978
rect 439274 225922 439342 225978
rect 439398 225922 456970 225978
rect 457026 225922 457094 225978
rect 457150 225922 457218 225978
rect 457274 225922 457342 225978
rect 457398 225922 492970 225978
rect 493026 225922 493094 225978
rect 493150 225922 493218 225978
rect 493274 225922 493342 225978
rect 493398 225922 510970 225978
rect 511026 225922 511094 225978
rect 511150 225922 511218 225978
rect 511274 225922 511342 225978
rect 511398 225922 528970 225978
rect 529026 225922 529094 225978
rect 529150 225922 529218 225978
rect 529274 225922 529342 225978
rect 529398 225922 546970 225978
rect 547026 225922 547094 225978
rect 547150 225922 547218 225978
rect 547274 225922 547342 225978
rect 547398 225922 564970 225978
rect 565026 225922 565094 225978
rect 565150 225922 565218 225978
rect 565274 225922 565342 225978
rect 565398 225922 582970 225978
rect 583026 225922 583094 225978
rect 583150 225922 583218 225978
rect 583274 225922 583342 225978
rect 583398 225922 597456 225978
rect 597512 225922 597580 225978
rect 597636 225922 597704 225978
rect 597760 225922 597828 225978
rect 597884 225922 597980 225978
rect -1916 225826 597980 225922
rect -1916 220350 597980 220446
rect -1916 220294 -860 220350
rect -804 220294 -736 220350
rect -680 220294 -612 220350
rect -556 220294 -488 220350
rect -432 220294 3250 220350
rect 3306 220294 3374 220350
rect 3430 220294 3498 220350
rect 3554 220294 3622 220350
rect 3678 220294 21250 220350
rect 21306 220294 21374 220350
rect 21430 220294 21498 220350
rect 21554 220294 21622 220350
rect 21678 220294 39250 220350
rect 39306 220294 39374 220350
rect 39430 220294 39498 220350
rect 39554 220294 39622 220350
rect 39678 220294 57250 220350
rect 57306 220294 57374 220350
rect 57430 220294 57498 220350
rect 57554 220294 57622 220350
rect 57678 220294 64518 220350
rect 64574 220294 64642 220350
rect 64698 220294 75250 220350
rect 75306 220294 75374 220350
rect 75430 220294 75498 220350
rect 75554 220294 75622 220350
rect 75678 220294 93250 220350
rect 93306 220294 93374 220350
rect 93430 220294 93498 220350
rect 93554 220294 93622 220350
rect 93678 220294 95238 220350
rect 95294 220294 95362 220350
rect 95418 220294 111250 220350
rect 111306 220294 111374 220350
rect 111430 220294 111498 220350
rect 111554 220294 111622 220350
rect 111678 220294 125958 220350
rect 126014 220294 126082 220350
rect 126138 220294 129250 220350
rect 129306 220294 129374 220350
rect 129430 220294 129498 220350
rect 129554 220294 129622 220350
rect 129678 220294 147250 220350
rect 147306 220294 147374 220350
rect 147430 220294 147498 220350
rect 147554 220294 147622 220350
rect 147678 220294 156678 220350
rect 156734 220294 156802 220350
rect 156858 220294 165250 220350
rect 165306 220294 165374 220350
rect 165430 220294 165498 220350
rect 165554 220294 165622 220350
rect 165678 220294 183250 220350
rect 183306 220294 183374 220350
rect 183430 220294 183498 220350
rect 183554 220294 183622 220350
rect 183678 220294 187398 220350
rect 187454 220294 187522 220350
rect 187578 220294 201250 220350
rect 201306 220294 201374 220350
rect 201430 220294 201498 220350
rect 201554 220294 201622 220350
rect 201678 220294 218118 220350
rect 218174 220294 218242 220350
rect 218298 220294 219250 220350
rect 219306 220294 219374 220350
rect 219430 220294 219498 220350
rect 219554 220294 219622 220350
rect 219678 220294 237250 220350
rect 237306 220294 237374 220350
rect 237430 220294 237498 220350
rect 237554 220294 237622 220350
rect 237678 220294 255250 220350
rect 255306 220294 255374 220350
rect 255430 220294 255498 220350
rect 255554 220294 255622 220350
rect 255678 220294 273250 220350
rect 273306 220294 273374 220350
rect 273430 220294 273498 220350
rect 273554 220294 273622 220350
rect 273678 220294 291250 220350
rect 291306 220294 291374 220350
rect 291430 220294 291498 220350
rect 291554 220294 291622 220350
rect 291678 220294 309250 220350
rect 309306 220294 309374 220350
rect 309430 220294 309498 220350
rect 309554 220294 309622 220350
rect 309678 220294 327250 220350
rect 327306 220294 327374 220350
rect 327430 220294 327498 220350
rect 327554 220294 327622 220350
rect 327678 220294 345250 220350
rect 345306 220294 345374 220350
rect 345430 220294 345498 220350
rect 345554 220294 345622 220350
rect 345678 220294 363250 220350
rect 363306 220294 363374 220350
rect 363430 220294 363498 220350
rect 363554 220294 363622 220350
rect 363678 220294 381250 220350
rect 381306 220294 381374 220350
rect 381430 220294 381498 220350
rect 381554 220294 381622 220350
rect 381678 220294 399250 220350
rect 399306 220294 399374 220350
rect 399430 220294 399498 220350
rect 399554 220294 399622 220350
rect 399678 220294 417250 220350
rect 417306 220294 417374 220350
rect 417430 220294 417498 220350
rect 417554 220294 417622 220350
rect 417678 220294 435250 220350
rect 435306 220294 435374 220350
rect 435430 220294 435498 220350
rect 435554 220294 435622 220350
rect 435678 220294 453250 220350
rect 453306 220294 453374 220350
rect 453430 220294 453498 220350
rect 453554 220294 453622 220350
rect 453678 220294 471250 220350
rect 471306 220294 471374 220350
rect 471430 220294 471498 220350
rect 471554 220294 471622 220350
rect 471678 220294 489250 220350
rect 489306 220294 489374 220350
rect 489430 220294 489498 220350
rect 489554 220294 489622 220350
rect 489678 220294 507250 220350
rect 507306 220294 507374 220350
rect 507430 220294 507498 220350
rect 507554 220294 507622 220350
rect 507678 220294 525250 220350
rect 525306 220294 525374 220350
rect 525430 220294 525498 220350
rect 525554 220294 525622 220350
rect 525678 220294 543250 220350
rect 543306 220294 543374 220350
rect 543430 220294 543498 220350
rect 543554 220294 543622 220350
rect 543678 220294 561250 220350
rect 561306 220294 561374 220350
rect 561430 220294 561498 220350
rect 561554 220294 561622 220350
rect 561678 220294 579250 220350
rect 579306 220294 579374 220350
rect 579430 220294 579498 220350
rect 579554 220294 579622 220350
rect 579678 220294 596496 220350
rect 596552 220294 596620 220350
rect 596676 220294 596744 220350
rect 596800 220294 596868 220350
rect 596924 220294 597980 220350
rect -1916 220226 597980 220294
rect -1916 220170 -860 220226
rect -804 220170 -736 220226
rect -680 220170 -612 220226
rect -556 220170 -488 220226
rect -432 220170 3250 220226
rect 3306 220170 3374 220226
rect 3430 220170 3498 220226
rect 3554 220170 3622 220226
rect 3678 220170 21250 220226
rect 21306 220170 21374 220226
rect 21430 220170 21498 220226
rect 21554 220170 21622 220226
rect 21678 220170 39250 220226
rect 39306 220170 39374 220226
rect 39430 220170 39498 220226
rect 39554 220170 39622 220226
rect 39678 220170 57250 220226
rect 57306 220170 57374 220226
rect 57430 220170 57498 220226
rect 57554 220170 57622 220226
rect 57678 220170 64518 220226
rect 64574 220170 64642 220226
rect 64698 220170 75250 220226
rect 75306 220170 75374 220226
rect 75430 220170 75498 220226
rect 75554 220170 75622 220226
rect 75678 220170 93250 220226
rect 93306 220170 93374 220226
rect 93430 220170 93498 220226
rect 93554 220170 93622 220226
rect 93678 220170 95238 220226
rect 95294 220170 95362 220226
rect 95418 220170 111250 220226
rect 111306 220170 111374 220226
rect 111430 220170 111498 220226
rect 111554 220170 111622 220226
rect 111678 220170 125958 220226
rect 126014 220170 126082 220226
rect 126138 220170 129250 220226
rect 129306 220170 129374 220226
rect 129430 220170 129498 220226
rect 129554 220170 129622 220226
rect 129678 220170 147250 220226
rect 147306 220170 147374 220226
rect 147430 220170 147498 220226
rect 147554 220170 147622 220226
rect 147678 220170 156678 220226
rect 156734 220170 156802 220226
rect 156858 220170 165250 220226
rect 165306 220170 165374 220226
rect 165430 220170 165498 220226
rect 165554 220170 165622 220226
rect 165678 220170 183250 220226
rect 183306 220170 183374 220226
rect 183430 220170 183498 220226
rect 183554 220170 183622 220226
rect 183678 220170 187398 220226
rect 187454 220170 187522 220226
rect 187578 220170 201250 220226
rect 201306 220170 201374 220226
rect 201430 220170 201498 220226
rect 201554 220170 201622 220226
rect 201678 220170 218118 220226
rect 218174 220170 218242 220226
rect 218298 220170 219250 220226
rect 219306 220170 219374 220226
rect 219430 220170 219498 220226
rect 219554 220170 219622 220226
rect 219678 220170 237250 220226
rect 237306 220170 237374 220226
rect 237430 220170 237498 220226
rect 237554 220170 237622 220226
rect 237678 220170 255250 220226
rect 255306 220170 255374 220226
rect 255430 220170 255498 220226
rect 255554 220170 255622 220226
rect 255678 220170 273250 220226
rect 273306 220170 273374 220226
rect 273430 220170 273498 220226
rect 273554 220170 273622 220226
rect 273678 220170 291250 220226
rect 291306 220170 291374 220226
rect 291430 220170 291498 220226
rect 291554 220170 291622 220226
rect 291678 220170 309250 220226
rect 309306 220170 309374 220226
rect 309430 220170 309498 220226
rect 309554 220170 309622 220226
rect 309678 220170 327250 220226
rect 327306 220170 327374 220226
rect 327430 220170 327498 220226
rect 327554 220170 327622 220226
rect 327678 220170 345250 220226
rect 345306 220170 345374 220226
rect 345430 220170 345498 220226
rect 345554 220170 345622 220226
rect 345678 220170 363250 220226
rect 363306 220170 363374 220226
rect 363430 220170 363498 220226
rect 363554 220170 363622 220226
rect 363678 220170 381250 220226
rect 381306 220170 381374 220226
rect 381430 220170 381498 220226
rect 381554 220170 381622 220226
rect 381678 220170 399250 220226
rect 399306 220170 399374 220226
rect 399430 220170 399498 220226
rect 399554 220170 399622 220226
rect 399678 220170 417250 220226
rect 417306 220170 417374 220226
rect 417430 220170 417498 220226
rect 417554 220170 417622 220226
rect 417678 220170 435250 220226
rect 435306 220170 435374 220226
rect 435430 220170 435498 220226
rect 435554 220170 435622 220226
rect 435678 220170 453250 220226
rect 453306 220170 453374 220226
rect 453430 220170 453498 220226
rect 453554 220170 453622 220226
rect 453678 220170 471250 220226
rect 471306 220170 471374 220226
rect 471430 220170 471498 220226
rect 471554 220170 471622 220226
rect 471678 220170 489250 220226
rect 489306 220170 489374 220226
rect 489430 220170 489498 220226
rect 489554 220170 489622 220226
rect 489678 220170 507250 220226
rect 507306 220170 507374 220226
rect 507430 220170 507498 220226
rect 507554 220170 507622 220226
rect 507678 220170 525250 220226
rect 525306 220170 525374 220226
rect 525430 220170 525498 220226
rect 525554 220170 525622 220226
rect 525678 220170 543250 220226
rect 543306 220170 543374 220226
rect 543430 220170 543498 220226
rect 543554 220170 543622 220226
rect 543678 220170 561250 220226
rect 561306 220170 561374 220226
rect 561430 220170 561498 220226
rect 561554 220170 561622 220226
rect 561678 220170 579250 220226
rect 579306 220170 579374 220226
rect 579430 220170 579498 220226
rect 579554 220170 579622 220226
rect 579678 220170 596496 220226
rect 596552 220170 596620 220226
rect 596676 220170 596744 220226
rect 596800 220170 596868 220226
rect 596924 220170 597980 220226
rect -1916 220102 597980 220170
rect -1916 220046 -860 220102
rect -804 220046 -736 220102
rect -680 220046 -612 220102
rect -556 220046 -488 220102
rect -432 220046 3250 220102
rect 3306 220046 3374 220102
rect 3430 220046 3498 220102
rect 3554 220046 3622 220102
rect 3678 220046 21250 220102
rect 21306 220046 21374 220102
rect 21430 220046 21498 220102
rect 21554 220046 21622 220102
rect 21678 220046 39250 220102
rect 39306 220046 39374 220102
rect 39430 220046 39498 220102
rect 39554 220046 39622 220102
rect 39678 220046 57250 220102
rect 57306 220046 57374 220102
rect 57430 220046 57498 220102
rect 57554 220046 57622 220102
rect 57678 220046 64518 220102
rect 64574 220046 64642 220102
rect 64698 220046 75250 220102
rect 75306 220046 75374 220102
rect 75430 220046 75498 220102
rect 75554 220046 75622 220102
rect 75678 220046 93250 220102
rect 93306 220046 93374 220102
rect 93430 220046 93498 220102
rect 93554 220046 93622 220102
rect 93678 220046 95238 220102
rect 95294 220046 95362 220102
rect 95418 220046 111250 220102
rect 111306 220046 111374 220102
rect 111430 220046 111498 220102
rect 111554 220046 111622 220102
rect 111678 220046 125958 220102
rect 126014 220046 126082 220102
rect 126138 220046 129250 220102
rect 129306 220046 129374 220102
rect 129430 220046 129498 220102
rect 129554 220046 129622 220102
rect 129678 220046 147250 220102
rect 147306 220046 147374 220102
rect 147430 220046 147498 220102
rect 147554 220046 147622 220102
rect 147678 220046 156678 220102
rect 156734 220046 156802 220102
rect 156858 220046 165250 220102
rect 165306 220046 165374 220102
rect 165430 220046 165498 220102
rect 165554 220046 165622 220102
rect 165678 220046 183250 220102
rect 183306 220046 183374 220102
rect 183430 220046 183498 220102
rect 183554 220046 183622 220102
rect 183678 220046 187398 220102
rect 187454 220046 187522 220102
rect 187578 220046 201250 220102
rect 201306 220046 201374 220102
rect 201430 220046 201498 220102
rect 201554 220046 201622 220102
rect 201678 220046 218118 220102
rect 218174 220046 218242 220102
rect 218298 220046 219250 220102
rect 219306 220046 219374 220102
rect 219430 220046 219498 220102
rect 219554 220046 219622 220102
rect 219678 220046 237250 220102
rect 237306 220046 237374 220102
rect 237430 220046 237498 220102
rect 237554 220046 237622 220102
rect 237678 220046 255250 220102
rect 255306 220046 255374 220102
rect 255430 220046 255498 220102
rect 255554 220046 255622 220102
rect 255678 220046 273250 220102
rect 273306 220046 273374 220102
rect 273430 220046 273498 220102
rect 273554 220046 273622 220102
rect 273678 220046 291250 220102
rect 291306 220046 291374 220102
rect 291430 220046 291498 220102
rect 291554 220046 291622 220102
rect 291678 220046 309250 220102
rect 309306 220046 309374 220102
rect 309430 220046 309498 220102
rect 309554 220046 309622 220102
rect 309678 220046 327250 220102
rect 327306 220046 327374 220102
rect 327430 220046 327498 220102
rect 327554 220046 327622 220102
rect 327678 220046 345250 220102
rect 345306 220046 345374 220102
rect 345430 220046 345498 220102
rect 345554 220046 345622 220102
rect 345678 220046 363250 220102
rect 363306 220046 363374 220102
rect 363430 220046 363498 220102
rect 363554 220046 363622 220102
rect 363678 220046 381250 220102
rect 381306 220046 381374 220102
rect 381430 220046 381498 220102
rect 381554 220046 381622 220102
rect 381678 220046 399250 220102
rect 399306 220046 399374 220102
rect 399430 220046 399498 220102
rect 399554 220046 399622 220102
rect 399678 220046 417250 220102
rect 417306 220046 417374 220102
rect 417430 220046 417498 220102
rect 417554 220046 417622 220102
rect 417678 220046 435250 220102
rect 435306 220046 435374 220102
rect 435430 220046 435498 220102
rect 435554 220046 435622 220102
rect 435678 220046 453250 220102
rect 453306 220046 453374 220102
rect 453430 220046 453498 220102
rect 453554 220046 453622 220102
rect 453678 220046 471250 220102
rect 471306 220046 471374 220102
rect 471430 220046 471498 220102
rect 471554 220046 471622 220102
rect 471678 220046 489250 220102
rect 489306 220046 489374 220102
rect 489430 220046 489498 220102
rect 489554 220046 489622 220102
rect 489678 220046 507250 220102
rect 507306 220046 507374 220102
rect 507430 220046 507498 220102
rect 507554 220046 507622 220102
rect 507678 220046 525250 220102
rect 525306 220046 525374 220102
rect 525430 220046 525498 220102
rect 525554 220046 525622 220102
rect 525678 220046 543250 220102
rect 543306 220046 543374 220102
rect 543430 220046 543498 220102
rect 543554 220046 543622 220102
rect 543678 220046 561250 220102
rect 561306 220046 561374 220102
rect 561430 220046 561498 220102
rect 561554 220046 561622 220102
rect 561678 220046 579250 220102
rect 579306 220046 579374 220102
rect 579430 220046 579498 220102
rect 579554 220046 579622 220102
rect 579678 220046 596496 220102
rect 596552 220046 596620 220102
rect 596676 220046 596744 220102
rect 596800 220046 596868 220102
rect 596924 220046 597980 220102
rect -1916 219978 597980 220046
rect -1916 219922 -860 219978
rect -804 219922 -736 219978
rect -680 219922 -612 219978
rect -556 219922 -488 219978
rect -432 219922 3250 219978
rect 3306 219922 3374 219978
rect 3430 219922 3498 219978
rect 3554 219922 3622 219978
rect 3678 219922 21250 219978
rect 21306 219922 21374 219978
rect 21430 219922 21498 219978
rect 21554 219922 21622 219978
rect 21678 219922 39250 219978
rect 39306 219922 39374 219978
rect 39430 219922 39498 219978
rect 39554 219922 39622 219978
rect 39678 219922 57250 219978
rect 57306 219922 57374 219978
rect 57430 219922 57498 219978
rect 57554 219922 57622 219978
rect 57678 219922 64518 219978
rect 64574 219922 64642 219978
rect 64698 219922 75250 219978
rect 75306 219922 75374 219978
rect 75430 219922 75498 219978
rect 75554 219922 75622 219978
rect 75678 219922 93250 219978
rect 93306 219922 93374 219978
rect 93430 219922 93498 219978
rect 93554 219922 93622 219978
rect 93678 219922 95238 219978
rect 95294 219922 95362 219978
rect 95418 219922 111250 219978
rect 111306 219922 111374 219978
rect 111430 219922 111498 219978
rect 111554 219922 111622 219978
rect 111678 219922 125958 219978
rect 126014 219922 126082 219978
rect 126138 219922 129250 219978
rect 129306 219922 129374 219978
rect 129430 219922 129498 219978
rect 129554 219922 129622 219978
rect 129678 219922 147250 219978
rect 147306 219922 147374 219978
rect 147430 219922 147498 219978
rect 147554 219922 147622 219978
rect 147678 219922 156678 219978
rect 156734 219922 156802 219978
rect 156858 219922 165250 219978
rect 165306 219922 165374 219978
rect 165430 219922 165498 219978
rect 165554 219922 165622 219978
rect 165678 219922 183250 219978
rect 183306 219922 183374 219978
rect 183430 219922 183498 219978
rect 183554 219922 183622 219978
rect 183678 219922 187398 219978
rect 187454 219922 187522 219978
rect 187578 219922 201250 219978
rect 201306 219922 201374 219978
rect 201430 219922 201498 219978
rect 201554 219922 201622 219978
rect 201678 219922 218118 219978
rect 218174 219922 218242 219978
rect 218298 219922 219250 219978
rect 219306 219922 219374 219978
rect 219430 219922 219498 219978
rect 219554 219922 219622 219978
rect 219678 219922 237250 219978
rect 237306 219922 237374 219978
rect 237430 219922 237498 219978
rect 237554 219922 237622 219978
rect 237678 219922 255250 219978
rect 255306 219922 255374 219978
rect 255430 219922 255498 219978
rect 255554 219922 255622 219978
rect 255678 219922 273250 219978
rect 273306 219922 273374 219978
rect 273430 219922 273498 219978
rect 273554 219922 273622 219978
rect 273678 219922 291250 219978
rect 291306 219922 291374 219978
rect 291430 219922 291498 219978
rect 291554 219922 291622 219978
rect 291678 219922 309250 219978
rect 309306 219922 309374 219978
rect 309430 219922 309498 219978
rect 309554 219922 309622 219978
rect 309678 219922 327250 219978
rect 327306 219922 327374 219978
rect 327430 219922 327498 219978
rect 327554 219922 327622 219978
rect 327678 219922 345250 219978
rect 345306 219922 345374 219978
rect 345430 219922 345498 219978
rect 345554 219922 345622 219978
rect 345678 219922 363250 219978
rect 363306 219922 363374 219978
rect 363430 219922 363498 219978
rect 363554 219922 363622 219978
rect 363678 219922 381250 219978
rect 381306 219922 381374 219978
rect 381430 219922 381498 219978
rect 381554 219922 381622 219978
rect 381678 219922 399250 219978
rect 399306 219922 399374 219978
rect 399430 219922 399498 219978
rect 399554 219922 399622 219978
rect 399678 219922 417250 219978
rect 417306 219922 417374 219978
rect 417430 219922 417498 219978
rect 417554 219922 417622 219978
rect 417678 219922 435250 219978
rect 435306 219922 435374 219978
rect 435430 219922 435498 219978
rect 435554 219922 435622 219978
rect 435678 219922 453250 219978
rect 453306 219922 453374 219978
rect 453430 219922 453498 219978
rect 453554 219922 453622 219978
rect 453678 219922 471250 219978
rect 471306 219922 471374 219978
rect 471430 219922 471498 219978
rect 471554 219922 471622 219978
rect 471678 219922 489250 219978
rect 489306 219922 489374 219978
rect 489430 219922 489498 219978
rect 489554 219922 489622 219978
rect 489678 219922 507250 219978
rect 507306 219922 507374 219978
rect 507430 219922 507498 219978
rect 507554 219922 507622 219978
rect 507678 219922 525250 219978
rect 525306 219922 525374 219978
rect 525430 219922 525498 219978
rect 525554 219922 525622 219978
rect 525678 219922 543250 219978
rect 543306 219922 543374 219978
rect 543430 219922 543498 219978
rect 543554 219922 543622 219978
rect 543678 219922 561250 219978
rect 561306 219922 561374 219978
rect 561430 219922 561498 219978
rect 561554 219922 561622 219978
rect 561678 219922 579250 219978
rect 579306 219922 579374 219978
rect 579430 219922 579498 219978
rect 579554 219922 579622 219978
rect 579678 219922 596496 219978
rect 596552 219922 596620 219978
rect 596676 219922 596744 219978
rect 596800 219922 596868 219978
rect 596924 219922 597980 219978
rect -1916 219826 597980 219922
rect -1916 208412 597980 208446
rect -1916 208356 364022 208412
rect 364078 208356 364146 208412
rect 364202 208356 364270 208412
rect 364326 208356 364394 208412
rect 364450 208356 364518 208412
rect 364574 208356 364642 208412
rect 364698 208356 364766 208412
rect 364822 208356 364890 208412
rect 364946 208356 365014 208412
rect 365070 208356 365138 208412
rect 365194 208356 384022 208412
rect 384078 208356 384146 208412
rect 384202 208356 384270 208412
rect 384326 208356 384394 208412
rect 384450 208356 384518 208412
rect 384574 208356 384642 208412
rect 384698 208356 384766 208412
rect 384822 208356 384890 208412
rect 384946 208356 385014 208412
rect 385070 208356 385138 208412
rect 385194 208356 404022 208412
rect 404078 208356 404146 208412
rect 404202 208356 404270 208412
rect 404326 208356 404394 208412
rect 404450 208356 404518 208412
rect 404574 208356 404642 208412
rect 404698 208356 404766 208412
rect 404822 208356 404890 208412
rect 404946 208356 405014 208412
rect 405070 208356 405138 208412
rect 405194 208356 424022 208412
rect 424078 208356 424146 208412
rect 424202 208356 424270 208412
rect 424326 208356 424394 208412
rect 424450 208356 424518 208412
rect 424574 208356 424642 208412
rect 424698 208356 424766 208412
rect 424822 208356 424890 208412
rect 424946 208356 425014 208412
rect 425070 208356 425138 208412
rect 425194 208356 444022 208412
rect 444078 208356 444146 208412
rect 444202 208356 444270 208412
rect 444326 208356 444394 208412
rect 444450 208356 444518 208412
rect 444574 208356 444642 208412
rect 444698 208356 444766 208412
rect 444822 208356 444890 208412
rect 444946 208356 445014 208412
rect 445070 208356 445138 208412
rect 445194 208356 464022 208412
rect 464078 208356 464146 208412
rect 464202 208356 464270 208412
rect 464326 208356 464394 208412
rect 464450 208356 464518 208412
rect 464574 208356 464642 208412
rect 464698 208356 464766 208412
rect 464822 208356 464890 208412
rect 464946 208356 465014 208412
rect 465070 208356 465138 208412
rect 465194 208356 484022 208412
rect 484078 208356 484146 208412
rect 484202 208356 484270 208412
rect 484326 208356 484394 208412
rect 484450 208356 484518 208412
rect 484574 208356 484642 208412
rect 484698 208356 484766 208412
rect 484822 208356 484890 208412
rect 484946 208356 485014 208412
rect 485070 208356 485138 208412
rect 485194 208356 504022 208412
rect 504078 208356 504146 208412
rect 504202 208356 504270 208412
rect 504326 208356 504394 208412
rect 504450 208356 504518 208412
rect 504574 208356 504642 208412
rect 504698 208356 504766 208412
rect 504822 208356 504890 208412
rect 504946 208356 505014 208412
rect 505070 208356 505138 208412
rect 505194 208356 524022 208412
rect 524078 208356 524146 208412
rect 524202 208356 524270 208412
rect 524326 208356 524394 208412
rect 524450 208356 524518 208412
rect 524574 208356 524642 208412
rect 524698 208356 524766 208412
rect 524822 208356 524890 208412
rect 524946 208356 525014 208412
rect 525070 208356 525138 208412
rect 525194 208356 544022 208412
rect 544078 208356 544146 208412
rect 544202 208356 544270 208412
rect 544326 208356 544394 208412
rect 544450 208356 544518 208412
rect 544574 208356 544642 208412
rect 544698 208356 544766 208412
rect 544822 208356 544890 208412
rect 544946 208356 545014 208412
rect 545070 208356 545138 208412
rect 545194 208356 597980 208412
rect -1916 208350 597980 208356
rect -1916 208294 -1820 208350
rect -1764 208294 -1696 208350
rect -1640 208294 -1572 208350
rect -1516 208294 -1448 208350
rect -1392 208294 6970 208350
rect 7026 208294 7094 208350
rect 7150 208294 7218 208350
rect 7274 208294 7342 208350
rect 7398 208294 24970 208350
rect 25026 208294 25094 208350
rect 25150 208294 25218 208350
rect 25274 208294 25342 208350
rect 25398 208294 42970 208350
rect 43026 208294 43094 208350
rect 43150 208294 43218 208350
rect 43274 208294 43342 208350
rect 43398 208294 79878 208350
rect 79934 208294 80002 208350
rect 80058 208294 110598 208350
rect 110654 208294 110722 208350
rect 110778 208294 141318 208350
rect 141374 208294 141442 208350
rect 141498 208294 172038 208350
rect 172094 208294 172162 208350
rect 172218 208294 202758 208350
rect 202814 208294 202882 208350
rect 202938 208294 233478 208350
rect 233534 208294 233602 208350
rect 233658 208294 240970 208350
rect 241026 208294 241094 208350
rect 241150 208294 241218 208350
rect 241274 208294 241342 208350
rect 241398 208294 258970 208350
rect 259026 208294 259094 208350
rect 259150 208294 259218 208350
rect 259274 208294 259342 208350
rect 259398 208294 276970 208350
rect 277026 208294 277094 208350
rect 277150 208294 277218 208350
rect 277274 208294 277342 208350
rect 277398 208294 294970 208350
rect 295026 208294 295094 208350
rect 295150 208294 295218 208350
rect 295274 208294 295342 208350
rect 295398 208294 312970 208350
rect 313026 208294 313094 208350
rect 313150 208294 313218 208350
rect 313274 208294 313342 208350
rect 313398 208294 330970 208350
rect 331026 208294 331094 208350
rect 331150 208294 331218 208350
rect 331274 208294 331342 208350
rect 331398 208294 348970 208350
rect 349026 208294 349094 208350
rect 349150 208294 349218 208350
rect 349274 208294 349342 208350
rect 349398 208294 564970 208350
rect 565026 208294 565094 208350
rect 565150 208294 565218 208350
rect 565274 208294 565342 208350
rect 565398 208294 582970 208350
rect 583026 208294 583094 208350
rect 583150 208294 583218 208350
rect 583274 208294 583342 208350
rect 583398 208294 597456 208350
rect 597512 208294 597580 208350
rect 597636 208294 597704 208350
rect 597760 208294 597828 208350
rect 597884 208294 597980 208350
rect -1916 208288 597980 208294
rect -1916 208232 364022 208288
rect 364078 208232 364146 208288
rect 364202 208232 364270 208288
rect 364326 208232 364394 208288
rect 364450 208232 364518 208288
rect 364574 208232 364642 208288
rect 364698 208232 364766 208288
rect 364822 208232 364890 208288
rect 364946 208232 365014 208288
rect 365070 208232 365138 208288
rect 365194 208232 384022 208288
rect 384078 208232 384146 208288
rect 384202 208232 384270 208288
rect 384326 208232 384394 208288
rect 384450 208232 384518 208288
rect 384574 208232 384642 208288
rect 384698 208232 384766 208288
rect 384822 208232 384890 208288
rect 384946 208232 385014 208288
rect 385070 208232 385138 208288
rect 385194 208232 404022 208288
rect 404078 208232 404146 208288
rect 404202 208232 404270 208288
rect 404326 208232 404394 208288
rect 404450 208232 404518 208288
rect 404574 208232 404642 208288
rect 404698 208232 404766 208288
rect 404822 208232 404890 208288
rect 404946 208232 405014 208288
rect 405070 208232 405138 208288
rect 405194 208232 424022 208288
rect 424078 208232 424146 208288
rect 424202 208232 424270 208288
rect 424326 208232 424394 208288
rect 424450 208232 424518 208288
rect 424574 208232 424642 208288
rect 424698 208232 424766 208288
rect 424822 208232 424890 208288
rect 424946 208232 425014 208288
rect 425070 208232 425138 208288
rect 425194 208232 444022 208288
rect 444078 208232 444146 208288
rect 444202 208232 444270 208288
rect 444326 208232 444394 208288
rect 444450 208232 444518 208288
rect 444574 208232 444642 208288
rect 444698 208232 444766 208288
rect 444822 208232 444890 208288
rect 444946 208232 445014 208288
rect 445070 208232 445138 208288
rect 445194 208232 464022 208288
rect 464078 208232 464146 208288
rect 464202 208232 464270 208288
rect 464326 208232 464394 208288
rect 464450 208232 464518 208288
rect 464574 208232 464642 208288
rect 464698 208232 464766 208288
rect 464822 208232 464890 208288
rect 464946 208232 465014 208288
rect 465070 208232 465138 208288
rect 465194 208232 484022 208288
rect 484078 208232 484146 208288
rect 484202 208232 484270 208288
rect 484326 208232 484394 208288
rect 484450 208232 484518 208288
rect 484574 208232 484642 208288
rect 484698 208232 484766 208288
rect 484822 208232 484890 208288
rect 484946 208232 485014 208288
rect 485070 208232 485138 208288
rect 485194 208232 504022 208288
rect 504078 208232 504146 208288
rect 504202 208232 504270 208288
rect 504326 208232 504394 208288
rect 504450 208232 504518 208288
rect 504574 208232 504642 208288
rect 504698 208232 504766 208288
rect 504822 208232 504890 208288
rect 504946 208232 505014 208288
rect 505070 208232 505138 208288
rect 505194 208232 524022 208288
rect 524078 208232 524146 208288
rect 524202 208232 524270 208288
rect 524326 208232 524394 208288
rect 524450 208232 524518 208288
rect 524574 208232 524642 208288
rect 524698 208232 524766 208288
rect 524822 208232 524890 208288
rect 524946 208232 525014 208288
rect 525070 208232 525138 208288
rect 525194 208232 544022 208288
rect 544078 208232 544146 208288
rect 544202 208232 544270 208288
rect 544326 208232 544394 208288
rect 544450 208232 544518 208288
rect 544574 208232 544642 208288
rect 544698 208232 544766 208288
rect 544822 208232 544890 208288
rect 544946 208232 545014 208288
rect 545070 208232 545138 208288
rect 545194 208232 597980 208288
rect -1916 208226 597980 208232
rect -1916 208170 -1820 208226
rect -1764 208170 -1696 208226
rect -1640 208170 -1572 208226
rect -1516 208170 -1448 208226
rect -1392 208170 6970 208226
rect 7026 208170 7094 208226
rect 7150 208170 7218 208226
rect 7274 208170 7342 208226
rect 7398 208170 24970 208226
rect 25026 208170 25094 208226
rect 25150 208170 25218 208226
rect 25274 208170 25342 208226
rect 25398 208170 42970 208226
rect 43026 208170 43094 208226
rect 43150 208170 43218 208226
rect 43274 208170 43342 208226
rect 43398 208170 79878 208226
rect 79934 208170 80002 208226
rect 80058 208170 110598 208226
rect 110654 208170 110722 208226
rect 110778 208170 141318 208226
rect 141374 208170 141442 208226
rect 141498 208170 172038 208226
rect 172094 208170 172162 208226
rect 172218 208170 202758 208226
rect 202814 208170 202882 208226
rect 202938 208170 233478 208226
rect 233534 208170 233602 208226
rect 233658 208170 240970 208226
rect 241026 208170 241094 208226
rect 241150 208170 241218 208226
rect 241274 208170 241342 208226
rect 241398 208170 258970 208226
rect 259026 208170 259094 208226
rect 259150 208170 259218 208226
rect 259274 208170 259342 208226
rect 259398 208170 276970 208226
rect 277026 208170 277094 208226
rect 277150 208170 277218 208226
rect 277274 208170 277342 208226
rect 277398 208170 294970 208226
rect 295026 208170 295094 208226
rect 295150 208170 295218 208226
rect 295274 208170 295342 208226
rect 295398 208170 312970 208226
rect 313026 208170 313094 208226
rect 313150 208170 313218 208226
rect 313274 208170 313342 208226
rect 313398 208170 330970 208226
rect 331026 208170 331094 208226
rect 331150 208170 331218 208226
rect 331274 208170 331342 208226
rect 331398 208170 348970 208226
rect 349026 208170 349094 208226
rect 349150 208170 349218 208226
rect 349274 208170 349342 208226
rect 349398 208170 564970 208226
rect 565026 208170 565094 208226
rect 565150 208170 565218 208226
rect 565274 208170 565342 208226
rect 565398 208170 582970 208226
rect 583026 208170 583094 208226
rect 583150 208170 583218 208226
rect 583274 208170 583342 208226
rect 583398 208170 597456 208226
rect 597512 208170 597580 208226
rect 597636 208170 597704 208226
rect 597760 208170 597828 208226
rect 597884 208170 597980 208226
rect -1916 208164 597980 208170
rect -1916 208108 364022 208164
rect 364078 208108 364146 208164
rect 364202 208108 364270 208164
rect 364326 208108 364394 208164
rect 364450 208108 364518 208164
rect 364574 208108 364642 208164
rect 364698 208108 364766 208164
rect 364822 208108 364890 208164
rect 364946 208108 365014 208164
rect 365070 208108 365138 208164
rect 365194 208108 384022 208164
rect 384078 208108 384146 208164
rect 384202 208108 384270 208164
rect 384326 208108 384394 208164
rect 384450 208108 384518 208164
rect 384574 208108 384642 208164
rect 384698 208108 384766 208164
rect 384822 208108 384890 208164
rect 384946 208108 385014 208164
rect 385070 208108 385138 208164
rect 385194 208108 404022 208164
rect 404078 208108 404146 208164
rect 404202 208108 404270 208164
rect 404326 208108 404394 208164
rect 404450 208108 404518 208164
rect 404574 208108 404642 208164
rect 404698 208108 404766 208164
rect 404822 208108 404890 208164
rect 404946 208108 405014 208164
rect 405070 208108 405138 208164
rect 405194 208108 424022 208164
rect 424078 208108 424146 208164
rect 424202 208108 424270 208164
rect 424326 208108 424394 208164
rect 424450 208108 424518 208164
rect 424574 208108 424642 208164
rect 424698 208108 424766 208164
rect 424822 208108 424890 208164
rect 424946 208108 425014 208164
rect 425070 208108 425138 208164
rect 425194 208108 444022 208164
rect 444078 208108 444146 208164
rect 444202 208108 444270 208164
rect 444326 208108 444394 208164
rect 444450 208108 444518 208164
rect 444574 208108 444642 208164
rect 444698 208108 444766 208164
rect 444822 208108 444890 208164
rect 444946 208108 445014 208164
rect 445070 208108 445138 208164
rect 445194 208108 464022 208164
rect 464078 208108 464146 208164
rect 464202 208108 464270 208164
rect 464326 208108 464394 208164
rect 464450 208108 464518 208164
rect 464574 208108 464642 208164
rect 464698 208108 464766 208164
rect 464822 208108 464890 208164
rect 464946 208108 465014 208164
rect 465070 208108 465138 208164
rect 465194 208108 484022 208164
rect 484078 208108 484146 208164
rect 484202 208108 484270 208164
rect 484326 208108 484394 208164
rect 484450 208108 484518 208164
rect 484574 208108 484642 208164
rect 484698 208108 484766 208164
rect 484822 208108 484890 208164
rect 484946 208108 485014 208164
rect 485070 208108 485138 208164
rect 485194 208108 504022 208164
rect 504078 208108 504146 208164
rect 504202 208108 504270 208164
rect 504326 208108 504394 208164
rect 504450 208108 504518 208164
rect 504574 208108 504642 208164
rect 504698 208108 504766 208164
rect 504822 208108 504890 208164
rect 504946 208108 505014 208164
rect 505070 208108 505138 208164
rect 505194 208108 524022 208164
rect 524078 208108 524146 208164
rect 524202 208108 524270 208164
rect 524326 208108 524394 208164
rect 524450 208108 524518 208164
rect 524574 208108 524642 208164
rect 524698 208108 524766 208164
rect 524822 208108 524890 208164
rect 524946 208108 525014 208164
rect 525070 208108 525138 208164
rect 525194 208108 544022 208164
rect 544078 208108 544146 208164
rect 544202 208108 544270 208164
rect 544326 208108 544394 208164
rect 544450 208108 544518 208164
rect 544574 208108 544642 208164
rect 544698 208108 544766 208164
rect 544822 208108 544890 208164
rect 544946 208108 545014 208164
rect 545070 208108 545138 208164
rect 545194 208108 597980 208164
rect -1916 208102 597980 208108
rect -1916 208046 -1820 208102
rect -1764 208046 -1696 208102
rect -1640 208046 -1572 208102
rect -1516 208046 -1448 208102
rect -1392 208046 6970 208102
rect 7026 208046 7094 208102
rect 7150 208046 7218 208102
rect 7274 208046 7342 208102
rect 7398 208046 24970 208102
rect 25026 208046 25094 208102
rect 25150 208046 25218 208102
rect 25274 208046 25342 208102
rect 25398 208046 42970 208102
rect 43026 208046 43094 208102
rect 43150 208046 43218 208102
rect 43274 208046 43342 208102
rect 43398 208046 79878 208102
rect 79934 208046 80002 208102
rect 80058 208046 110598 208102
rect 110654 208046 110722 208102
rect 110778 208046 141318 208102
rect 141374 208046 141442 208102
rect 141498 208046 172038 208102
rect 172094 208046 172162 208102
rect 172218 208046 202758 208102
rect 202814 208046 202882 208102
rect 202938 208046 233478 208102
rect 233534 208046 233602 208102
rect 233658 208046 240970 208102
rect 241026 208046 241094 208102
rect 241150 208046 241218 208102
rect 241274 208046 241342 208102
rect 241398 208046 258970 208102
rect 259026 208046 259094 208102
rect 259150 208046 259218 208102
rect 259274 208046 259342 208102
rect 259398 208046 276970 208102
rect 277026 208046 277094 208102
rect 277150 208046 277218 208102
rect 277274 208046 277342 208102
rect 277398 208046 294970 208102
rect 295026 208046 295094 208102
rect 295150 208046 295218 208102
rect 295274 208046 295342 208102
rect 295398 208046 312970 208102
rect 313026 208046 313094 208102
rect 313150 208046 313218 208102
rect 313274 208046 313342 208102
rect 313398 208046 330970 208102
rect 331026 208046 331094 208102
rect 331150 208046 331218 208102
rect 331274 208046 331342 208102
rect 331398 208046 348970 208102
rect 349026 208046 349094 208102
rect 349150 208046 349218 208102
rect 349274 208046 349342 208102
rect 349398 208046 564970 208102
rect 565026 208046 565094 208102
rect 565150 208046 565218 208102
rect 565274 208046 565342 208102
rect 565398 208046 582970 208102
rect 583026 208046 583094 208102
rect 583150 208046 583218 208102
rect 583274 208046 583342 208102
rect 583398 208046 597456 208102
rect 597512 208046 597580 208102
rect 597636 208046 597704 208102
rect 597760 208046 597828 208102
rect 597884 208046 597980 208102
rect -1916 208040 597980 208046
rect -1916 207984 364022 208040
rect 364078 207984 364146 208040
rect 364202 207984 364270 208040
rect 364326 207984 364394 208040
rect 364450 207984 364518 208040
rect 364574 207984 364642 208040
rect 364698 207984 364766 208040
rect 364822 207984 364890 208040
rect 364946 207984 365014 208040
rect 365070 207984 365138 208040
rect 365194 207984 384022 208040
rect 384078 207984 384146 208040
rect 384202 207984 384270 208040
rect 384326 207984 384394 208040
rect 384450 207984 384518 208040
rect 384574 207984 384642 208040
rect 384698 207984 384766 208040
rect 384822 207984 384890 208040
rect 384946 207984 385014 208040
rect 385070 207984 385138 208040
rect 385194 207984 404022 208040
rect 404078 207984 404146 208040
rect 404202 207984 404270 208040
rect 404326 207984 404394 208040
rect 404450 207984 404518 208040
rect 404574 207984 404642 208040
rect 404698 207984 404766 208040
rect 404822 207984 404890 208040
rect 404946 207984 405014 208040
rect 405070 207984 405138 208040
rect 405194 207984 424022 208040
rect 424078 207984 424146 208040
rect 424202 207984 424270 208040
rect 424326 207984 424394 208040
rect 424450 207984 424518 208040
rect 424574 207984 424642 208040
rect 424698 207984 424766 208040
rect 424822 207984 424890 208040
rect 424946 207984 425014 208040
rect 425070 207984 425138 208040
rect 425194 207984 444022 208040
rect 444078 207984 444146 208040
rect 444202 207984 444270 208040
rect 444326 207984 444394 208040
rect 444450 207984 444518 208040
rect 444574 207984 444642 208040
rect 444698 207984 444766 208040
rect 444822 207984 444890 208040
rect 444946 207984 445014 208040
rect 445070 207984 445138 208040
rect 445194 207984 464022 208040
rect 464078 207984 464146 208040
rect 464202 207984 464270 208040
rect 464326 207984 464394 208040
rect 464450 207984 464518 208040
rect 464574 207984 464642 208040
rect 464698 207984 464766 208040
rect 464822 207984 464890 208040
rect 464946 207984 465014 208040
rect 465070 207984 465138 208040
rect 465194 207984 484022 208040
rect 484078 207984 484146 208040
rect 484202 207984 484270 208040
rect 484326 207984 484394 208040
rect 484450 207984 484518 208040
rect 484574 207984 484642 208040
rect 484698 207984 484766 208040
rect 484822 207984 484890 208040
rect 484946 207984 485014 208040
rect 485070 207984 485138 208040
rect 485194 207984 504022 208040
rect 504078 207984 504146 208040
rect 504202 207984 504270 208040
rect 504326 207984 504394 208040
rect 504450 207984 504518 208040
rect 504574 207984 504642 208040
rect 504698 207984 504766 208040
rect 504822 207984 504890 208040
rect 504946 207984 505014 208040
rect 505070 207984 505138 208040
rect 505194 207984 524022 208040
rect 524078 207984 524146 208040
rect 524202 207984 524270 208040
rect 524326 207984 524394 208040
rect 524450 207984 524518 208040
rect 524574 207984 524642 208040
rect 524698 207984 524766 208040
rect 524822 207984 524890 208040
rect 524946 207984 525014 208040
rect 525070 207984 525138 208040
rect 525194 207984 544022 208040
rect 544078 207984 544146 208040
rect 544202 207984 544270 208040
rect 544326 207984 544394 208040
rect 544450 207984 544518 208040
rect 544574 207984 544642 208040
rect 544698 207984 544766 208040
rect 544822 207984 544890 208040
rect 544946 207984 545014 208040
rect 545070 207984 545138 208040
rect 545194 207984 597980 208040
rect -1916 207978 597980 207984
rect -1916 207922 -1820 207978
rect -1764 207922 -1696 207978
rect -1640 207922 -1572 207978
rect -1516 207922 -1448 207978
rect -1392 207922 6970 207978
rect 7026 207922 7094 207978
rect 7150 207922 7218 207978
rect 7274 207922 7342 207978
rect 7398 207922 24970 207978
rect 25026 207922 25094 207978
rect 25150 207922 25218 207978
rect 25274 207922 25342 207978
rect 25398 207922 42970 207978
rect 43026 207922 43094 207978
rect 43150 207922 43218 207978
rect 43274 207922 43342 207978
rect 43398 207922 79878 207978
rect 79934 207922 80002 207978
rect 80058 207922 110598 207978
rect 110654 207922 110722 207978
rect 110778 207922 141318 207978
rect 141374 207922 141442 207978
rect 141498 207922 172038 207978
rect 172094 207922 172162 207978
rect 172218 207922 202758 207978
rect 202814 207922 202882 207978
rect 202938 207922 233478 207978
rect 233534 207922 233602 207978
rect 233658 207922 240970 207978
rect 241026 207922 241094 207978
rect 241150 207922 241218 207978
rect 241274 207922 241342 207978
rect 241398 207922 258970 207978
rect 259026 207922 259094 207978
rect 259150 207922 259218 207978
rect 259274 207922 259342 207978
rect 259398 207922 276970 207978
rect 277026 207922 277094 207978
rect 277150 207922 277218 207978
rect 277274 207922 277342 207978
rect 277398 207922 294970 207978
rect 295026 207922 295094 207978
rect 295150 207922 295218 207978
rect 295274 207922 295342 207978
rect 295398 207922 312970 207978
rect 313026 207922 313094 207978
rect 313150 207922 313218 207978
rect 313274 207922 313342 207978
rect 313398 207922 330970 207978
rect 331026 207922 331094 207978
rect 331150 207922 331218 207978
rect 331274 207922 331342 207978
rect 331398 207922 348970 207978
rect 349026 207922 349094 207978
rect 349150 207922 349218 207978
rect 349274 207922 349342 207978
rect 349398 207922 564970 207978
rect 565026 207922 565094 207978
rect 565150 207922 565218 207978
rect 565274 207922 565342 207978
rect 565398 207922 582970 207978
rect 583026 207922 583094 207978
rect 583150 207922 583218 207978
rect 583274 207922 583342 207978
rect 583398 207922 597456 207978
rect 597512 207922 597580 207978
rect 597636 207922 597704 207978
rect 597760 207922 597828 207978
rect 597884 207922 597980 207978
rect -1916 207916 597980 207922
rect -1916 207860 364022 207916
rect 364078 207860 364146 207916
rect 364202 207860 364270 207916
rect 364326 207860 364394 207916
rect 364450 207860 364518 207916
rect 364574 207860 364642 207916
rect 364698 207860 364766 207916
rect 364822 207860 364890 207916
rect 364946 207860 365014 207916
rect 365070 207860 365138 207916
rect 365194 207860 384022 207916
rect 384078 207860 384146 207916
rect 384202 207860 384270 207916
rect 384326 207860 384394 207916
rect 384450 207860 384518 207916
rect 384574 207860 384642 207916
rect 384698 207860 384766 207916
rect 384822 207860 384890 207916
rect 384946 207860 385014 207916
rect 385070 207860 385138 207916
rect 385194 207860 404022 207916
rect 404078 207860 404146 207916
rect 404202 207860 404270 207916
rect 404326 207860 404394 207916
rect 404450 207860 404518 207916
rect 404574 207860 404642 207916
rect 404698 207860 404766 207916
rect 404822 207860 404890 207916
rect 404946 207860 405014 207916
rect 405070 207860 405138 207916
rect 405194 207860 424022 207916
rect 424078 207860 424146 207916
rect 424202 207860 424270 207916
rect 424326 207860 424394 207916
rect 424450 207860 424518 207916
rect 424574 207860 424642 207916
rect 424698 207860 424766 207916
rect 424822 207860 424890 207916
rect 424946 207860 425014 207916
rect 425070 207860 425138 207916
rect 425194 207860 444022 207916
rect 444078 207860 444146 207916
rect 444202 207860 444270 207916
rect 444326 207860 444394 207916
rect 444450 207860 444518 207916
rect 444574 207860 444642 207916
rect 444698 207860 444766 207916
rect 444822 207860 444890 207916
rect 444946 207860 445014 207916
rect 445070 207860 445138 207916
rect 445194 207860 464022 207916
rect 464078 207860 464146 207916
rect 464202 207860 464270 207916
rect 464326 207860 464394 207916
rect 464450 207860 464518 207916
rect 464574 207860 464642 207916
rect 464698 207860 464766 207916
rect 464822 207860 464890 207916
rect 464946 207860 465014 207916
rect 465070 207860 465138 207916
rect 465194 207860 484022 207916
rect 484078 207860 484146 207916
rect 484202 207860 484270 207916
rect 484326 207860 484394 207916
rect 484450 207860 484518 207916
rect 484574 207860 484642 207916
rect 484698 207860 484766 207916
rect 484822 207860 484890 207916
rect 484946 207860 485014 207916
rect 485070 207860 485138 207916
rect 485194 207860 504022 207916
rect 504078 207860 504146 207916
rect 504202 207860 504270 207916
rect 504326 207860 504394 207916
rect 504450 207860 504518 207916
rect 504574 207860 504642 207916
rect 504698 207860 504766 207916
rect 504822 207860 504890 207916
rect 504946 207860 505014 207916
rect 505070 207860 505138 207916
rect 505194 207860 524022 207916
rect 524078 207860 524146 207916
rect 524202 207860 524270 207916
rect 524326 207860 524394 207916
rect 524450 207860 524518 207916
rect 524574 207860 524642 207916
rect 524698 207860 524766 207916
rect 524822 207860 524890 207916
rect 524946 207860 525014 207916
rect 525070 207860 525138 207916
rect 525194 207860 544022 207916
rect 544078 207860 544146 207916
rect 544202 207860 544270 207916
rect 544326 207860 544394 207916
rect 544450 207860 544518 207916
rect 544574 207860 544642 207916
rect 544698 207860 544766 207916
rect 544822 207860 544890 207916
rect 544946 207860 545014 207916
rect 545070 207860 545138 207916
rect 545194 207860 597980 207916
rect -1916 207826 597980 207860
rect -1916 202412 597980 202446
rect -1916 202356 354022 202412
rect 354078 202356 354146 202412
rect 354202 202356 354270 202412
rect 354326 202356 354394 202412
rect 354450 202356 354518 202412
rect 354574 202356 354642 202412
rect 354698 202356 354766 202412
rect 354822 202356 354890 202412
rect 354946 202356 355014 202412
rect 355070 202356 355138 202412
rect 355194 202356 374022 202412
rect 374078 202356 374146 202412
rect 374202 202356 374270 202412
rect 374326 202356 374394 202412
rect 374450 202356 374518 202412
rect 374574 202356 374642 202412
rect 374698 202356 374766 202412
rect 374822 202356 374890 202412
rect 374946 202356 375014 202412
rect 375070 202356 375138 202412
rect 375194 202356 394022 202412
rect 394078 202356 394146 202412
rect 394202 202356 394270 202412
rect 394326 202356 394394 202412
rect 394450 202356 394518 202412
rect 394574 202356 394642 202412
rect 394698 202356 394766 202412
rect 394822 202356 394890 202412
rect 394946 202356 395014 202412
rect 395070 202356 395138 202412
rect 395194 202356 414022 202412
rect 414078 202356 414146 202412
rect 414202 202356 414270 202412
rect 414326 202356 414394 202412
rect 414450 202356 414518 202412
rect 414574 202356 414642 202412
rect 414698 202356 414766 202412
rect 414822 202356 414890 202412
rect 414946 202356 415014 202412
rect 415070 202356 415138 202412
rect 415194 202356 434022 202412
rect 434078 202356 434146 202412
rect 434202 202356 434270 202412
rect 434326 202356 434394 202412
rect 434450 202356 434518 202412
rect 434574 202356 434642 202412
rect 434698 202356 434766 202412
rect 434822 202356 434890 202412
rect 434946 202356 435014 202412
rect 435070 202356 435138 202412
rect 435194 202356 454022 202412
rect 454078 202356 454146 202412
rect 454202 202356 454270 202412
rect 454326 202356 454394 202412
rect 454450 202356 454518 202412
rect 454574 202356 454642 202412
rect 454698 202356 454766 202412
rect 454822 202356 454890 202412
rect 454946 202356 455014 202412
rect 455070 202356 455138 202412
rect 455194 202356 474022 202412
rect 474078 202356 474146 202412
rect 474202 202356 474270 202412
rect 474326 202356 474394 202412
rect 474450 202356 474518 202412
rect 474574 202356 474642 202412
rect 474698 202356 474766 202412
rect 474822 202356 474890 202412
rect 474946 202356 475014 202412
rect 475070 202356 475138 202412
rect 475194 202356 494022 202412
rect 494078 202356 494146 202412
rect 494202 202356 494270 202412
rect 494326 202356 494394 202412
rect 494450 202356 494518 202412
rect 494574 202356 494642 202412
rect 494698 202356 494766 202412
rect 494822 202356 494890 202412
rect 494946 202356 495014 202412
rect 495070 202356 495138 202412
rect 495194 202356 514022 202412
rect 514078 202356 514146 202412
rect 514202 202356 514270 202412
rect 514326 202356 514394 202412
rect 514450 202356 514518 202412
rect 514574 202356 514642 202412
rect 514698 202356 514766 202412
rect 514822 202356 514890 202412
rect 514946 202356 515014 202412
rect 515070 202356 515138 202412
rect 515194 202356 534022 202412
rect 534078 202356 534146 202412
rect 534202 202356 534270 202412
rect 534326 202356 534394 202412
rect 534450 202356 534518 202412
rect 534574 202356 534642 202412
rect 534698 202356 534766 202412
rect 534822 202356 534890 202412
rect 534946 202356 535014 202412
rect 535070 202356 535138 202412
rect 535194 202356 597980 202412
rect -1916 202350 597980 202356
rect -1916 202294 -860 202350
rect -804 202294 -736 202350
rect -680 202294 -612 202350
rect -556 202294 -488 202350
rect -432 202294 3250 202350
rect 3306 202294 3374 202350
rect 3430 202294 3498 202350
rect 3554 202294 3622 202350
rect 3678 202294 21250 202350
rect 21306 202294 21374 202350
rect 21430 202294 21498 202350
rect 21554 202294 21622 202350
rect 21678 202294 39250 202350
rect 39306 202294 39374 202350
rect 39430 202294 39498 202350
rect 39554 202294 39622 202350
rect 39678 202294 57250 202350
rect 57306 202294 57374 202350
rect 57430 202294 57498 202350
rect 57554 202294 57622 202350
rect 57678 202294 64518 202350
rect 64574 202294 64642 202350
rect 64698 202294 95238 202350
rect 95294 202294 95362 202350
rect 95418 202294 125958 202350
rect 126014 202294 126082 202350
rect 126138 202294 156678 202350
rect 156734 202294 156802 202350
rect 156858 202294 187398 202350
rect 187454 202294 187522 202350
rect 187578 202294 218118 202350
rect 218174 202294 218242 202350
rect 218298 202294 255250 202350
rect 255306 202294 255374 202350
rect 255430 202294 255498 202350
rect 255554 202294 255622 202350
rect 255678 202294 273250 202350
rect 273306 202294 273374 202350
rect 273430 202294 273498 202350
rect 273554 202294 273622 202350
rect 273678 202294 291250 202350
rect 291306 202294 291374 202350
rect 291430 202294 291498 202350
rect 291554 202294 291622 202350
rect 291678 202294 309250 202350
rect 309306 202294 309374 202350
rect 309430 202294 309498 202350
rect 309554 202294 309622 202350
rect 309678 202294 327250 202350
rect 327306 202294 327374 202350
rect 327430 202294 327498 202350
rect 327554 202294 327622 202350
rect 327678 202294 345250 202350
rect 345306 202294 345374 202350
rect 345430 202294 345498 202350
rect 345554 202294 345622 202350
rect 345678 202294 561250 202350
rect 561306 202294 561374 202350
rect 561430 202294 561498 202350
rect 561554 202294 561622 202350
rect 561678 202294 579250 202350
rect 579306 202294 579374 202350
rect 579430 202294 579498 202350
rect 579554 202294 579622 202350
rect 579678 202294 596496 202350
rect 596552 202294 596620 202350
rect 596676 202294 596744 202350
rect 596800 202294 596868 202350
rect 596924 202294 597980 202350
rect -1916 202288 597980 202294
rect -1916 202232 354022 202288
rect 354078 202232 354146 202288
rect 354202 202232 354270 202288
rect 354326 202232 354394 202288
rect 354450 202232 354518 202288
rect 354574 202232 354642 202288
rect 354698 202232 354766 202288
rect 354822 202232 354890 202288
rect 354946 202232 355014 202288
rect 355070 202232 355138 202288
rect 355194 202232 374022 202288
rect 374078 202232 374146 202288
rect 374202 202232 374270 202288
rect 374326 202232 374394 202288
rect 374450 202232 374518 202288
rect 374574 202232 374642 202288
rect 374698 202232 374766 202288
rect 374822 202232 374890 202288
rect 374946 202232 375014 202288
rect 375070 202232 375138 202288
rect 375194 202232 394022 202288
rect 394078 202232 394146 202288
rect 394202 202232 394270 202288
rect 394326 202232 394394 202288
rect 394450 202232 394518 202288
rect 394574 202232 394642 202288
rect 394698 202232 394766 202288
rect 394822 202232 394890 202288
rect 394946 202232 395014 202288
rect 395070 202232 395138 202288
rect 395194 202232 414022 202288
rect 414078 202232 414146 202288
rect 414202 202232 414270 202288
rect 414326 202232 414394 202288
rect 414450 202232 414518 202288
rect 414574 202232 414642 202288
rect 414698 202232 414766 202288
rect 414822 202232 414890 202288
rect 414946 202232 415014 202288
rect 415070 202232 415138 202288
rect 415194 202232 434022 202288
rect 434078 202232 434146 202288
rect 434202 202232 434270 202288
rect 434326 202232 434394 202288
rect 434450 202232 434518 202288
rect 434574 202232 434642 202288
rect 434698 202232 434766 202288
rect 434822 202232 434890 202288
rect 434946 202232 435014 202288
rect 435070 202232 435138 202288
rect 435194 202232 454022 202288
rect 454078 202232 454146 202288
rect 454202 202232 454270 202288
rect 454326 202232 454394 202288
rect 454450 202232 454518 202288
rect 454574 202232 454642 202288
rect 454698 202232 454766 202288
rect 454822 202232 454890 202288
rect 454946 202232 455014 202288
rect 455070 202232 455138 202288
rect 455194 202232 474022 202288
rect 474078 202232 474146 202288
rect 474202 202232 474270 202288
rect 474326 202232 474394 202288
rect 474450 202232 474518 202288
rect 474574 202232 474642 202288
rect 474698 202232 474766 202288
rect 474822 202232 474890 202288
rect 474946 202232 475014 202288
rect 475070 202232 475138 202288
rect 475194 202232 494022 202288
rect 494078 202232 494146 202288
rect 494202 202232 494270 202288
rect 494326 202232 494394 202288
rect 494450 202232 494518 202288
rect 494574 202232 494642 202288
rect 494698 202232 494766 202288
rect 494822 202232 494890 202288
rect 494946 202232 495014 202288
rect 495070 202232 495138 202288
rect 495194 202232 514022 202288
rect 514078 202232 514146 202288
rect 514202 202232 514270 202288
rect 514326 202232 514394 202288
rect 514450 202232 514518 202288
rect 514574 202232 514642 202288
rect 514698 202232 514766 202288
rect 514822 202232 514890 202288
rect 514946 202232 515014 202288
rect 515070 202232 515138 202288
rect 515194 202232 534022 202288
rect 534078 202232 534146 202288
rect 534202 202232 534270 202288
rect 534326 202232 534394 202288
rect 534450 202232 534518 202288
rect 534574 202232 534642 202288
rect 534698 202232 534766 202288
rect 534822 202232 534890 202288
rect 534946 202232 535014 202288
rect 535070 202232 535138 202288
rect 535194 202232 597980 202288
rect -1916 202226 597980 202232
rect -1916 202170 -860 202226
rect -804 202170 -736 202226
rect -680 202170 -612 202226
rect -556 202170 -488 202226
rect -432 202170 3250 202226
rect 3306 202170 3374 202226
rect 3430 202170 3498 202226
rect 3554 202170 3622 202226
rect 3678 202170 21250 202226
rect 21306 202170 21374 202226
rect 21430 202170 21498 202226
rect 21554 202170 21622 202226
rect 21678 202170 39250 202226
rect 39306 202170 39374 202226
rect 39430 202170 39498 202226
rect 39554 202170 39622 202226
rect 39678 202170 57250 202226
rect 57306 202170 57374 202226
rect 57430 202170 57498 202226
rect 57554 202170 57622 202226
rect 57678 202170 64518 202226
rect 64574 202170 64642 202226
rect 64698 202170 95238 202226
rect 95294 202170 95362 202226
rect 95418 202170 125958 202226
rect 126014 202170 126082 202226
rect 126138 202170 156678 202226
rect 156734 202170 156802 202226
rect 156858 202170 187398 202226
rect 187454 202170 187522 202226
rect 187578 202170 218118 202226
rect 218174 202170 218242 202226
rect 218298 202170 255250 202226
rect 255306 202170 255374 202226
rect 255430 202170 255498 202226
rect 255554 202170 255622 202226
rect 255678 202170 273250 202226
rect 273306 202170 273374 202226
rect 273430 202170 273498 202226
rect 273554 202170 273622 202226
rect 273678 202170 291250 202226
rect 291306 202170 291374 202226
rect 291430 202170 291498 202226
rect 291554 202170 291622 202226
rect 291678 202170 309250 202226
rect 309306 202170 309374 202226
rect 309430 202170 309498 202226
rect 309554 202170 309622 202226
rect 309678 202170 327250 202226
rect 327306 202170 327374 202226
rect 327430 202170 327498 202226
rect 327554 202170 327622 202226
rect 327678 202170 345250 202226
rect 345306 202170 345374 202226
rect 345430 202170 345498 202226
rect 345554 202170 345622 202226
rect 345678 202170 561250 202226
rect 561306 202170 561374 202226
rect 561430 202170 561498 202226
rect 561554 202170 561622 202226
rect 561678 202170 579250 202226
rect 579306 202170 579374 202226
rect 579430 202170 579498 202226
rect 579554 202170 579622 202226
rect 579678 202170 596496 202226
rect 596552 202170 596620 202226
rect 596676 202170 596744 202226
rect 596800 202170 596868 202226
rect 596924 202170 597980 202226
rect -1916 202164 597980 202170
rect -1916 202108 354022 202164
rect 354078 202108 354146 202164
rect 354202 202108 354270 202164
rect 354326 202108 354394 202164
rect 354450 202108 354518 202164
rect 354574 202108 354642 202164
rect 354698 202108 354766 202164
rect 354822 202108 354890 202164
rect 354946 202108 355014 202164
rect 355070 202108 355138 202164
rect 355194 202108 374022 202164
rect 374078 202108 374146 202164
rect 374202 202108 374270 202164
rect 374326 202108 374394 202164
rect 374450 202108 374518 202164
rect 374574 202108 374642 202164
rect 374698 202108 374766 202164
rect 374822 202108 374890 202164
rect 374946 202108 375014 202164
rect 375070 202108 375138 202164
rect 375194 202108 394022 202164
rect 394078 202108 394146 202164
rect 394202 202108 394270 202164
rect 394326 202108 394394 202164
rect 394450 202108 394518 202164
rect 394574 202108 394642 202164
rect 394698 202108 394766 202164
rect 394822 202108 394890 202164
rect 394946 202108 395014 202164
rect 395070 202108 395138 202164
rect 395194 202108 414022 202164
rect 414078 202108 414146 202164
rect 414202 202108 414270 202164
rect 414326 202108 414394 202164
rect 414450 202108 414518 202164
rect 414574 202108 414642 202164
rect 414698 202108 414766 202164
rect 414822 202108 414890 202164
rect 414946 202108 415014 202164
rect 415070 202108 415138 202164
rect 415194 202108 434022 202164
rect 434078 202108 434146 202164
rect 434202 202108 434270 202164
rect 434326 202108 434394 202164
rect 434450 202108 434518 202164
rect 434574 202108 434642 202164
rect 434698 202108 434766 202164
rect 434822 202108 434890 202164
rect 434946 202108 435014 202164
rect 435070 202108 435138 202164
rect 435194 202108 454022 202164
rect 454078 202108 454146 202164
rect 454202 202108 454270 202164
rect 454326 202108 454394 202164
rect 454450 202108 454518 202164
rect 454574 202108 454642 202164
rect 454698 202108 454766 202164
rect 454822 202108 454890 202164
rect 454946 202108 455014 202164
rect 455070 202108 455138 202164
rect 455194 202108 474022 202164
rect 474078 202108 474146 202164
rect 474202 202108 474270 202164
rect 474326 202108 474394 202164
rect 474450 202108 474518 202164
rect 474574 202108 474642 202164
rect 474698 202108 474766 202164
rect 474822 202108 474890 202164
rect 474946 202108 475014 202164
rect 475070 202108 475138 202164
rect 475194 202108 494022 202164
rect 494078 202108 494146 202164
rect 494202 202108 494270 202164
rect 494326 202108 494394 202164
rect 494450 202108 494518 202164
rect 494574 202108 494642 202164
rect 494698 202108 494766 202164
rect 494822 202108 494890 202164
rect 494946 202108 495014 202164
rect 495070 202108 495138 202164
rect 495194 202108 514022 202164
rect 514078 202108 514146 202164
rect 514202 202108 514270 202164
rect 514326 202108 514394 202164
rect 514450 202108 514518 202164
rect 514574 202108 514642 202164
rect 514698 202108 514766 202164
rect 514822 202108 514890 202164
rect 514946 202108 515014 202164
rect 515070 202108 515138 202164
rect 515194 202108 534022 202164
rect 534078 202108 534146 202164
rect 534202 202108 534270 202164
rect 534326 202108 534394 202164
rect 534450 202108 534518 202164
rect 534574 202108 534642 202164
rect 534698 202108 534766 202164
rect 534822 202108 534890 202164
rect 534946 202108 535014 202164
rect 535070 202108 535138 202164
rect 535194 202108 597980 202164
rect -1916 202102 597980 202108
rect -1916 202046 -860 202102
rect -804 202046 -736 202102
rect -680 202046 -612 202102
rect -556 202046 -488 202102
rect -432 202046 3250 202102
rect 3306 202046 3374 202102
rect 3430 202046 3498 202102
rect 3554 202046 3622 202102
rect 3678 202046 21250 202102
rect 21306 202046 21374 202102
rect 21430 202046 21498 202102
rect 21554 202046 21622 202102
rect 21678 202046 39250 202102
rect 39306 202046 39374 202102
rect 39430 202046 39498 202102
rect 39554 202046 39622 202102
rect 39678 202046 57250 202102
rect 57306 202046 57374 202102
rect 57430 202046 57498 202102
rect 57554 202046 57622 202102
rect 57678 202046 64518 202102
rect 64574 202046 64642 202102
rect 64698 202046 95238 202102
rect 95294 202046 95362 202102
rect 95418 202046 125958 202102
rect 126014 202046 126082 202102
rect 126138 202046 156678 202102
rect 156734 202046 156802 202102
rect 156858 202046 187398 202102
rect 187454 202046 187522 202102
rect 187578 202046 218118 202102
rect 218174 202046 218242 202102
rect 218298 202046 255250 202102
rect 255306 202046 255374 202102
rect 255430 202046 255498 202102
rect 255554 202046 255622 202102
rect 255678 202046 273250 202102
rect 273306 202046 273374 202102
rect 273430 202046 273498 202102
rect 273554 202046 273622 202102
rect 273678 202046 291250 202102
rect 291306 202046 291374 202102
rect 291430 202046 291498 202102
rect 291554 202046 291622 202102
rect 291678 202046 309250 202102
rect 309306 202046 309374 202102
rect 309430 202046 309498 202102
rect 309554 202046 309622 202102
rect 309678 202046 327250 202102
rect 327306 202046 327374 202102
rect 327430 202046 327498 202102
rect 327554 202046 327622 202102
rect 327678 202046 345250 202102
rect 345306 202046 345374 202102
rect 345430 202046 345498 202102
rect 345554 202046 345622 202102
rect 345678 202046 561250 202102
rect 561306 202046 561374 202102
rect 561430 202046 561498 202102
rect 561554 202046 561622 202102
rect 561678 202046 579250 202102
rect 579306 202046 579374 202102
rect 579430 202046 579498 202102
rect 579554 202046 579622 202102
rect 579678 202046 596496 202102
rect 596552 202046 596620 202102
rect 596676 202046 596744 202102
rect 596800 202046 596868 202102
rect 596924 202046 597980 202102
rect -1916 202040 597980 202046
rect -1916 201984 354022 202040
rect 354078 201984 354146 202040
rect 354202 201984 354270 202040
rect 354326 201984 354394 202040
rect 354450 201984 354518 202040
rect 354574 201984 354642 202040
rect 354698 201984 354766 202040
rect 354822 201984 354890 202040
rect 354946 201984 355014 202040
rect 355070 201984 355138 202040
rect 355194 201984 374022 202040
rect 374078 201984 374146 202040
rect 374202 201984 374270 202040
rect 374326 201984 374394 202040
rect 374450 201984 374518 202040
rect 374574 201984 374642 202040
rect 374698 201984 374766 202040
rect 374822 201984 374890 202040
rect 374946 201984 375014 202040
rect 375070 201984 375138 202040
rect 375194 201984 394022 202040
rect 394078 201984 394146 202040
rect 394202 201984 394270 202040
rect 394326 201984 394394 202040
rect 394450 201984 394518 202040
rect 394574 201984 394642 202040
rect 394698 201984 394766 202040
rect 394822 201984 394890 202040
rect 394946 201984 395014 202040
rect 395070 201984 395138 202040
rect 395194 201984 414022 202040
rect 414078 201984 414146 202040
rect 414202 201984 414270 202040
rect 414326 201984 414394 202040
rect 414450 201984 414518 202040
rect 414574 201984 414642 202040
rect 414698 201984 414766 202040
rect 414822 201984 414890 202040
rect 414946 201984 415014 202040
rect 415070 201984 415138 202040
rect 415194 201984 434022 202040
rect 434078 201984 434146 202040
rect 434202 201984 434270 202040
rect 434326 201984 434394 202040
rect 434450 201984 434518 202040
rect 434574 201984 434642 202040
rect 434698 201984 434766 202040
rect 434822 201984 434890 202040
rect 434946 201984 435014 202040
rect 435070 201984 435138 202040
rect 435194 201984 454022 202040
rect 454078 201984 454146 202040
rect 454202 201984 454270 202040
rect 454326 201984 454394 202040
rect 454450 201984 454518 202040
rect 454574 201984 454642 202040
rect 454698 201984 454766 202040
rect 454822 201984 454890 202040
rect 454946 201984 455014 202040
rect 455070 201984 455138 202040
rect 455194 201984 474022 202040
rect 474078 201984 474146 202040
rect 474202 201984 474270 202040
rect 474326 201984 474394 202040
rect 474450 201984 474518 202040
rect 474574 201984 474642 202040
rect 474698 201984 474766 202040
rect 474822 201984 474890 202040
rect 474946 201984 475014 202040
rect 475070 201984 475138 202040
rect 475194 201984 494022 202040
rect 494078 201984 494146 202040
rect 494202 201984 494270 202040
rect 494326 201984 494394 202040
rect 494450 201984 494518 202040
rect 494574 201984 494642 202040
rect 494698 201984 494766 202040
rect 494822 201984 494890 202040
rect 494946 201984 495014 202040
rect 495070 201984 495138 202040
rect 495194 201984 514022 202040
rect 514078 201984 514146 202040
rect 514202 201984 514270 202040
rect 514326 201984 514394 202040
rect 514450 201984 514518 202040
rect 514574 201984 514642 202040
rect 514698 201984 514766 202040
rect 514822 201984 514890 202040
rect 514946 201984 515014 202040
rect 515070 201984 515138 202040
rect 515194 201984 534022 202040
rect 534078 201984 534146 202040
rect 534202 201984 534270 202040
rect 534326 201984 534394 202040
rect 534450 201984 534518 202040
rect 534574 201984 534642 202040
rect 534698 201984 534766 202040
rect 534822 201984 534890 202040
rect 534946 201984 535014 202040
rect 535070 201984 535138 202040
rect 535194 201984 597980 202040
rect -1916 201978 597980 201984
rect -1916 201922 -860 201978
rect -804 201922 -736 201978
rect -680 201922 -612 201978
rect -556 201922 -488 201978
rect -432 201922 3250 201978
rect 3306 201922 3374 201978
rect 3430 201922 3498 201978
rect 3554 201922 3622 201978
rect 3678 201922 21250 201978
rect 21306 201922 21374 201978
rect 21430 201922 21498 201978
rect 21554 201922 21622 201978
rect 21678 201922 39250 201978
rect 39306 201922 39374 201978
rect 39430 201922 39498 201978
rect 39554 201922 39622 201978
rect 39678 201922 57250 201978
rect 57306 201922 57374 201978
rect 57430 201922 57498 201978
rect 57554 201922 57622 201978
rect 57678 201922 64518 201978
rect 64574 201922 64642 201978
rect 64698 201922 95238 201978
rect 95294 201922 95362 201978
rect 95418 201922 125958 201978
rect 126014 201922 126082 201978
rect 126138 201922 156678 201978
rect 156734 201922 156802 201978
rect 156858 201922 187398 201978
rect 187454 201922 187522 201978
rect 187578 201922 218118 201978
rect 218174 201922 218242 201978
rect 218298 201922 255250 201978
rect 255306 201922 255374 201978
rect 255430 201922 255498 201978
rect 255554 201922 255622 201978
rect 255678 201922 273250 201978
rect 273306 201922 273374 201978
rect 273430 201922 273498 201978
rect 273554 201922 273622 201978
rect 273678 201922 291250 201978
rect 291306 201922 291374 201978
rect 291430 201922 291498 201978
rect 291554 201922 291622 201978
rect 291678 201922 309250 201978
rect 309306 201922 309374 201978
rect 309430 201922 309498 201978
rect 309554 201922 309622 201978
rect 309678 201922 327250 201978
rect 327306 201922 327374 201978
rect 327430 201922 327498 201978
rect 327554 201922 327622 201978
rect 327678 201922 345250 201978
rect 345306 201922 345374 201978
rect 345430 201922 345498 201978
rect 345554 201922 345622 201978
rect 345678 201922 561250 201978
rect 561306 201922 561374 201978
rect 561430 201922 561498 201978
rect 561554 201922 561622 201978
rect 561678 201922 579250 201978
rect 579306 201922 579374 201978
rect 579430 201922 579498 201978
rect 579554 201922 579622 201978
rect 579678 201922 596496 201978
rect 596552 201922 596620 201978
rect 596676 201922 596744 201978
rect 596800 201922 596868 201978
rect 596924 201922 597980 201978
rect -1916 201916 597980 201922
rect -1916 201860 354022 201916
rect 354078 201860 354146 201916
rect 354202 201860 354270 201916
rect 354326 201860 354394 201916
rect 354450 201860 354518 201916
rect 354574 201860 354642 201916
rect 354698 201860 354766 201916
rect 354822 201860 354890 201916
rect 354946 201860 355014 201916
rect 355070 201860 355138 201916
rect 355194 201860 374022 201916
rect 374078 201860 374146 201916
rect 374202 201860 374270 201916
rect 374326 201860 374394 201916
rect 374450 201860 374518 201916
rect 374574 201860 374642 201916
rect 374698 201860 374766 201916
rect 374822 201860 374890 201916
rect 374946 201860 375014 201916
rect 375070 201860 375138 201916
rect 375194 201860 394022 201916
rect 394078 201860 394146 201916
rect 394202 201860 394270 201916
rect 394326 201860 394394 201916
rect 394450 201860 394518 201916
rect 394574 201860 394642 201916
rect 394698 201860 394766 201916
rect 394822 201860 394890 201916
rect 394946 201860 395014 201916
rect 395070 201860 395138 201916
rect 395194 201860 414022 201916
rect 414078 201860 414146 201916
rect 414202 201860 414270 201916
rect 414326 201860 414394 201916
rect 414450 201860 414518 201916
rect 414574 201860 414642 201916
rect 414698 201860 414766 201916
rect 414822 201860 414890 201916
rect 414946 201860 415014 201916
rect 415070 201860 415138 201916
rect 415194 201860 434022 201916
rect 434078 201860 434146 201916
rect 434202 201860 434270 201916
rect 434326 201860 434394 201916
rect 434450 201860 434518 201916
rect 434574 201860 434642 201916
rect 434698 201860 434766 201916
rect 434822 201860 434890 201916
rect 434946 201860 435014 201916
rect 435070 201860 435138 201916
rect 435194 201860 454022 201916
rect 454078 201860 454146 201916
rect 454202 201860 454270 201916
rect 454326 201860 454394 201916
rect 454450 201860 454518 201916
rect 454574 201860 454642 201916
rect 454698 201860 454766 201916
rect 454822 201860 454890 201916
rect 454946 201860 455014 201916
rect 455070 201860 455138 201916
rect 455194 201860 474022 201916
rect 474078 201860 474146 201916
rect 474202 201860 474270 201916
rect 474326 201860 474394 201916
rect 474450 201860 474518 201916
rect 474574 201860 474642 201916
rect 474698 201860 474766 201916
rect 474822 201860 474890 201916
rect 474946 201860 475014 201916
rect 475070 201860 475138 201916
rect 475194 201860 494022 201916
rect 494078 201860 494146 201916
rect 494202 201860 494270 201916
rect 494326 201860 494394 201916
rect 494450 201860 494518 201916
rect 494574 201860 494642 201916
rect 494698 201860 494766 201916
rect 494822 201860 494890 201916
rect 494946 201860 495014 201916
rect 495070 201860 495138 201916
rect 495194 201860 514022 201916
rect 514078 201860 514146 201916
rect 514202 201860 514270 201916
rect 514326 201860 514394 201916
rect 514450 201860 514518 201916
rect 514574 201860 514642 201916
rect 514698 201860 514766 201916
rect 514822 201860 514890 201916
rect 514946 201860 515014 201916
rect 515070 201860 515138 201916
rect 515194 201860 534022 201916
rect 534078 201860 534146 201916
rect 534202 201860 534270 201916
rect 534326 201860 534394 201916
rect 534450 201860 534518 201916
rect 534574 201860 534642 201916
rect 534698 201860 534766 201916
rect 534822 201860 534890 201916
rect 534946 201860 535014 201916
rect 535070 201860 535138 201916
rect 535194 201860 597980 201916
rect -1916 201826 597980 201860
rect -1916 190350 66564 190446
rect -1916 190294 -1820 190350
rect -1764 190294 -1696 190350
rect -1640 190294 -1572 190350
rect -1516 190294 -1448 190350
rect -1392 190294 6970 190350
rect 7026 190294 7094 190350
rect 7150 190294 7218 190350
rect 7274 190294 7342 190350
rect 7398 190294 24970 190350
rect 25026 190294 25094 190350
rect 25150 190294 25218 190350
rect 25274 190294 25342 190350
rect 25398 190294 42970 190350
rect 43026 190294 43094 190350
rect 43150 190294 43218 190350
rect 43274 190294 43342 190350
rect 43398 190294 66564 190350
rect -1916 190226 66564 190294
rect -1916 190170 -1820 190226
rect -1764 190170 -1696 190226
rect -1640 190170 -1572 190226
rect -1516 190170 -1448 190226
rect -1392 190170 6970 190226
rect 7026 190170 7094 190226
rect 7150 190170 7218 190226
rect 7274 190170 7342 190226
rect 7398 190170 24970 190226
rect 25026 190170 25094 190226
rect 25150 190170 25218 190226
rect 25274 190170 25342 190226
rect 25398 190170 42970 190226
rect 43026 190170 43094 190226
rect 43150 190170 43218 190226
rect 43274 190170 43342 190226
rect 43398 190170 66564 190226
rect -1916 190102 66564 190170
rect -1916 190046 -1820 190102
rect -1764 190046 -1696 190102
rect -1640 190046 -1572 190102
rect -1516 190046 -1448 190102
rect -1392 190046 6970 190102
rect 7026 190046 7094 190102
rect 7150 190046 7218 190102
rect 7274 190046 7342 190102
rect 7398 190046 24970 190102
rect 25026 190046 25094 190102
rect 25150 190046 25218 190102
rect 25274 190046 25342 190102
rect 25398 190046 42970 190102
rect 43026 190046 43094 190102
rect 43150 190046 43218 190102
rect 43274 190046 43342 190102
rect 43398 190046 66564 190102
rect -1916 189978 66564 190046
rect -1916 189922 -1820 189978
rect -1764 189922 -1696 189978
rect -1640 189922 -1572 189978
rect -1516 189922 -1448 189978
rect -1392 189922 6970 189978
rect 7026 189922 7094 189978
rect 7150 189922 7218 189978
rect 7274 189922 7342 189978
rect 7398 189922 24970 189978
rect 25026 189922 25094 189978
rect 25150 189922 25218 189978
rect 25274 189922 25342 189978
rect 25398 189922 42970 189978
rect 43026 189922 43094 189978
rect 43150 189922 43218 189978
rect 43274 189922 43342 189978
rect 43398 189922 66564 189978
rect -1916 189826 66564 189922
rect 239468 190350 350740 190446
rect 239468 190294 240970 190350
rect 241026 190294 241094 190350
rect 241150 190294 241218 190350
rect 241274 190294 241342 190350
rect 241398 190294 258970 190350
rect 259026 190294 259094 190350
rect 259150 190294 259218 190350
rect 259274 190294 259342 190350
rect 259398 190294 276970 190350
rect 277026 190294 277094 190350
rect 277150 190294 277218 190350
rect 277274 190294 277342 190350
rect 277398 190294 294970 190350
rect 295026 190294 295094 190350
rect 295150 190294 295218 190350
rect 295274 190294 295342 190350
rect 295398 190294 312970 190350
rect 313026 190294 313094 190350
rect 313150 190294 313218 190350
rect 313274 190294 313342 190350
rect 313398 190294 330970 190350
rect 331026 190294 331094 190350
rect 331150 190294 331218 190350
rect 331274 190294 331342 190350
rect 331398 190294 348970 190350
rect 349026 190294 349094 190350
rect 349150 190294 349218 190350
rect 349274 190294 349342 190350
rect 349398 190294 350740 190350
rect 239468 190226 350740 190294
rect 239468 190170 240970 190226
rect 241026 190170 241094 190226
rect 241150 190170 241218 190226
rect 241274 190170 241342 190226
rect 241398 190170 258970 190226
rect 259026 190170 259094 190226
rect 259150 190170 259218 190226
rect 259274 190170 259342 190226
rect 259398 190170 276970 190226
rect 277026 190170 277094 190226
rect 277150 190170 277218 190226
rect 277274 190170 277342 190226
rect 277398 190170 294970 190226
rect 295026 190170 295094 190226
rect 295150 190170 295218 190226
rect 295274 190170 295342 190226
rect 295398 190170 312970 190226
rect 313026 190170 313094 190226
rect 313150 190170 313218 190226
rect 313274 190170 313342 190226
rect 313398 190170 330970 190226
rect 331026 190170 331094 190226
rect 331150 190170 331218 190226
rect 331274 190170 331342 190226
rect 331398 190170 348970 190226
rect 349026 190170 349094 190226
rect 349150 190170 349218 190226
rect 349274 190170 349342 190226
rect 349398 190170 350740 190226
rect 239468 190102 350740 190170
rect 239468 190046 240970 190102
rect 241026 190046 241094 190102
rect 241150 190046 241218 190102
rect 241274 190046 241342 190102
rect 241398 190046 258970 190102
rect 259026 190046 259094 190102
rect 259150 190046 259218 190102
rect 259274 190046 259342 190102
rect 259398 190046 276970 190102
rect 277026 190046 277094 190102
rect 277150 190046 277218 190102
rect 277274 190046 277342 190102
rect 277398 190046 294970 190102
rect 295026 190046 295094 190102
rect 295150 190046 295218 190102
rect 295274 190046 295342 190102
rect 295398 190046 312970 190102
rect 313026 190046 313094 190102
rect 313150 190046 313218 190102
rect 313274 190046 313342 190102
rect 313398 190046 330970 190102
rect 331026 190046 331094 190102
rect 331150 190046 331218 190102
rect 331274 190046 331342 190102
rect 331398 190046 348970 190102
rect 349026 190046 349094 190102
rect 349150 190046 349218 190102
rect 349274 190046 349342 190102
rect 349398 190046 350740 190102
rect 239468 189978 350740 190046
rect 239468 189922 240970 189978
rect 241026 189922 241094 189978
rect 241150 189922 241218 189978
rect 241274 189922 241342 189978
rect 241398 189922 258970 189978
rect 259026 189922 259094 189978
rect 259150 189922 259218 189978
rect 259274 189922 259342 189978
rect 259398 189922 276970 189978
rect 277026 189922 277094 189978
rect 277150 189922 277218 189978
rect 277274 189922 277342 189978
rect 277398 189922 294970 189978
rect 295026 189922 295094 189978
rect 295150 189922 295218 189978
rect 295274 189922 295342 189978
rect 295398 189922 312970 189978
rect 313026 189922 313094 189978
rect 313150 189922 313218 189978
rect 313274 189922 313342 189978
rect 313398 189922 330970 189978
rect 331026 189922 331094 189978
rect 331150 189922 331218 189978
rect 331274 189922 331342 189978
rect 331398 189922 348970 189978
rect 349026 189922 349094 189978
rect 349150 189922 349218 189978
rect 349274 189922 349342 189978
rect 349398 189922 350740 189978
rect 239468 189826 350740 189922
rect 545484 190350 597980 190446
rect 545484 190294 564970 190350
rect 565026 190294 565094 190350
rect 565150 190294 565218 190350
rect 565274 190294 565342 190350
rect 565398 190294 582970 190350
rect 583026 190294 583094 190350
rect 583150 190294 583218 190350
rect 583274 190294 583342 190350
rect 583398 190294 597456 190350
rect 597512 190294 597580 190350
rect 597636 190294 597704 190350
rect 597760 190294 597828 190350
rect 597884 190294 597980 190350
rect 545484 190226 597980 190294
rect 545484 190170 564970 190226
rect 565026 190170 565094 190226
rect 565150 190170 565218 190226
rect 565274 190170 565342 190226
rect 565398 190170 582970 190226
rect 583026 190170 583094 190226
rect 583150 190170 583218 190226
rect 583274 190170 583342 190226
rect 583398 190170 597456 190226
rect 597512 190170 597580 190226
rect 597636 190170 597704 190226
rect 597760 190170 597828 190226
rect 597884 190170 597980 190226
rect 545484 190102 597980 190170
rect 545484 190046 564970 190102
rect 565026 190046 565094 190102
rect 565150 190046 565218 190102
rect 565274 190046 565342 190102
rect 565398 190046 582970 190102
rect 583026 190046 583094 190102
rect 583150 190046 583218 190102
rect 583274 190046 583342 190102
rect 583398 190046 597456 190102
rect 597512 190046 597580 190102
rect 597636 190046 597704 190102
rect 597760 190046 597828 190102
rect 597884 190046 597980 190102
rect 545484 189978 597980 190046
rect 545484 189922 564970 189978
rect 565026 189922 565094 189978
rect 565150 189922 565218 189978
rect 565274 189922 565342 189978
rect 565398 189922 582970 189978
rect 583026 189922 583094 189978
rect 583150 189922 583218 189978
rect 583274 189922 583342 189978
rect 583398 189922 597456 189978
rect 597512 189922 597580 189978
rect 597636 189922 597704 189978
rect 597760 189922 597828 189978
rect 597884 189922 597980 189978
rect 545484 189826 597980 189922
rect -1916 184350 66564 184446
rect -1916 184294 -860 184350
rect -804 184294 -736 184350
rect -680 184294 -612 184350
rect -556 184294 -488 184350
rect -432 184294 3250 184350
rect 3306 184294 3374 184350
rect 3430 184294 3498 184350
rect 3554 184294 3622 184350
rect 3678 184294 21250 184350
rect 21306 184294 21374 184350
rect 21430 184294 21498 184350
rect 21554 184294 21622 184350
rect 21678 184294 39250 184350
rect 39306 184294 39374 184350
rect 39430 184294 39498 184350
rect 39554 184294 39622 184350
rect 39678 184294 57250 184350
rect 57306 184294 57374 184350
rect 57430 184294 57498 184350
rect 57554 184294 57622 184350
rect 57678 184294 64518 184350
rect 64574 184294 64642 184350
rect 64698 184294 66564 184350
rect -1916 184226 66564 184294
rect -1916 184170 -860 184226
rect -804 184170 -736 184226
rect -680 184170 -612 184226
rect -556 184170 -488 184226
rect -432 184170 3250 184226
rect 3306 184170 3374 184226
rect 3430 184170 3498 184226
rect 3554 184170 3622 184226
rect 3678 184170 21250 184226
rect 21306 184170 21374 184226
rect 21430 184170 21498 184226
rect 21554 184170 21622 184226
rect 21678 184170 39250 184226
rect 39306 184170 39374 184226
rect 39430 184170 39498 184226
rect 39554 184170 39622 184226
rect 39678 184170 57250 184226
rect 57306 184170 57374 184226
rect 57430 184170 57498 184226
rect 57554 184170 57622 184226
rect 57678 184170 64518 184226
rect 64574 184170 64642 184226
rect 64698 184170 66564 184226
rect -1916 184102 66564 184170
rect -1916 184046 -860 184102
rect -804 184046 -736 184102
rect -680 184046 -612 184102
rect -556 184046 -488 184102
rect -432 184046 3250 184102
rect 3306 184046 3374 184102
rect 3430 184046 3498 184102
rect 3554 184046 3622 184102
rect 3678 184046 21250 184102
rect 21306 184046 21374 184102
rect 21430 184046 21498 184102
rect 21554 184046 21622 184102
rect 21678 184046 39250 184102
rect 39306 184046 39374 184102
rect 39430 184046 39498 184102
rect 39554 184046 39622 184102
rect 39678 184046 57250 184102
rect 57306 184046 57374 184102
rect 57430 184046 57498 184102
rect 57554 184046 57622 184102
rect 57678 184046 64518 184102
rect 64574 184046 64642 184102
rect 64698 184046 66564 184102
rect -1916 183978 66564 184046
rect -1916 183922 -860 183978
rect -804 183922 -736 183978
rect -680 183922 -612 183978
rect -556 183922 -488 183978
rect -432 183922 3250 183978
rect 3306 183922 3374 183978
rect 3430 183922 3498 183978
rect 3554 183922 3622 183978
rect 3678 183922 21250 183978
rect 21306 183922 21374 183978
rect 21430 183922 21498 183978
rect 21554 183922 21622 183978
rect 21678 183922 39250 183978
rect 39306 183922 39374 183978
rect 39430 183922 39498 183978
rect 39554 183922 39622 183978
rect 39678 183922 57250 183978
rect 57306 183922 57374 183978
rect 57430 183922 57498 183978
rect 57554 183922 57622 183978
rect 57678 183922 64518 183978
rect 64574 183922 64642 183978
rect 64698 183922 66564 183978
rect -1916 183826 66564 183922
rect 239468 184350 350740 184446
rect 239468 184294 255250 184350
rect 255306 184294 255374 184350
rect 255430 184294 255498 184350
rect 255554 184294 255622 184350
rect 255678 184294 273250 184350
rect 273306 184294 273374 184350
rect 273430 184294 273498 184350
rect 273554 184294 273622 184350
rect 273678 184294 291250 184350
rect 291306 184294 291374 184350
rect 291430 184294 291498 184350
rect 291554 184294 291622 184350
rect 291678 184294 309250 184350
rect 309306 184294 309374 184350
rect 309430 184294 309498 184350
rect 309554 184294 309622 184350
rect 309678 184294 327250 184350
rect 327306 184294 327374 184350
rect 327430 184294 327498 184350
rect 327554 184294 327622 184350
rect 327678 184294 345250 184350
rect 345306 184294 345374 184350
rect 345430 184294 345498 184350
rect 345554 184294 345622 184350
rect 345678 184294 350740 184350
rect 239468 184226 350740 184294
rect 239468 184170 255250 184226
rect 255306 184170 255374 184226
rect 255430 184170 255498 184226
rect 255554 184170 255622 184226
rect 255678 184170 273250 184226
rect 273306 184170 273374 184226
rect 273430 184170 273498 184226
rect 273554 184170 273622 184226
rect 273678 184170 291250 184226
rect 291306 184170 291374 184226
rect 291430 184170 291498 184226
rect 291554 184170 291622 184226
rect 291678 184170 309250 184226
rect 309306 184170 309374 184226
rect 309430 184170 309498 184226
rect 309554 184170 309622 184226
rect 309678 184170 327250 184226
rect 327306 184170 327374 184226
rect 327430 184170 327498 184226
rect 327554 184170 327622 184226
rect 327678 184170 345250 184226
rect 345306 184170 345374 184226
rect 345430 184170 345498 184226
rect 345554 184170 345622 184226
rect 345678 184170 350740 184226
rect 239468 184102 350740 184170
rect 239468 184046 255250 184102
rect 255306 184046 255374 184102
rect 255430 184046 255498 184102
rect 255554 184046 255622 184102
rect 255678 184046 273250 184102
rect 273306 184046 273374 184102
rect 273430 184046 273498 184102
rect 273554 184046 273622 184102
rect 273678 184046 291250 184102
rect 291306 184046 291374 184102
rect 291430 184046 291498 184102
rect 291554 184046 291622 184102
rect 291678 184046 309250 184102
rect 309306 184046 309374 184102
rect 309430 184046 309498 184102
rect 309554 184046 309622 184102
rect 309678 184046 327250 184102
rect 327306 184046 327374 184102
rect 327430 184046 327498 184102
rect 327554 184046 327622 184102
rect 327678 184046 345250 184102
rect 345306 184046 345374 184102
rect 345430 184046 345498 184102
rect 345554 184046 345622 184102
rect 345678 184046 350740 184102
rect 239468 183978 350740 184046
rect 239468 183922 255250 183978
rect 255306 183922 255374 183978
rect 255430 183922 255498 183978
rect 255554 183922 255622 183978
rect 255678 183922 273250 183978
rect 273306 183922 273374 183978
rect 273430 183922 273498 183978
rect 273554 183922 273622 183978
rect 273678 183922 291250 183978
rect 291306 183922 291374 183978
rect 291430 183922 291498 183978
rect 291554 183922 291622 183978
rect 291678 183922 309250 183978
rect 309306 183922 309374 183978
rect 309430 183922 309498 183978
rect 309554 183922 309622 183978
rect 309678 183922 327250 183978
rect 327306 183922 327374 183978
rect 327430 183922 327498 183978
rect 327554 183922 327622 183978
rect 327678 183922 345250 183978
rect 345306 183922 345374 183978
rect 345430 183922 345498 183978
rect 345554 183922 345622 183978
rect 345678 183922 350740 183978
rect 239468 183826 350740 183922
rect 545484 184350 597980 184446
rect 545484 184294 561250 184350
rect 561306 184294 561374 184350
rect 561430 184294 561498 184350
rect 561554 184294 561622 184350
rect 561678 184294 579250 184350
rect 579306 184294 579374 184350
rect 579430 184294 579498 184350
rect 579554 184294 579622 184350
rect 579678 184294 596496 184350
rect 596552 184294 596620 184350
rect 596676 184294 596744 184350
rect 596800 184294 596868 184350
rect 596924 184294 597980 184350
rect 545484 184226 597980 184294
rect 545484 184170 561250 184226
rect 561306 184170 561374 184226
rect 561430 184170 561498 184226
rect 561554 184170 561622 184226
rect 561678 184170 579250 184226
rect 579306 184170 579374 184226
rect 579430 184170 579498 184226
rect 579554 184170 579622 184226
rect 579678 184170 596496 184226
rect 596552 184170 596620 184226
rect 596676 184170 596744 184226
rect 596800 184170 596868 184226
rect 596924 184170 597980 184226
rect 545484 184102 597980 184170
rect 545484 184046 561250 184102
rect 561306 184046 561374 184102
rect 561430 184046 561498 184102
rect 561554 184046 561622 184102
rect 561678 184046 579250 184102
rect 579306 184046 579374 184102
rect 579430 184046 579498 184102
rect 579554 184046 579622 184102
rect 579678 184046 596496 184102
rect 596552 184046 596620 184102
rect 596676 184046 596744 184102
rect 596800 184046 596868 184102
rect 596924 184046 597980 184102
rect 545484 183978 597980 184046
rect 545484 183922 561250 183978
rect 561306 183922 561374 183978
rect 561430 183922 561498 183978
rect 561554 183922 561622 183978
rect 561678 183922 579250 183978
rect 579306 183922 579374 183978
rect 579430 183922 579498 183978
rect 579554 183922 579622 183978
rect 579678 183922 596496 183978
rect 596552 183922 596620 183978
rect 596676 183922 596744 183978
rect 596800 183922 596868 183978
rect 596924 183922 597980 183978
rect 545484 183826 597980 183922
rect -1916 172350 66564 172446
rect -1916 172294 -1820 172350
rect -1764 172294 -1696 172350
rect -1640 172294 -1572 172350
rect -1516 172294 -1448 172350
rect -1392 172294 6970 172350
rect 7026 172294 7094 172350
rect 7150 172294 7218 172350
rect 7274 172294 7342 172350
rect 7398 172294 24970 172350
rect 25026 172294 25094 172350
rect 25150 172294 25218 172350
rect 25274 172294 25342 172350
rect 25398 172294 42970 172350
rect 43026 172294 43094 172350
rect 43150 172294 43218 172350
rect 43274 172294 43342 172350
rect 43398 172294 66564 172350
rect -1916 172226 66564 172294
rect -1916 172170 -1820 172226
rect -1764 172170 -1696 172226
rect -1640 172170 -1572 172226
rect -1516 172170 -1448 172226
rect -1392 172170 6970 172226
rect 7026 172170 7094 172226
rect 7150 172170 7218 172226
rect 7274 172170 7342 172226
rect 7398 172170 24970 172226
rect 25026 172170 25094 172226
rect 25150 172170 25218 172226
rect 25274 172170 25342 172226
rect 25398 172170 42970 172226
rect 43026 172170 43094 172226
rect 43150 172170 43218 172226
rect 43274 172170 43342 172226
rect 43398 172170 66564 172226
rect -1916 172102 66564 172170
rect -1916 172046 -1820 172102
rect -1764 172046 -1696 172102
rect -1640 172046 -1572 172102
rect -1516 172046 -1448 172102
rect -1392 172046 6970 172102
rect 7026 172046 7094 172102
rect 7150 172046 7218 172102
rect 7274 172046 7342 172102
rect 7398 172046 24970 172102
rect 25026 172046 25094 172102
rect 25150 172046 25218 172102
rect 25274 172046 25342 172102
rect 25398 172046 42970 172102
rect 43026 172046 43094 172102
rect 43150 172046 43218 172102
rect 43274 172046 43342 172102
rect 43398 172046 66564 172102
rect -1916 171978 66564 172046
rect -1916 171922 -1820 171978
rect -1764 171922 -1696 171978
rect -1640 171922 -1572 171978
rect -1516 171922 -1448 171978
rect -1392 171922 6970 171978
rect 7026 171922 7094 171978
rect 7150 171922 7218 171978
rect 7274 171922 7342 171978
rect 7398 171922 24970 171978
rect 25026 171922 25094 171978
rect 25150 171922 25218 171978
rect 25274 171922 25342 171978
rect 25398 171922 42970 171978
rect 43026 171922 43094 171978
rect 43150 171922 43218 171978
rect 43274 171922 43342 171978
rect 43398 171922 66564 171978
rect -1916 171826 66564 171922
rect 239468 172350 350740 172446
rect 239468 172294 240970 172350
rect 241026 172294 241094 172350
rect 241150 172294 241218 172350
rect 241274 172294 241342 172350
rect 241398 172294 258970 172350
rect 259026 172294 259094 172350
rect 259150 172294 259218 172350
rect 259274 172294 259342 172350
rect 259398 172294 276970 172350
rect 277026 172294 277094 172350
rect 277150 172294 277218 172350
rect 277274 172294 277342 172350
rect 277398 172294 294970 172350
rect 295026 172294 295094 172350
rect 295150 172294 295218 172350
rect 295274 172294 295342 172350
rect 295398 172294 312970 172350
rect 313026 172294 313094 172350
rect 313150 172294 313218 172350
rect 313274 172294 313342 172350
rect 313398 172294 330970 172350
rect 331026 172294 331094 172350
rect 331150 172294 331218 172350
rect 331274 172294 331342 172350
rect 331398 172294 348970 172350
rect 349026 172294 349094 172350
rect 349150 172294 349218 172350
rect 349274 172294 349342 172350
rect 349398 172294 350740 172350
rect 239468 172226 350740 172294
rect 239468 172170 240970 172226
rect 241026 172170 241094 172226
rect 241150 172170 241218 172226
rect 241274 172170 241342 172226
rect 241398 172170 258970 172226
rect 259026 172170 259094 172226
rect 259150 172170 259218 172226
rect 259274 172170 259342 172226
rect 259398 172170 276970 172226
rect 277026 172170 277094 172226
rect 277150 172170 277218 172226
rect 277274 172170 277342 172226
rect 277398 172170 294970 172226
rect 295026 172170 295094 172226
rect 295150 172170 295218 172226
rect 295274 172170 295342 172226
rect 295398 172170 312970 172226
rect 313026 172170 313094 172226
rect 313150 172170 313218 172226
rect 313274 172170 313342 172226
rect 313398 172170 330970 172226
rect 331026 172170 331094 172226
rect 331150 172170 331218 172226
rect 331274 172170 331342 172226
rect 331398 172170 348970 172226
rect 349026 172170 349094 172226
rect 349150 172170 349218 172226
rect 349274 172170 349342 172226
rect 349398 172170 350740 172226
rect 239468 172102 350740 172170
rect 239468 172046 240970 172102
rect 241026 172046 241094 172102
rect 241150 172046 241218 172102
rect 241274 172046 241342 172102
rect 241398 172046 258970 172102
rect 259026 172046 259094 172102
rect 259150 172046 259218 172102
rect 259274 172046 259342 172102
rect 259398 172046 276970 172102
rect 277026 172046 277094 172102
rect 277150 172046 277218 172102
rect 277274 172046 277342 172102
rect 277398 172046 294970 172102
rect 295026 172046 295094 172102
rect 295150 172046 295218 172102
rect 295274 172046 295342 172102
rect 295398 172046 312970 172102
rect 313026 172046 313094 172102
rect 313150 172046 313218 172102
rect 313274 172046 313342 172102
rect 313398 172046 330970 172102
rect 331026 172046 331094 172102
rect 331150 172046 331218 172102
rect 331274 172046 331342 172102
rect 331398 172046 348970 172102
rect 349026 172046 349094 172102
rect 349150 172046 349218 172102
rect 349274 172046 349342 172102
rect 349398 172046 350740 172102
rect 239468 171978 350740 172046
rect 239468 171922 240970 171978
rect 241026 171922 241094 171978
rect 241150 171922 241218 171978
rect 241274 171922 241342 171978
rect 241398 171922 258970 171978
rect 259026 171922 259094 171978
rect 259150 171922 259218 171978
rect 259274 171922 259342 171978
rect 259398 171922 276970 171978
rect 277026 171922 277094 171978
rect 277150 171922 277218 171978
rect 277274 171922 277342 171978
rect 277398 171922 294970 171978
rect 295026 171922 295094 171978
rect 295150 171922 295218 171978
rect 295274 171922 295342 171978
rect 295398 171922 312970 171978
rect 313026 171922 313094 171978
rect 313150 171922 313218 171978
rect 313274 171922 313342 171978
rect 313398 171922 330970 171978
rect 331026 171922 331094 171978
rect 331150 171922 331218 171978
rect 331274 171922 331342 171978
rect 331398 171922 348970 171978
rect 349026 171922 349094 171978
rect 349150 171922 349218 171978
rect 349274 171922 349342 171978
rect 349398 171922 350740 171978
rect 239468 171826 350740 171922
rect 545484 172350 597980 172446
rect 545484 172294 564970 172350
rect 565026 172294 565094 172350
rect 565150 172294 565218 172350
rect 565274 172294 565342 172350
rect 565398 172294 582970 172350
rect 583026 172294 583094 172350
rect 583150 172294 583218 172350
rect 583274 172294 583342 172350
rect 583398 172294 597456 172350
rect 597512 172294 597580 172350
rect 597636 172294 597704 172350
rect 597760 172294 597828 172350
rect 597884 172294 597980 172350
rect 545484 172226 597980 172294
rect 545484 172170 564970 172226
rect 565026 172170 565094 172226
rect 565150 172170 565218 172226
rect 565274 172170 565342 172226
rect 565398 172170 582970 172226
rect 583026 172170 583094 172226
rect 583150 172170 583218 172226
rect 583274 172170 583342 172226
rect 583398 172170 597456 172226
rect 597512 172170 597580 172226
rect 597636 172170 597704 172226
rect 597760 172170 597828 172226
rect 597884 172170 597980 172226
rect 545484 172102 597980 172170
rect 545484 172046 564970 172102
rect 565026 172046 565094 172102
rect 565150 172046 565218 172102
rect 565274 172046 565342 172102
rect 565398 172046 582970 172102
rect 583026 172046 583094 172102
rect 583150 172046 583218 172102
rect 583274 172046 583342 172102
rect 583398 172046 597456 172102
rect 597512 172046 597580 172102
rect 597636 172046 597704 172102
rect 597760 172046 597828 172102
rect 597884 172046 597980 172102
rect 545484 171978 597980 172046
rect 545484 171922 564970 171978
rect 565026 171922 565094 171978
rect 565150 171922 565218 171978
rect 565274 171922 565342 171978
rect 565398 171922 582970 171978
rect 583026 171922 583094 171978
rect 583150 171922 583218 171978
rect 583274 171922 583342 171978
rect 583398 171922 597456 171978
rect 597512 171922 597580 171978
rect 597636 171922 597704 171978
rect 597760 171922 597828 171978
rect 597884 171922 597980 171978
rect 545484 171826 597980 171922
rect -1916 166350 66564 166446
rect -1916 166294 -860 166350
rect -804 166294 -736 166350
rect -680 166294 -612 166350
rect -556 166294 -488 166350
rect -432 166294 3250 166350
rect 3306 166294 3374 166350
rect 3430 166294 3498 166350
rect 3554 166294 3622 166350
rect 3678 166294 21250 166350
rect 21306 166294 21374 166350
rect 21430 166294 21498 166350
rect 21554 166294 21622 166350
rect 21678 166294 39250 166350
rect 39306 166294 39374 166350
rect 39430 166294 39498 166350
rect 39554 166294 39622 166350
rect 39678 166294 57250 166350
rect 57306 166294 57374 166350
rect 57430 166294 57498 166350
rect 57554 166294 57622 166350
rect 57678 166294 64518 166350
rect 64574 166294 64642 166350
rect 64698 166294 66564 166350
rect -1916 166226 66564 166294
rect -1916 166170 -860 166226
rect -804 166170 -736 166226
rect -680 166170 -612 166226
rect -556 166170 -488 166226
rect -432 166170 3250 166226
rect 3306 166170 3374 166226
rect 3430 166170 3498 166226
rect 3554 166170 3622 166226
rect 3678 166170 21250 166226
rect 21306 166170 21374 166226
rect 21430 166170 21498 166226
rect 21554 166170 21622 166226
rect 21678 166170 39250 166226
rect 39306 166170 39374 166226
rect 39430 166170 39498 166226
rect 39554 166170 39622 166226
rect 39678 166170 57250 166226
rect 57306 166170 57374 166226
rect 57430 166170 57498 166226
rect 57554 166170 57622 166226
rect 57678 166170 64518 166226
rect 64574 166170 64642 166226
rect 64698 166170 66564 166226
rect -1916 166102 66564 166170
rect -1916 166046 -860 166102
rect -804 166046 -736 166102
rect -680 166046 -612 166102
rect -556 166046 -488 166102
rect -432 166046 3250 166102
rect 3306 166046 3374 166102
rect 3430 166046 3498 166102
rect 3554 166046 3622 166102
rect 3678 166046 21250 166102
rect 21306 166046 21374 166102
rect 21430 166046 21498 166102
rect 21554 166046 21622 166102
rect 21678 166046 39250 166102
rect 39306 166046 39374 166102
rect 39430 166046 39498 166102
rect 39554 166046 39622 166102
rect 39678 166046 57250 166102
rect 57306 166046 57374 166102
rect 57430 166046 57498 166102
rect 57554 166046 57622 166102
rect 57678 166046 64518 166102
rect 64574 166046 64642 166102
rect 64698 166046 66564 166102
rect -1916 165978 66564 166046
rect -1916 165922 -860 165978
rect -804 165922 -736 165978
rect -680 165922 -612 165978
rect -556 165922 -488 165978
rect -432 165922 3250 165978
rect 3306 165922 3374 165978
rect 3430 165922 3498 165978
rect 3554 165922 3622 165978
rect 3678 165922 21250 165978
rect 21306 165922 21374 165978
rect 21430 165922 21498 165978
rect 21554 165922 21622 165978
rect 21678 165922 39250 165978
rect 39306 165922 39374 165978
rect 39430 165922 39498 165978
rect 39554 165922 39622 165978
rect 39678 165922 57250 165978
rect 57306 165922 57374 165978
rect 57430 165922 57498 165978
rect 57554 165922 57622 165978
rect 57678 165922 64518 165978
rect 64574 165922 64642 165978
rect 64698 165922 66564 165978
rect -1916 165826 66564 165922
rect 239468 166412 350740 166446
rect 239468 166356 284022 166412
rect 284078 166356 284146 166412
rect 284202 166356 284270 166412
rect 284326 166356 284394 166412
rect 284450 166356 284518 166412
rect 284574 166356 284642 166412
rect 284698 166356 284766 166412
rect 284822 166356 284890 166412
rect 284946 166356 285014 166412
rect 285070 166356 285138 166412
rect 285194 166356 304022 166412
rect 304078 166356 304146 166412
rect 304202 166356 304270 166412
rect 304326 166356 304394 166412
rect 304450 166356 304518 166412
rect 304574 166356 304642 166412
rect 304698 166356 304766 166412
rect 304822 166356 304890 166412
rect 304946 166356 305014 166412
rect 305070 166356 305138 166412
rect 305194 166356 350740 166412
rect 239468 166350 350740 166356
rect 239468 166294 255250 166350
rect 255306 166294 255374 166350
rect 255430 166294 255498 166350
rect 255554 166294 255622 166350
rect 255678 166294 273250 166350
rect 273306 166294 273374 166350
rect 273430 166294 273498 166350
rect 273554 166294 273622 166350
rect 273678 166294 291250 166350
rect 291306 166294 291374 166350
rect 291430 166294 291498 166350
rect 291554 166294 291622 166350
rect 291678 166294 309250 166350
rect 309306 166294 309374 166350
rect 309430 166294 309498 166350
rect 309554 166294 309622 166350
rect 309678 166294 327250 166350
rect 327306 166294 327374 166350
rect 327430 166294 327498 166350
rect 327554 166294 327622 166350
rect 327678 166294 345250 166350
rect 345306 166294 345374 166350
rect 345430 166294 345498 166350
rect 345554 166294 345622 166350
rect 345678 166294 350740 166350
rect 239468 166288 350740 166294
rect 239468 166232 284022 166288
rect 284078 166232 284146 166288
rect 284202 166232 284270 166288
rect 284326 166232 284394 166288
rect 284450 166232 284518 166288
rect 284574 166232 284642 166288
rect 284698 166232 284766 166288
rect 284822 166232 284890 166288
rect 284946 166232 285014 166288
rect 285070 166232 285138 166288
rect 285194 166232 304022 166288
rect 304078 166232 304146 166288
rect 304202 166232 304270 166288
rect 304326 166232 304394 166288
rect 304450 166232 304518 166288
rect 304574 166232 304642 166288
rect 304698 166232 304766 166288
rect 304822 166232 304890 166288
rect 304946 166232 305014 166288
rect 305070 166232 305138 166288
rect 305194 166232 350740 166288
rect 239468 166226 350740 166232
rect 239468 166170 255250 166226
rect 255306 166170 255374 166226
rect 255430 166170 255498 166226
rect 255554 166170 255622 166226
rect 255678 166170 273250 166226
rect 273306 166170 273374 166226
rect 273430 166170 273498 166226
rect 273554 166170 273622 166226
rect 273678 166170 291250 166226
rect 291306 166170 291374 166226
rect 291430 166170 291498 166226
rect 291554 166170 291622 166226
rect 291678 166170 309250 166226
rect 309306 166170 309374 166226
rect 309430 166170 309498 166226
rect 309554 166170 309622 166226
rect 309678 166170 327250 166226
rect 327306 166170 327374 166226
rect 327430 166170 327498 166226
rect 327554 166170 327622 166226
rect 327678 166170 345250 166226
rect 345306 166170 345374 166226
rect 345430 166170 345498 166226
rect 345554 166170 345622 166226
rect 345678 166170 350740 166226
rect 239468 166164 350740 166170
rect 239468 166108 284022 166164
rect 284078 166108 284146 166164
rect 284202 166108 284270 166164
rect 284326 166108 284394 166164
rect 284450 166108 284518 166164
rect 284574 166108 284642 166164
rect 284698 166108 284766 166164
rect 284822 166108 284890 166164
rect 284946 166108 285014 166164
rect 285070 166108 285138 166164
rect 285194 166108 304022 166164
rect 304078 166108 304146 166164
rect 304202 166108 304270 166164
rect 304326 166108 304394 166164
rect 304450 166108 304518 166164
rect 304574 166108 304642 166164
rect 304698 166108 304766 166164
rect 304822 166108 304890 166164
rect 304946 166108 305014 166164
rect 305070 166108 305138 166164
rect 305194 166108 350740 166164
rect 239468 166102 350740 166108
rect 239468 166046 255250 166102
rect 255306 166046 255374 166102
rect 255430 166046 255498 166102
rect 255554 166046 255622 166102
rect 255678 166046 273250 166102
rect 273306 166046 273374 166102
rect 273430 166046 273498 166102
rect 273554 166046 273622 166102
rect 273678 166046 291250 166102
rect 291306 166046 291374 166102
rect 291430 166046 291498 166102
rect 291554 166046 291622 166102
rect 291678 166046 309250 166102
rect 309306 166046 309374 166102
rect 309430 166046 309498 166102
rect 309554 166046 309622 166102
rect 309678 166046 327250 166102
rect 327306 166046 327374 166102
rect 327430 166046 327498 166102
rect 327554 166046 327622 166102
rect 327678 166046 345250 166102
rect 345306 166046 345374 166102
rect 345430 166046 345498 166102
rect 345554 166046 345622 166102
rect 345678 166046 350740 166102
rect 239468 166040 350740 166046
rect 239468 165984 284022 166040
rect 284078 165984 284146 166040
rect 284202 165984 284270 166040
rect 284326 165984 284394 166040
rect 284450 165984 284518 166040
rect 284574 165984 284642 166040
rect 284698 165984 284766 166040
rect 284822 165984 284890 166040
rect 284946 165984 285014 166040
rect 285070 165984 285138 166040
rect 285194 165984 304022 166040
rect 304078 165984 304146 166040
rect 304202 165984 304270 166040
rect 304326 165984 304394 166040
rect 304450 165984 304518 166040
rect 304574 165984 304642 166040
rect 304698 165984 304766 166040
rect 304822 165984 304890 166040
rect 304946 165984 305014 166040
rect 305070 165984 305138 166040
rect 305194 165984 350740 166040
rect 239468 165978 350740 165984
rect 239468 165922 255250 165978
rect 255306 165922 255374 165978
rect 255430 165922 255498 165978
rect 255554 165922 255622 165978
rect 255678 165922 273250 165978
rect 273306 165922 273374 165978
rect 273430 165922 273498 165978
rect 273554 165922 273622 165978
rect 273678 165922 291250 165978
rect 291306 165922 291374 165978
rect 291430 165922 291498 165978
rect 291554 165922 291622 165978
rect 291678 165922 309250 165978
rect 309306 165922 309374 165978
rect 309430 165922 309498 165978
rect 309554 165922 309622 165978
rect 309678 165922 327250 165978
rect 327306 165922 327374 165978
rect 327430 165922 327498 165978
rect 327554 165922 327622 165978
rect 327678 165922 345250 165978
rect 345306 165922 345374 165978
rect 345430 165922 345498 165978
rect 345554 165922 345622 165978
rect 345678 165922 350740 165978
rect 239468 165916 350740 165922
rect 239468 165860 284022 165916
rect 284078 165860 284146 165916
rect 284202 165860 284270 165916
rect 284326 165860 284394 165916
rect 284450 165860 284518 165916
rect 284574 165860 284642 165916
rect 284698 165860 284766 165916
rect 284822 165860 284890 165916
rect 284946 165860 285014 165916
rect 285070 165860 285138 165916
rect 285194 165860 304022 165916
rect 304078 165860 304146 165916
rect 304202 165860 304270 165916
rect 304326 165860 304394 165916
rect 304450 165860 304518 165916
rect 304574 165860 304642 165916
rect 304698 165860 304766 165916
rect 304822 165860 304890 165916
rect 304946 165860 305014 165916
rect 305070 165860 305138 165916
rect 305194 165860 350740 165916
rect 239468 165826 350740 165860
rect 545484 166350 597980 166446
rect 545484 166294 561250 166350
rect 561306 166294 561374 166350
rect 561430 166294 561498 166350
rect 561554 166294 561622 166350
rect 561678 166294 579250 166350
rect 579306 166294 579374 166350
rect 579430 166294 579498 166350
rect 579554 166294 579622 166350
rect 579678 166294 596496 166350
rect 596552 166294 596620 166350
rect 596676 166294 596744 166350
rect 596800 166294 596868 166350
rect 596924 166294 597980 166350
rect 545484 166226 597980 166294
rect 545484 166170 561250 166226
rect 561306 166170 561374 166226
rect 561430 166170 561498 166226
rect 561554 166170 561622 166226
rect 561678 166170 579250 166226
rect 579306 166170 579374 166226
rect 579430 166170 579498 166226
rect 579554 166170 579622 166226
rect 579678 166170 596496 166226
rect 596552 166170 596620 166226
rect 596676 166170 596744 166226
rect 596800 166170 596868 166226
rect 596924 166170 597980 166226
rect 545484 166102 597980 166170
rect 545484 166046 561250 166102
rect 561306 166046 561374 166102
rect 561430 166046 561498 166102
rect 561554 166046 561622 166102
rect 561678 166046 579250 166102
rect 579306 166046 579374 166102
rect 579430 166046 579498 166102
rect 579554 166046 579622 166102
rect 579678 166046 596496 166102
rect 596552 166046 596620 166102
rect 596676 166046 596744 166102
rect 596800 166046 596868 166102
rect 596924 166046 597980 166102
rect 545484 165978 597980 166046
rect 545484 165922 561250 165978
rect 561306 165922 561374 165978
rect 561430 165922 561498 165978
rect 561554 165922 561622 165978
rect 561678 165922 579250 165978
rect 579306 165922 579374 165978
rect 579430 165922 579498 165978
rect 579554 165922 579622 165978
rect 579678 165922 596496 165978
rect 596552 165922 596620 165978
rect 596676 165922 596744 165978
rect 596800 165922 596868 165978
rect 596924 165922 597980 165978
rect 545484 165826 597980 165922
rect -1916 154350 66564 154446
rect -1916 154294 -1820 154350
rect -1764 154294 -1696 154350
rect -1640 154294 -1572 154350
rect -1516 154294 -1448 154350
rect -1392 154294 6970 154350
rect 7026 154294 7094 154350
rect 7150 154294 7218 154350
rect 7274 154294 7342 154350
rect 7398 154294 24970 154350
rect 25026 154294 25094 154350
rect 25150 154294 25218 154350
rect 25274 154294 25342 154350
rect 25398 154294 42970 154350
rect 43026 154294 43094 154350
rect 43150 154294 43218 154350
rect 43274 154294 43342 154350
rect 43398 154294 66564 154350
rect -1916 154226 66564 154294
rect -1916 154170 -1820 154226
rect -1764 154170 -1696 154226
rect -1640 154170 -1572 154226
rect -1516 154170 -1448 154226
rect -1392 154170 6970 154226
rect 7026 154170 7094 154226
rect 7150 154170 7218 154226
rect 7274 154170 7342 154226
rect 7398 154170 24970 154226
rect 25026 154170 25094 154226
rect 25150 154170 25218 154226
rect 25274 154170 25342 154226
rect 25398 154170 42970 154226
rect 43026 154170 43094 154226
rect 43150 154170 43218 154226
rect 43274 154170 43342 154226
rect 43398 154170 66564 154226
rect -1916 154102 66564 154170
rect -1916 154046 -1820 154102
rect -1764 154046 -1696 154102
rect -1640 154046 -1572 154102
rect -1516 154046 -1448 154102
rect -1392 154046 6970 154102
rect 7026 154046 7094 154102
rect 7150 154046 7218 154102
rect 7274 154046 7342 154102
rect 7398 154046 24970 154102
rect 25026 154046 25094 154102
rect 25150 154046 25218 154102
rect 25274 154046 25342 154102
rect 25398 154046 42970 154102
rect 43026 154046 43094 154102
rect 43150 154046 43218 154102
rect 43274 154046 43342 154102
rect 43398 154046 66564 154102
rect -1916 153978 66564 154046
rect -1916 153922 -1820 153978
rect -1764 153922 -1696 153978
rect -1640 153922 -1572 153978
rect -1516 153922 -1448 153978
rect -1392 153922 6970 153978
rect 7026 153922 7094 153978
rect 7150 153922 7218 153978
rect 7274 153922 7342 153978
rect 7398 153922 24970 153978
rect 25026 153922 25094 153978
rect 25150 153922 25218 153978
rect 25274 153922 25342 153978
rect 25398 153922 42970 153978
rect 43026 153922 43094 153978
rect 43150 153922 43218 153978
rect 43274 153922 43342 153978
rect 43398 153922 66564 153978
rect -1916 153826 66564 153922
rect 239468 154412 350740 154446
rect 239468 154356 294022 154412
rect 294078 154356 294146 154412
rect 294202 154356 294270 154412
rect 294326 154356 294394 154412
rect 294450 154356 294518 154412
rect 294574 154356 294642 154412
rect 294698 154356 294766 154412
rect 294822 154356 294890 154412
rect 294946 154356 295014 154412
rect 295070 154356 295138 154412
rect 295194 154356 314022 154412
rect 314078 154356 314146 154412
rect 314202 154356 314270 154412
rect 314326 154356 314394 154412
rect 314450 154356 314518 154412
rect 314574 154356 314642 154412
rect 314698 154356 314766 154412
rect 314822 154356 314890 154412
rect 314946 154356 315014 154412
rect 315070 154356 315138 154412
rect 315194 154356 350740 154412
rect 239468 154350 350740 154356
rect 239468 154294 240970 154350
rect 241026 154294 241094 154350
rect 241150 154294 241218 154350
rect 241274 154294 241342 154350
rect 241398 154294 258970 154350
rect 259026 154294 259094 154350
rect 259150 154294 259218 154350
rect 259274 154294 259342 154350
rect 259398 154294 276970 154350
rect 277026 154294 277094 154350
rect 277150 154294 277218 154350
rect 277274 154294 277342 154350
rect 277398 154294 330970 154350
rect 331026 154294 331094 154350
rect 331150 154294 331218 154350
rect 331274 154294 331342 154350
rect 331398 154294 348970 154350
rect 349026 154294 349094 154350
rect 349150 154294 349218 154350
rect 349274 154294 349342 154350
rect 349398 154294 350740 154350
rect 239468 154288 350740 154294
rect 239468 154232 294022 154288
rect 294078 154232 294146 154288
rect 294202 154232 294270 154288
rect 294326 154232 294394 154288
rect 294450 154232 294518 154288
rect 294574 154232 294642 154288
rect 294698 154232 294766 154288
rect 294822 154232 294890 154288
rect 294946 154232 295014 154288
rect 295070 154232 295138 154288
rect 295194 154232 314022 154288
rect 314078 154232 314146 154288
rect 314202 154232 314270 154288
rect 314326 154232 314394 154288
rect 314450 154232 314518 154288
rect 314574 154232 314642 154288
rect 314698 154232 314766 154288
rect 314822 154232 314890 154288
rect 314946 154232 315014 154288
rect 315070 154232 315138 154288
rect 315194 154232 350740 154288
rect 239468 154226 350740 154232
rect 239468 154170 240970 154226
rect 241026 154170 241094 154226
rect 241150 154170 241218 154226
rect 241274 154170 241342 154226
rect 241398 154170 258970 154226
rect 259026 154170 259094 154226
rect 259150 154170 259218 154226
rect 259274 154170 259342 154226
rect 259398 154170 276970 154226
rect 277026 154170 277094 154226
rect 277150 154170 277218 154226
rect 277274 154170 277342 154226
rect 277398 154170 330970 154226
rect 331026 154170 331094 154226
rect 331150 154170 331218 154226
rect 331274 154170 331342 154226
rect 331398 154170 348970 154226
rect 349026 154170 349094 154226
rect 349150 154170 349218 154226
rect 349274 154170 349342 154226
rect 349398 154170 350740 154226
rect 239468 154164 350740 154170
rect 239468 154108 294022 154164
rect 294078 154108 294146 154164
rect 294202 154108 294270 154164
rect 294326 154108 294394 154164
rect 294450 154108 294518 154164
rect 294574 154108 294642 154164
rect 294698 154108 294766 154164
rect 294822 154108 294890 154164
rect 294946 154108 295014 154164
rect 295070 154108 295138 154164
rect 295194 154108 314022 154164
rect 314078 154108 314146 154164
rect 314202 154108 314270 154164
rect 314326 154108 314394 154164
rect 314450 154108 314518 154164
rect 314574 154108 314642 154164
rect 314698 154108 314766 154164
rect 314822 154108 314890 154164
rect 314946 154108 315014 154164
rect 315070 154108 315138 154164
rect 315194 154108 350740 154164
rect 239468 154102 350740 154108
rect 239468 154046 240970 154102
rect 241026 154046 241094 154102
rect 241150 154046 241218 154102
rect 241274 154046 241342 154102
rect 241398 154046 258970 154102
rect 259026 154046 259094 154102
rect 259150 154046 259218 154102
rect 259274 154046 259342 154102
rect 259398 154046 276970 154102
rect 277026 154046 277094 154102
rect 277150 154046 277218 154102
rect 277274 154046 277342 154102
rect 277398 154046 330970 154102
rect 331026 154046 331094 154102
rect 331150 154046 331218 154102
rect 331274 154046 331342 154102
rect 331398 154046 348970 154102
rect 349026 154046 349094 154102
rect 349150 154046 349218 154102
rect 349274 154046 349342 154102
rect 349398 154046 350740 154102
rect 239468 154040 350740 154046
rect 239468 153984 294022 154040
rect 294078 153984 294146 154040
rect 294202 153984 294270 154040
rect 294326 153984 294394 154040
rect 294450 153984 294518 154040
rect 294574 153984 294642 154040
rect 294698 153984 294766 154040
rect 294822 153984 294890 154040
rect 294946 153984 295014 154040
rect 295070 153984 295138 154040
rect 295194 153984 314022 154040
rect 314078 153984 314146 154040
rect 314202 153984 314270 154040
rect 314326 153984 314394 154040
rect 314450 153984 314518 154040
rect 314574 153984 314642 154040
rect 314698 153984 314766 154040
rect 314822 153984 314890 154040
rect 314946 153984 315014 154040
rect 315070 153984 315138 154040
rect 315194 153984 350740 154040
rect 239468 153978 350740 153984
rect 239468 153922 240970 153978
rect 241026 153922 241094 153978
rect 241150 153922 241218 153978
rect 241274 153922 241342 153978
rect 241398 153922 258970 153978
rect 259026 153922 259094 153978
rect 259150 153922 259218 153978
rect 259274 153922 259342 153978
rect 259398 153922 276970 153978
rect 277026 153922 277094 153978
rect 277150 153922 277218 153978
rect 277274 153922 277342 153978
rect 277398 153922 330970 153978
rect 331026 153922 331094 153978
rect 331150 153922 331218 153978
rect 331274 153922 331342 153978
rect 331398 153922 348970 153978
rect 349026 153922 349094 153978
rect 349150 153922 349218 153978
rect 349274 153922 349342 153978
rect 349398 153922 350740 153978
rect 239468 153916 350740 153922
rect 239468 153860 294022 153916
rect 294078 153860 294146 153916
rect 294202 153860 294270 153916
rect 294326 153860 294394 153916
rect 294450 153860 294518 153916
rect 294574 153860 294642 153916
rect 294698 153860 294766 153916
rect 294822 153860 294890 153916
rect 294946 153860 295014 153916
rect 295070 153860 295138 153916
rect 295194 153860 314022 153916
rect 314078 153860 314146 153916
rect 314202 153860 314270 153916
rect 314326 153860 314394 153916
rect 314450 153860 314518 153916
rect 314574 153860 314642 153916
rect 314698 153860 314766 153916
rect 314822 153860 314890 153916
rect 314946 153860 315014 153916
rect 315070 153860 315138 153916
rect 315194 153860 350740 153916
rect 239468 153826 350740 153860
rect 545484 154350 597980 154446
rect 545484 154294 564970 154350
rect 565026 154294 565094 154350
rect 565150 154294 565218 154350
rect 565274 154294 565342 154350
rect 565398 154294 582970 154350
rect 583026 154294 583094 154350
rect 583150 154294 583218 154350
rect 583274 154294 583342 154350
rect 583398 154294 597456 154350
rect 597512 154294 597580 154350
rect 597636 154294 597704 154350
rect 597760 154294 597828 154350
rect 597884 154294 597980 154350
rect 545484 154226 597980 154294
rect 545484 154170 564970 154226
rect 565026 154170 565094 154226
rect 565150 154170 565218 154226
rect 565274 154170 565342 154226
rect 565398 154170 582970 154226
rect 583026 154170 583094 154226
rect 583150 154170 583218 154226
rect 583274 154170 583342 154226
rect 583398 154170 597456 154226
rect 597512 154170 597580 154226
rect 597636 154170 597704 154226
rect 597760 154170 597828 154226
rect 597884 154170 597980 154226
rect 545484 154102 597980 154170
rect 545484 154046 564970 154102
rect 565026 154046 565094 154102
rect 565150 154046 565218 154102
rect 565274 154046 565342 154102
rect 565398 154046 582970 154102
rect 583026 154046 583094 154102
rect 583150 154046 583218 154102
rect 583274 154046 583342 154102
rect 583398 154046 597456 154102
rect 597512 154046 597580 154102
rect 597636 154046 597704 154102
rect 597760 154046 597828 154102
rect 597884 154046 597980 154102
rect 545484 153978 597980 154046
rect 545484 153922 564970 153978
rect 565026 153922 565094 153978
rect 565150 153922 565218 153978
rect 565274 153922 565342 153978
rect 565398 153922 582970 153978
rect 583026 153922 583094 153978
rect 583150 153922 583218 153978
rect 583274 153922 583342 153978
rect 583398 153922 597456 153978
rect 597512 153922 597580 153978
rect 597636 153922 597704 153978
rect 597760 153922 597828 153978
rect 597884 153922 597980 153978
rect 545484 153826 597980 153922
rect -1916 148350 66564 148446
rect -1916 148294 -860 148350
rect -804 148294 -736 148350
rect -680 148294 -612 148350
rect -556 148294 -488 148350
rect -432 148294 3250 148350
rect 3306 148294 3374 148350
rect 3430 148294 3498 148350
rect 3554 148294 3622 148350
rect 3678 148294 21250 148350
rect 21306 148294 21374 148350
rect 21430 148294 21498 148350
rect 21554 148294 21622 148350
rect 21678 148294 39250 148350
rect 39306 148294 39374 148350
rect 39430 148294 39498 148350
rect 39554 148294 39622 148350
rect 39678 148294 57250 148350
rect 57306 148294 57374 148350
rect 57430 148294 57498 148350
rect 57554 148294 57622 148350
rect 57678 148294 64518 148350
rect 64574 148294 64642 148350
rect 64698 148294 66564 148350
rect -1916 148226 66564 148294
rect -1916 148170 -860 148226
rect -804 148170 -736 148226
rect -680 148170 -612 148226
rect -556 148170 -488 148226
rect -432 148170 3250 148226
rect 3306 148170 3374 148226
rect 3430 148170 3498 148226
rect 3554 148170 3622 148226
rect 3678 148170 21250 148226
rect 21306 148170 21374 148226
rect 21430 148170 21498 148226
rect 21554 148170 21622 148226
rect 21678 148170 39250 148226
rect 39306 148170 39374 148226
rect 39430 148170 39498 148226
rect 39554 148170 39622 148226
rect 39678 148170 57250 148226
rect 57306 148170 57374 148226
rect 57430 148170 57498 148226
rect 57554 148170 57622 148226
rect 57678 148170 64518 148226
rect 64574 148170 64642 148226
rect 64698 148170 66564 148226
rect -1916 148102 66564 148170
rect -1916 148046 -860 148102
rect -804 148046 -736 148102
rect -680 148046 -612 148102
rect -556 148046 -488 148102
rect -432 148046 3250 148102
rect 3306 148046 3374 148102
rect 3430 148046 3498 148102
rect 3554 148046 3622 148102
rect 3678 148046 21250 148102
rect 21306 148046 21374 148102
rect 21430 148046 21498 148102
rect 21554 148046 21622 148102
rect 21678 148046 39250 148102
rect 39306 148046 39374 148102
rect 39430 148046 39498 148102
rect 39554 148046 39622 148102
rect 39678 148046 57250 148102
rect 57306 148046 57374 148102
rect 57430 148046 57498 148102
rect 57554 148046 57622 148102
rect 57678 148046 64518 148102
rect 64574 148046 64642 148102
rect 64698 148046 66564 148102
rect -1916 147978 66564 148046
rect -1916 147922 -860 147978
rect -804 147922 -736 147978
rect -680 147922 -612 147978
rect -556 147922 -488 147978
rect -432 147922 3250 147978
rect 3306 147922 3374 147978
rect 3430 147922 3498 147978
rect 3554 147922 3622 147978
rect 3678 147922 21250 147978
rect 21306 147922 21374 147978
rect 21430 147922 21498 147978
rect 21554 147922 21622 147978
rect 21678 147922 39250 147978
rect 39306 147922 39374 147978
rect 39430 147922 39498 147978
rect 39554 147922 39622 147978
rect 39678 147922 57250 147978
rect 57306 147922 57374 147978
rect 57430 147922 57498 147978
rect 57554 147922 57622 147978
rect 57678 147922 64518 147978
rect 64574 147922 64642 147978
rect 64698 147922 66564 147978
rect -1916 147826 66564 147922
rect 239468 148412 350740 148446
rect 239468 148356 284022 148412
rect 284078 148356 284146 148412
rect 284202 148356 284270 148412
rect 284326 148356 284394 148412
rect 284450 148356 284518 148412
rect 284574 148356 284642 148412
rect 284698 148356 284766 148412
rect 284822 148356 284890 148412
rect 284946 148356 285014 148412
rect 285070 148356 285138 148412
rect 285194 148356 304022 148412
rect 304078 148356 304146 148412
rect 304202 148356 304270 148412
rect 304326 148356 304394 148412
rect 304450 148356 304518 148412
rect 304574 148356 304642 148412
rect 304698 148356 304766 148412
rect 304822 148356 304890 148412
rect 304946 148356 305014 148412
rect 305070 148356 305138 148412
rect 305194 148356 350740 148412
rect 239468 148350 350740 148356
rect 239468 148294 255250 148350
rect 255306 148294 255374 148350
rect 255430 148294 255498 148350
rect 255554 148294 255622 148350
rect 255678 148294 273250 148350
rect 273306 148294 273374 148350
rect 273430 148294 273498 148350
rect 273554 148294 273622 148350
rect 273678 148294 327250 148350
rect 327306 148294 327374 148350
rect 327430 148294 327498 148350
rect 327554 148294 327622 148350
rect 327678 148294 345250 148350
rect 345306 148294 345374 148350
rect 345430 148294 345498 148350
rect 345554 148294 345622 148350
rect 345678 148294 350740 148350
rect 239468 148288 350740 148294
rect 239468 148232 284022 148288
rect 284078 148232 284146 148288
rect 284202 148232 284270 148288
rect 284326 148232 284394 148288
rect 284450 148232 284518 148288
rect 284574 148232 284642 148288
rect 284698 148232 284766 148288
rect 284822 148232 284890 148288
rect 284946 148232 285014 148288
rect 285070 148232 285138 148288
rect 285194 148232 304022 148288
rect 304078 148232 304146 148288
rect 304202 148232 304270 148288
rect 304326 148232 304394 148288
rect 304450 148232 304518 148288
rect 304574 148232 304642 148288
rect 304698 148232 304766 148288
rect 304822 148232 304890 148288
rect 304946 148232 305014 148288
rect 305070 148232 305138 148288
rect 305194 148232 350740 148288
rect 239468 148226 350740 148232
rect 239468 148170 255250 148226
rect 255306 148170 255374 148226
rect 255430 148170 255498 148226
rect 255554 148170 255622 148226
rect 255678 148170 273250 148226
rect 273306 148170 273374 148226
rect 273430 148170 273498 148226
rect 273554 148170 273622 148226
rect 273678 148170 327250 148226
rect 327306 148170 327374 148226
rect 327430 148170 327498 148226
rect 327554 148170 327622 148226
rect 327678 148170 345250 148226
rect 345306 148170 345374 148226
rect 345430 148170 345498 148226
rect 345554 148170 345622 148226
rect 345678 148170 350740 148226
rect 239468 148164 350740 148170
rect 239468 148108 284022 148164
rect 284078 148108 284146 148164
rect 284202 148108 284270 148164
rect 284326 148108 284394 148164
rect 284450 148108 284518 148164
rect 284574 148108 284642 148164
rect 284698 148108 284766 148164
rect 284822 148108 284890 148164
rect 284946 148108 285014 148164
rect 285070 148108 285138 148164
rect 285194 148108 304022 148164
rect 304078 148108 304146 148164
rect 304202 148108 304270 148164
rect 304326 148108 304394 148164
rect 304450 148108 304518 148164
rect 304574 148108 304642 148164
rect 304698 148108 304766 148164
rect 304822 148108 304890 148164
rect 304946 148108 305014 148164
rect 305070 148108 305138 148164
rect 305194 148108 350740 148164
rect 239468 148102 350740 148108
rect 239468 148046 255250 148102
rect 255306 148046 255374 148102
rect 255430 148046 255498 148102
rect 255554 148046 255622 148102
rect 255678 148046 273250 148102
rect 273306 148046 273374 148102
rect 273430 148046 273498 148102
rect 273554 148046 273622 148102
rect 273678 148046 327250 148102
rect 327306 148046 327374 148102
rect 327430 148046 327498 148102
rect 327554 148046 327622 148102
rect 327678 148046 345250 148102
rect 345306 148046 345374 148102
rect 345430 148046 345498 148102
rect 345554 148046 345622 148102
rect 345678 148046 350740 148102
rect 239468 148040 350740 148046
rect 239468 147984 284022 148040
rect 284078 147984 284146 148040
rect 284202 147984 284270 148040
rect 284326 147984 284394 148040
rect 284450 147984 284518 148040
rect 284574 147984 284642 148040
rect 284698 147984 284766 148040
rect 284822 147984 284890 148040
rect 284946 147984 285014 148040
rect 285070 147984 285138 148040
rect 285194 147984 304022 148040
rect 304078 147984 304146 148040
rect 304202 147984 304270 148040
rect 304326 147984 304394 148040
rect 304450 147984 304518 148040
rect 304574 147984 304642 148040
rect 304698 147984 304766 148040
rect 304822 147984 304890 148040
rect 304946 147984 305014 148040
rect 305070 147984 305138 148040
rect 305194 147984 350740 148040
rect 239468 147978 350740 147984
rect 239468 147922 255250 147978
rect 255306 147922 255374 147978
rect 255430 147922 255498 147978
rect 255554 147922 255622 147978
rect 255678 147922 273250 147978
rect 273306 147922 273374 147978
rect 273430 147922 273498 147978
rect 273554 147922 273622 147978
rect 273678 147922 327250 147978
rect 327306 147922 327374 147978
rect 327430 147922 327498 147978
rect 327554 147922 327622 147978
rect 327678 147922 345250 147978
rect 345306 147922 345374 147978
rect 345430 147922 345498 147978
rect 345554 147922 345622 147978
rect 345678 147922 350740 147978
rect 239468 147916 350740 147922
rect 239468 147860 284022 147916
rect 284078 147860 284146 147916
rect 284202 147860 284270 147916
rect 284326 147860 284394 147916
rect 284450 147860 284518 147916
rect 284574 147860 284642 147916
rect 284698 147860 284766 147916
rect 284822 147860 284890 147916
rect 284946 147860 285014 147916
rect 285070 147860 285138 147916
rect 285194 147860 304022 147916
rect 304078 147860 304146 147916
rect 304202 147860 304270 147916
rect 304326 147860 304394 147916
rect 304450 147860 304518 147916
rect 304574 147860 304642 147916
rect 304698 147860 304766 147916
rect 304822 147860 304890 147916
rect 304946 147860 305014 147916
rect 305070 147860 305138 147916
rect 305194 147860 350740 147916
rect 239468 147826 350740 147860
rect 545484 148350 597980 148446
rect 545484 148294 561250 148350
rect 561306 148294 561374 148350
rect 561430 148294 561498 148350
rect 561554 148294 561622 148350
rect 561678 148294 579250 148350
rect 579306 148294 579374 148350
rect 579430 148294 579498 148350
rect 579554 148294 579622 148350
rect 579678 148294 596496 148350
rect 596552 148294 596620 148350
rect 596676 148294 596744 148350
rect 596800 148294 596868 148350
rect 596924 148294 597980 148350
rect 545484 148226 597980 148294
rect 545484 148170 561250 148226
rect 561306 148170 561374 148226
rect 561430 148170 561498 148226
rect 561554 148170 561622 148226
rect 561678 148170 579250 148226
rect 579306 148170 579374 148226
rect 579430 148170 579498 148226
rect 579554 148170 579622 148226
rect 579678 148170 596496 148226
rect 596552 148170 596620 148226
rect 596676 148170 596744 148226
rect 596800 148170 596868 148226
rect 596924 148170 597980 148226
rect 545484 148102 597980 148170
rect 545484 148046 561250 148102
rect 561306 148046 561374 148102
rect 561430 148046 561498 148102
rect 561554 148046 561622 148102
rect 561678 148046 579250 148102
rect 579306 148046 579374 148102
rect 579430 148046 579498 148102
rect 579554 148046 579622 148102
rect 579678 148046 596496 148102
rect 596552 148046 596620 148102
rect 596676 148046 596744 148102
rect 596800 148046 596868 148102
rect 596924 148046 597980 148102
rect 545484 147978 597980 148046
rect 545484 147922 561250 147978
rect 561306 147922 561374 147978
rect 561430 147922 561498 147978
rect 561554 147922 561622 147978
rect 561678 147922 579250 147978
rect 579306 147922 579374 147978
rect 579430 147922 579498 147978
rect 579554 147922 579622 147978
rect 579678 147922 596496 147978
rect 596552 147922 596620 147978
rect 596676 147922 596744 147978
rect 596800 147922 596868 147978
rect 596924 147922 597980 147978
rect 545484 147826 597980 147922
rect -1916 136350 66564 136446
rect -1916 136294 -1820 136350
rect -1764 136294 -1696 136350
rect -1640 136294 -1572 136350
rect -1516 136294 -1448 136350
rect -1392 136294 6970 136350
rect 7026 136294 7094 136350
rect 7150 136294 7218 136350
rect 7274 136294 7342 136350
rect 7398 136294 24970 136350
rect 25026 136294 25094 136350
rect 25150 136294 25218 136350
rect 25274 136294 25342 136350
rect 25398 136294 42970 136350
rect 43026 136294 43094 136350
rect 43150 136294 43218 136350
rect 43274 136294 43342 136350
rect 43398 136294 66564 136350
rect -1916 136226 66564 136294
rect -1916 136170 -1820 136226
rect -1764 136170 -1696 136226
rect -1640 136170 -1572 136226
rect -1516 136170 -1448 136226
rect -1392 136170 6970 136226
rect 7026 136170 7094 136226
rect 7150 136170 7218 136226
rect 7274 136170 7342 136226
rect 7398 136170 24970 136226
rect 25026 136170 25094 136226
rect 25150 136170 25218 136226
rect 25274 136170 25342 136226
rect 25398 136170 42970 136226
rect 43026 136170 43094 136226
rect 43150 136170 43218 136226
rect 43274 136170 43342 136226
rect 43398 136170 66564 136226
rect -1916 136102 66564 136170
rect -1916 136046 -1820 136102
rect -1764 136046 -1696 136102
rect -1640 136046 -1572 136102
rect -1516 136046 -1448 136102
rect -1392 136046 6970 136102
rect 7026 136046 7094 136102
rect 7150 136046 7218 136102
rect 7274 136046 7342 136102
rect 7398 136046 24970 136102
rect 25026 136046 25094 136102
rect 25150 136046 25218 136102
rect 25274 136046 25342 136102
rect 25398 136046 42970 136102
rect 43026 136046 43094 136102
rect 43150 136046 43218 136102
rect 43274 136046 43342 136102
rect 43398 136046 66564 136102
rect -1916 135978 66564 136046
rect -1916 135922 -1820 135978
rect -1764 135922 -1696 135978
rect -1640 135922 -1572 135978
rect -1516 135922 -1448 135978
rect -1392 135922 6970 135978
rect 7026 135922 7094 135978
rect 7150 135922 7218 135978
rect 7274 135922 7342 135978
rect 7398 135922 24970 135978
rect 25026 135922 25094 135978
rect 25150 135922 25218 135978
rect 25274 135922 25342 135978
rect 25398 135922 42970 135978
rect 43026 135922 43094 135978
rect 43150 135922 43218 135978
rect 43274 135922 43342 135978
rect 43398 135922 66564 135978
rect -1916 135826 66564 135922
rect 239468 136412 350740 136446
rect 239468 136356 294022 136412
rect 294078 136356 294146 136412
rect 294202 136356 294270 136412
rect 294326 136356 294394 136412
rect 294450 136356 294518 136412
rect 294574 136356 294642 136412
rect 294698 136356 294766 136412
rect 294822 136356 294890 136412
rect 294946 136356 295014 136412
rect 295070 136356 295138 136412
rect 295194 136356 314022 136412
rect 314078 136356 314146 136412
rect 314202 136356 314270 136412
rect 314326 136356 314394 136412
rect 314450 136356 314518 136412
rect 314574 136356 314642 136412
rect 314698 136356 314766 136412
rect 314822 136356 314890 136412
rect 314946 136356 315014 136412
rect 315070 136356 315138 136412
rect 315194 136356 350740 136412
rect 239468 136350 350740 136356
rect 239468 136294 240970 136350
rect 241026 136294 241094 136350
rect 241150 136294 241218 136350
rect 241274 136294 241342 136350
rect 241398 136294 258970 136350
rect 259026 136294 259094 136350
rect 259150 136294 259218 136350
rect 259274 136294 259342 136350
rect 259398 136294 276970 136350
rect 277026 136294 277094 136350
rect 277150 136294 277218 136350
rect 277274 136294 277342 136350
rect 277398 136294 330970 136350
rect 331026 136294 331094 136350
rect 331150 136294 331218 136350
rect 331274 136294 331342 136350
rect 331398 136294 348970 136350
rect 349026 136294 349094 136350
rect 349150 136294 349218 136350
rect 349274 136294 349342 136350
rect 349398 136294 350740 136350
rect 239468 136288 350740 136294
rect 239468 136232 294022 136288
rect 294078 136232 294146 136288
rect 294202 136232 294270 136288
rect 294326 136232 294394 136288
rect 294450 136232 294518 136288
rect 294574 136232 294642 136288
rect 294698 136232 294766 136288
rect 294822 136232 294890 136288
rect 294946 136232 295014 136288
rect 295070 136232 295138 136288
rect 295194 136232 314022 136288
rect 314078 136232 314146 136288
rect 314202 136232 314270 136288
rect 314326 136232 314394 136288
rect 314450 136232 314518 136288
rect 314574 136232 314642 136288
rect 314698 136232 314766 136288
rect 314822 136232 314890 136288
rect 314946 136232 315014 136288
rect 315070 136232 315138 136288
rect 315194 136232 350740 136288
rect 239468 136226 350740 136232
rect 239468 136170 240970 136226
rect 241026 136170 241094 136226
rect 241150 136170 241218 136226
rect 241274 136170 241342 136226
rect 241398 136170 258970 136226
rect 259026 136170 259094 136226
rect 259150 136170 259218 136226
rect 259274 136170 259342 136226
rect 259398 136170 276970 136226
rect 277026 136170 277094 136226
rect 277150 136170 277218 136226
rect 277274 136170 277342 136226
rect 277398 136170 330970 136226
rect 331026 136170 331094 136226
rect 331150 136170 331218 136226
rect 331274 136170 331342 136226
rect 331398 136170 348970 136226
rect 349026 136170 349094 136226
rect 349150 136170 349218 136226
rect 349274 136170 349342 136226
rect 349398 136170 350740 136226
rect 239468 136164 350740 136170
rect 239468 136108 294022 136164
rect 294078 136108 294146 136164
rect 294202 136108 294270 136164
rect 294326 136108 294394 136164
rect 294450 136108 294518 136164
rect 294574 136108 294642 136164
rect 294698 136108 294766 136164
rect 294822 136108 294890 136164
rect 294946 136108 295014 136164
rect 295070 136108 295138 136164
rect 295194 136108 314022 136164
rect 314078 136108 314146 136164
rect 314202 136108 314270 136164
rect 314326 136108 314394 136164
rect 314450 136108 314518 136164
rect 314574 136108 314642 136164
rect 314698 136108 314766 136164
rect 314822 136108 314890 136164
rect 314946 136108 315014 136164
rect 315070 136108 315138 136164
rect 315194 136108 350740 136164
rect 239468 136102 350740 136108
rect 239468 136046 240970 136102
rect 241026 136046 241094 136102
rect 241150 136046 241218 136102
rect 241274 136046 241342 136102
rect 241398 136046 258970 136102
rect 259026 136046 259094 136102
rect 259150 136046 259218 136102
rect 259274 136046 259342 136102
rect 259398 136046 276970 136102
rect 277026 136046 277094 136102
rect 277150 136046 277218 136102
rect 277274 136046 277342 136102
rect 277398 136046 330970 136102
rect 331026 136046 331094 136102
rect 331150 136046 331218 136102
rect 331274 136046 331342 136102
rect 331398 136046 348970 136102
rect 349026 136046 349094 136102
rect 349150 136046 349218 136102
rect 349274 136046 349342 136102
rect 349398 136046 350740 136102
rect 239468 136040 350740 136046
rect 239468 135984 294022 136040
rect 294078 135984 294146 136040
rect 294202 135984 294270 136040
rect 294326 135984 294394 136040
rect 294450 135984 294518 136040
rect 294574 135984 294642 136040
rect 294698 135984 294766 136040
rect 294822 135984 294890 136040
rect 294946 135984 295014 136040
rect 295070 135984 295138 136040
rect 295194 135984 314022 136040
rect 314078 135984 314146 136040
rect 314202 135984 314270 136040
rect 314326 135984 314394 136040
rect 314450 135984 314518 136040
rect 314574 135984 314642 136040
rect 314698 135984 314766 136040
rect 314822 135984 314890 136040
rect 314946 135984 315014 136040
rect 315070 135984 315138 136040
rect 315194 135984 350740 136040
rect 239468 135978 350740 135984
rect 239468 135922 240970 135978
rect 241026 135922 241094 135978
rect 241150 135922 241218 135978
rect 241274 135922 241342 135978
rect 241398 135922 258970 135978
rect 259026 135922 259094 135978
rect 259150 135922 259218 135978
rect 259274 135922 259342 135978
rect 259398 135922 276970 135978
rect 277026 135922 277094 135978
rect 277150 135922 277218 135978
rect 277274 135922 277342 135978
rect 277398 135922 330970 135978
rect 331026 135922 331094 135978
rect 331150 135922 331218 135978
rect 331274 135922 331342 135978
rect 331398 135922 348970 135978
rect 349026 135922 349094 135978
rect 349150 135922 349218 135978
rect 349274 135922 349342 135978
rect 349398 135922 350740 135978
rect 239468 135916 350740 135922
rect 239468 135860 294022 135916
rect 294078 135860 294146 135916
rect 294202 135860 294270 135916
rect 294326 135860 294394 135916
rect 294450 135860 294518 135916
rect 294574 135860 294642 135916
rect 294698 135860 294766 135916
rect 294822 135860 294890 135916
rect 294946 135860 295014 135916
rect 295070 135860 295138 135916
rect 295194 135860 314022 135916
rect 314078 135860 314146 135916
rect 314202 135860 314270 135916
rect 314326 135860 314394 135916
rect 314450 135860 314518 135916
rect 314574 135860 314642 135916
rect 314698 135860 314766 135916
rect 314822 135860 314890 135916
rect 314946 135860 315014 135916
rect 315070 135860 315138 135916
rect 315194 135860 350740 135916
rect 239468 135826 350740 135860
rect 545484 136350 597980 136446
rect 545484 136294 564970 136350
rect 565026 136294 565094 136350
rect 565150 136294 565218 136350
rect 565274 136294 565342 136350
rect 565398 136294 582970 136350
rect 583026 136294 583094 136350
rect 583150 136294 583218 136350
rect 583274 136294 583342 136350
rect 583398 136294 597456 136350
rect 597512 136294 597580 136350
rect 597636 136294 597704 136350
rect 597760 136294 597828 136350
rect 597884 136294 597980 136350
rect 545484 136226 597980 136294
rect 545484 136170 564970 136226
rect 565026 136170 565094 136226
rect 565150 136170 565218 136226
rect 565274 136170 565342 136226
rect 565398 136170 582970 136226
rect 583026 136170 583094 136226
rect 583150 136170 583218 136226
rect 583274 136170 583342 136226
rect 583398 136170 597456 136226
rect 597512 136170 597580 136226
rect 597636 136170 597704 136226
rect 597760 136170 597828 136226
rect 597884 136170 597980 136226
rect 545484 136102 597980 136170
rect 545484 136046 564970 136102
rect 565026 136046 565094 136102
rect 565150 136046 565218 136102
rect 565274 136046 565342 136102
rect 565398 136046 582970 136102
rect 583026 136046 583094 136102
rect 583150 136046 583218 136102
rect 583274 136046 583342 136102
rect 583398 136046 597456 136102
rect 597512 136046 597580 136102
rect 597636 136046 597704 136102
rect 597760 136046 597828 136102
rect 597884 136046 597980 136102
rect 545484 135978 597980 136046
rect 545484 135922 564970 135978
rect 565026 135922 565094 135978
rect 565150 135922 565218 135978
rect 565274 135922 565342 135978
rect 565398 135922 582970 135978
rect 583026 135922 583094 135978
rect 583150 135922 583218 135978
rect 583274 135922 583342 135978
rect 583398 135922 597456 135978
rect 597512 135922 597580 135978
rect 597636 135922 597704 135978
rect 597760 135922 597828 135978
rect 597884 135922 597980 135978
rect 545484 135826 597980 135922
rect -1916 130350 66564 130446
rect -1916 130294 -860 130350
rect -804 130294 -736 130350
rect -680 130294 -612 130350
rect -556 130294 -488 130350
rect -432 130294 3250 130350
rect 3306 130294 3374 130350
rect 3430 130294 3498 130350
rect 3554 130294 3622 130350
rect 3678 130294 21250 130350
rect 21306 130294 21374 130350
rect 21430 130294 21498 130350
rect 21554 130294 21622 130350
rect 21678 130294 39250 130350
rect 39306 130294 39374 130350
rect 39430 130294 39498 130350
rect 39554 130294 39622 130350
rect 39678 130294 57250 130350
rect 57306 130294 57374 130350
rect 57430 130294 57498 130350
rect 57554 130294 57622 130350
rect 57678 130294 64518 130350
rect 64574 130294 64642 130350
rect 64698 130294 66564 130350
rect -1916 130226 66564 130294
rect -1916 130170 -860 130226
rect -804 130170 -736 130226
rect -680 130170 -612 130226
rect -556 130170 -488 130226
rect -432 130170 3250 130226
rect 3306 130170 3374 130226
rect 3430 130170 3498 130226
rect 3554 130170 3622 130226
rect 3678 130170 21250 130226
rect 21306 130170 21374 130226
rect 21430 130170 21498 130226
rect 21554 130170 21622 130226
rect 21678 130170 39250 130226
rect 39306 130170 39374 130226
rect 39430 130170 39498 130226
rect 39554 130170 39622 130226
rect 39678 130170 57250 130226
rect 57306 130170 57374 130226
rect 57430 130170 57498 130226
rect 57554 130170 57622 130226
rect 57678 130170 64518 130226
rect 64574 130170 64642 130226
rect 64698 130170 66564 130226
rect -1916 130102 66564 130170
rect -1916 130046 -860 130102
rect -804 130046 -736 130102
rect -680 130046 -612 130102
rect -556 130046 -488 130102
rect -432 130046 3250 130102
rect 3306 130046 3374 130102
rect 3430 130046 3498 130102
rect 3554 130046 3622 130102
rect 3678 130046 21250 130102
rect 21306 130046 21374 130102
rect 21430 130046 21498 130102
rect 21554 130046 21622 130102
rect 21678 130046 39250 130102
rect 39306 130046 39374 130102
rect 39430 130046 39498 130102
rect 39554 130046 39622 130102
rect 39678 130046 57250 130102
rect 57306 130046 57374 130102
rect 57430 130046 57498 130102
rect 57554 130046 57622 130102
rect 57678 130046 64518 130102
rect 64574 130046 64642 130102
rect 64698 130046 66564 130102
rect -1916 129978 66564 130046
rect -1916 129922 -860 129978
rect -804 129922 -736 129978
rect -680 129922 -612 129978
rect -556 129922 -488 129978
rect -432 129922 3250 129978
rect 3306 129922 3374 129978
rect 3430 129922 3498 129978
rect 3554 129922 3622 129978
rect 3678 129922 21250 129978
rect 21306 129922 21374 129978
rect 21430 129922 21498 129978
rect 21554 129922 21622 129978
rect 21678 129922 39250 129978
rect 39306 129922 39374 129978
rect 39430 129922 39498 129978
rect 39554 129922 39622 129978
rect 39678 129922 57250 129978
rect 57306 129922 57374 129978
rect 57430 129922 57498 129978
rect 57554 129922 57622 129978
rect 57678 129922 64518 129978
rect 64574 129922 64642 129978
rect 64698 129922 66564 129978
rect -1916 129826 66564 129922
rect 239468 130412 350740 130446
rect 239468 130356 284022 130412
rect 284078 130356 284146 130412
rect 284202 130356 284270 130412
rect 284326 130356 284394 130412
rect 284450 130356 284518 130412
rect 284574 130356 284642 130412
rect 284698 130356 284766 130412
rect 284822 130356 284890 130412
rect 284946 130356 285014 130412
rect 285070 130356 285138 130412
rect 285194 130356 304022 130412
rect 304078 130356 304146 130412
rect 304202 130356 304270 130412
rect 304326 130356 304394 130412
rect 304450 130356 304518 130412
rect 304574 130356 304642 130412
rect 304698 130356 304766 130412
rect 304822 130356 304890 130412
rect 304946 130356 305014 130412
rect 305070 130356 305138 130412
rect 305194 130356 350740 130412
rect 239468 130350 350740 130356
rect 239468 130294 255250 130350
rect 255306 130294 255374 130350
rect 255430 130294 255498 130350
rect 255554 130294 255622 130350
rect 255678 130294 273250 130350
rect 273306 130294 273374 130350
rect 273430 130294 273498 130350
rect 273554 130294 273622 130350
rect 273678 130294 327250 130350
rect 327306 130294 327374 130350
rect 327430 130294 327498 130350
rect 327554 130294 327622 130350
rect 327678 130294 345250 130350
rect 345306 130294 345374 130350
rect 345430 130294 345498 130350
rect 345554 130294 345622 130350
rect 345678 130294 350740 130350
rect 239468 130288 350740 130294
rect 239468 130232 284022 130288
rect 284078 130232 284146 130288
rect 284202 130232 284270 130288
rect 284326 130232 284394 130288
rect 284450 130232 284518 130288
rect 284574 130232 284642 130288
rect 284698 130232 284766 130288
rect 284822 130232 284890 130288
rect 284946 130232 285014 130288
rect 285070 130232 285138 130288
rect 285194 130232 304022 130288
rect 304078 130232 304146 130288
rect 304202 130232 304270 130288
rect 304326 130232 304394 130288
rect 304450 130232 304518 130288
rect 304574 130232 304642 130288
rect 304698 130232 304766 130288
rect 304822 130232 304890 130288
rect 304946 130232 305014 130288
rect 305070 130232 305138 130288
rect 305194 130232 350740 130288
rect 239468 130226 350740 130232
rect 239468 130170 255250 130226
rect 255306 130170 255374 130226
rect 255430 130170 255498 130226
rect 255554 130170 255622 130226
rect 255678 130170 273250 130226
rect 273306 130170 273374 130226
rect 273430 130170 273498 130226
rect 273554 130170 273622 130226
rect 273678 130170 327250 130226
rect 327306 130170 327374 130226
rect 327430 130170 327498 130226
rect 327554 130170 327622 130226
rect 327678 130170 345250 130226
rect 345306 130170 345374 130226
rect 345430 130170 345498 130226
rect 345554 130170 345622 130226
rect 345678 130170 350740 130226
rect 239468 130164 350740 130170
rect 239468 130108 284022 130164
rect 284078 130108 284146 130164
rect 284202 130108 284270 130164
rect 284326 130108 284394 130164
rect 284450 130108 284518 130164
rect 284574 130108 284642 130164
rect 284698 130108 284766 130164
rect 284822 130108 284890 130164
rect 284946 130108 285014 130164
rect 285070 130108 285138 130164
rect 285194 130108 304022 130164
rect 304078 130108 304146 130164
rect 304202 130108 304270 130164
rect 304326 130108 304394 130164
rect 304450 130108 304518 130164
rect 304574 130108 304642 130164
rect 304698 130108 304766 130164
rect 304822 130108 304890 130164
rect 304946 130108 305014 130164
rect 305070 130108 305138 130164
rect 305194 130108 350740 130164
rect 239468 130102 350740 130108
rect 239468 130046 255250 130102
rect 255306 130046 255374 130102
rect 255430 130046 255498 130102
rect 255554 130046 255622 130102
rect 255678 130046 273250 130102
rect 273306 130046 273374 130102
rect 273430 130046 273498 130102
rect 273554 130046 273622 130102
rect 273678 130046 327250 130102
rect 327306 130046 327374 130102
rect 327430 130046 327498 130102
rect 327554 130046 327622 130102
rect 327678 130046 345250 130102
rect 345306 130046 345374 130102
rect 345430 130046 345498 130102
rect 345554 130046 345622 130102
rect 345678 130046 350740 130102
rect 239468 130040 350740 130046
rect 239468 129984 284022 130040
rect 284078 129984 284146 130040
rect 284202 129984 284270 130040
rect 284326 129984 284394 130040
rect 284450 129984 284518 130040
rect 284574 129984 284642 130040
rect 284698 129984 284766 130040
rect 284822 129984 284890 130040
rect 284946 129984 285014 130040
rect 285070 129984 285138 130040
rect 285194 129984 304022 130040
rect 304078 129984 304146 130040
rect 304202 129984 304270 130040
rect 304326 129984 304394 130040
rect 304450 129984 304518 130040
rect 304574 129984 304642 130040
rect 304698 129984 304766 130040
rect 304822 129984 304890 130040
rect 304946 129984 305014 130040
rect 305070 129984 305138 130040
rect 305194 129984 350740 130040
rect 239468 129978 350740 129984
rect 239468 129922 255250 129978
rect 255306 129922 255374 129978
rect 255430 129922 255498 129978
rect 255554 129922 255622 129978
rect 255678 129922 273250 129978
rect 273306 129922 273374 129978
rect 273430 129922 273498 129978
rect 273554 129922 273622 129978
rect 273678 129922 327250 129978
rect 327306 129922 327374 129978
rect 327430 129922 327498 129978
rect 327554 129922 327622 129978
rect 327678 129922 345250 129978
rect 345306 129922 345374 129978
rect 345430 129922 345498 129978
rect 345554 129922 345622 129978
rect 345678 129922 350740 129978
rect 239468 129916 350740 129922
rect 239468 129860 284022 129916
rect 284078 129860 284146 129916
rect 284202 129860 284270 129916
rect 284326 129860 284394 129916
rect 284450 129860 284518 129916
rect 284574 129860 284642 129916
rect 284698 129860 284766 129916
rect 284822 129860 284890 129916
rect 284946 129860 285014 129916
rect 285070 129860 285138 129916
rect 285194 129860 304022 129916
rect 304078 129860 304146 129916
rect 304202 129860 304270 129916
rect 304326 129860 304394 129916
rect 304450 129860 304518 129916
rect 304574 129860 304642 129916
rect 304698 129860 304766 129916
rect 304822 129860 304890 129916
rect 304946 129860 305014 129916
rect 305070 129860 305138 129916
rect 305194 129860 350740 129916
rect 239468 129826 350740 129860
rect 545484 130350 597980 130446
rect 545484 130294 561250 130350
rect 561306 130294 561374 130350
rect 561430 130294 561498 130350
rect 561554 130294 561622 130350
rect 561678 130294 579250 130350
rect 579306 130294 579374 130350
rect 579430 130294 579498 130350
rect 579554 130294 579622 130350
rect 579678 130294 596496 130350
rect 596552 130294 596620 130350
rect 596676 130294 596744 130350
rect 596800 130294 596868 130350
rect 596924 130294 597980 130350
rect 545484 130226 597980 130294
rect 545484 130170 561250 130226
rect 561306 130170 561374 130226
rect 561430 130170 561498 130226
rect 561554 130170 561622 130226
rect 561678 130170 579250 130226
rect 579306 130170 579374 130226
rect 579430 130170 579498 130226
rect 579554 130170 579622 130226
rect 579678 130170 596496 130226
rect 596552 130170 596620 130226
rect 596676 130170 596744 130226
rect 596800 130170 596868 130226
rect 596924 130170 597980 130226
rect 545484 130102 597980 130170
rect 545484 130046 561250 130102
rect 561306 130046 561374 130102
rect 561430 130046 561498 130102
rect 561554 130046 561622 130102
rect 561678 130046 579250 130102
rect 579306 130046 579374 130102
rect 579430 130046 579498 130102
rect 579554 130046 579622 130102
rect 579678 130046 596496 130102
rect 596552 130046 596620 130102
rect 596676 130046 596744 130102
rect 596800 130046 596868 130102
rect 596924 130046 597980 130102
rect 545484 129978 597980 130046
rect 545484 129922 561250 129978
rect 561306 129922 561374 129978
rect 561430 129922 561498 129978
rect 561554 129922 561622 129978
rect 561678 129922 579250 129978
rect 579306 129922 579374 129978
rect 579430 129922 579498 129978
rect 579554 129922 579622 129978
rect 579678 129922 596496 129978
rect 596552 129922 596620 129978
rect 596676 129922 596744 129978
rect 596800 129922 596868 129978
rect 596924 129922 597980 129978
rect 545484 129826 597980 129922
rect -1916 118350 66564 118446
rect -1916 118294 -1820 118350
rect -1764 118294 -1696 118350
rect -1640 118294 -1572 118350
rect -1516 118294 -1448 118350
rect -1392 118294 6970 118350
rect 7026 118294 7094 118350
rect 7150 118294 7218 118350
rect 7274 118294 7342 118350
rect 7398 118294 24970 118350
rect 25026 118294 25094 118350
rect 25150 118294 25218 118350
rect 25274 118294 25342 118350
rect 25398 118294 42970 118350
rect 43026 118294 43094 118350
rect 43150 118294 43218 118350
rect 43274 118294 43342 118350
rect 43398 118294 66564 118350
rect -1916 118226 66564 118294
rect -1916 118170 -1820 118226
rect -1764 118170 -1696 118226
rect -1640 118170 -1572 118226
rect -1516 118170 -1448 118226
rect -1392 118170 6970 118226
rect 7026 118170 7094 118226
rect 7150 118170 7218 118226
rect 7274 118170 7342 118226
rect 7398 118170 24970 118226
rect 25026 118170 25094 118226
rect 25150 118170 25218 118226
rect 25274 118170 25342 118226
rect 25398 118170 42970 118226
rect 43026 118170 43094 118226
rect 43150 118170 43218 118226
rect 43274 118170 43342 118226
rect 43398 118170 66564 118226
rect -1916 118102 66564 118170
rect -1916 118046 -1820 118102
rect -1764 118046 -1696 118102
rect -1640 118046 -1572 118102
rect -1516 118046 -1448 118102
rect -1392 118046 6970 118102
rect 7026 118046 7094 118102
rect 7150 118046 7218 118102
rect 7274 118046 7342 118102
rect 7398 118046 24970 118102
rect 25026 118046 25094 118102
rect 25150 118046 25218 118102
rect 25274 118046 25342 118102
rect 25398 118046 42970 118102
rect 43026 118046 43094 118102
rect 43150 118046 43218 118102
rect 43274 118046 43342 118102
rect 43398 118046 66564 118102
rect -1916 117978 66564 118046
rect -1916 117922 -1820 117978
rect -1764 117922 -1696 117978
rect -1640 117922 -1572 117978
rect -1516 117922 -1448 117978
rect -1392 117922 6970 117978
rect 7026 117922 7094 117978
rect 7150 117922 7218 117978
rect 7274 117922 7342 117978
rect 7398 117922 24970 117978
rect 25026 117922 25094 117978
rect 25150 117922 25218 117978
rect 25274 117922 25342 117978
rect 25398 117922 42970 117978
rect 43026 117922 43094 117978
rect 43150 117922 43218 117978
rect 43274 117922 43342 117978
rect 43398 117922 66564 117978
rect -1916 117826 66564 117922
rect 239468 118412 350740 118446
rect 239468 118356 294022 118412
rect 294078 118356 294146 118412
rect 294202 118356 294270 118412
rect 294326 118356 294394 118412
rect 294450 118356 294518 118412
rect 294574 118356 294642 118412
rect 294698 118356 294766 118412
rect 294822 118356 294890 118412
rect 294946 118356 295014 118412
rect 295070 118356 295138 118412
rect 295194 118356 314022 118412
rect 314078 118356 314146 118412
rect 314202 118356 314270 118412
rect 314326 118356 314394 118412
rect 314450 118356 314518 118412
rect 314574 118356 314642 118412
rect 314698 118356 314766 118412
rect 314822 118356 314890 118412
rect 314946 118356 315014 118412
rect 315070 118356 315138 118412
rect 315194 118356 350740 118412
rect 239468 118350 350740 118356
rect 239468 118294 240970 118350
rect 241026 118294 241094 118350
rect 241150 118294 241218 118350
rect 241274 118294 241342 118350
rect 241398 118294 258970 118350
rect 259026 118294 259094 118350
rect 259150 118294 259218 118350
rect 259274 118294 259342 118350
rect 259398 118294 276970 118350
rect 277026 118294 277094 118350
rect 277150 118294 277218 118350
rect 277274 118294 277342 118350
rect 277398 118294 330970 118350
rect 331026 118294 331094 118350
rect 331150 118294 331218 118350
rect 331274 118294 331342 118350
rect 331398 118294 348970 118350
rect 349026 118294 349094 118350
rect 349150 118294 349218 118350
rect 349274 118294 349342 118350
rect 349398 118294 350740 118350
rect 239468 118288 350740 118294
rect 239468 118232 294022 118288
rect 294078 118232 294146 118288
rect 294202 118232 294270 118288
rect 294326 118232 294394 118288
rect 294450 118232 294518 118288
rect 294574 118232 294642 118288
rect 294698 118232 294766 118288
rect 294822 118232 294890 118288
rect 294946 118232 295014 118288
rect 295070 118232 295138 118288
rect 295194 118232 314022 118288
rect 314078 118232 314146 118288
rect 314202 118232 314270 118288
rect 314326 118232 314394 118288
rect 314450 118232 314518 118288
rect 314574 118232 314642 118288
rect 314698 118232 314766 118288
rect 314822 118232 314890 118288
rect 314946 118232 315014 118288
rect 315070 118232 315138 118288
rect 315194 118232 350740 118288
rect 239468 118226 350740 118232
rect 239468 118170 240970 118226
rect 241026 118170 241094 118226
rect 241150 118170 241218 118226
rect 241274 118170 241342 118226
rect 241398 118170 258970 118226
rect 259026 118170 259094 118226
rect 259150 118170 259218 118226
rect 259274 118170 259342 118226
rect 259398 118170 276970 118226
rect 277026 118170 277094 118226
rect 277150 118170 277218 118226
rect 277274 118170 277342 118226
rect 277398 118170 330970 118226
rect 331026 118170 331094 118226
rect 331150 118170 331218 118226
rect 331274 118170 331342 118226
rect 331398 118170 348970 118226
rect 349026 118170 349094 118226
rect 349150 118170 349218 118226
rect 349274 118170 349342 118226
rect 349398 118170 350740 118226
rect 239468 118164 350740 118170
rect 239468 118108 294022 118164
rect 294078 118108 294146 118164
rect 294202 118108 294270 118164
rect 294326 118108 294394 118164
rect 294450 118108 294518 118164
rect 294574 118108 294642 118164
rect 294698 118108 294766 118164
rect 294822 118108 294890 118164
rect 294946 118108 295014 118164
rect 295070 118108 295138 118164
rect 295194 118108 314022 118164
rect 314078 118108 314146 118164
rect 314202 118108 314270 118164
rect 314326 118108 314394 118164
rect 314450 118108 314518 118164
rect 314574 118108 314642 118164
rect 314698 118108 314766 118164
rect 314822 118108 314890 118164
rect 314946 118108 315014 118164
rect 315070 118108 315138 118164
rect 315194 118108 350740 118164
rect 239468 118102 350740 118108
rect 239468 118046 240970 118102
rect 241026 118046 241094 118102
rect 241150 118046 241218 118102
rect 241274 118046 241342 118102
rect 241398 118046 258970 118102
rect 259026 118046 259094 118102
rect 259150 118046 259218 118102
rect 259274 118046 259342 118102
rect 259398 118046 276970 118102
rect 277026 118046 277094 118102
rect 277150 118046 277218 118102
rect 277274 118046 277342 118102
rect 277398 118046 330970 118102
rect 331026 118046 331094 118102
rect 331150 118046 331218 118102
rect 331274 118046 331342 118102
rect 331398 118046 348970 118102
rect 349026 118046 349094 118102
rect 349150 118046 349218 118102
rect 349274 118046 349342 118102
rect 349398 118046 350740 118102
rect 239468 118040 350740 118046
rect 239468 117984 294022 118040
rect 294078 117984 294146 118040
rect 294202 117984 294270 118040
rect 294326 117984 294394 118040
rect 294450 117984 294518 118040
rect 294574 117984 294642 118040
rect 294698 117984 294766 118040
rect 294822 117984 294890 118040
rect 294946 117984 295014 118040
rect 295070 117984 295138 118040
rect 295194 117984 314022 118040
rect 314078 117984 314146 118040
rect 314202 117984 314270 118040
rect 314326 117984 314394 118040
rect 314450 117984 314518 118040
rect 314574 117984 314642 118040
rect 314698 117984 314766 118040
rect 314822 117984 314890 118040
rect 314946 117984 315014 118040
rect 315070 117984 315138 118040
rect 315194 117984 350740 118040
rect 239468 117978 350740 117984
rect 239468 117922 240970 117978
rect 241026 117922 241094 117978
rect 241150 117922 241218 117978
rect 241274 117922 241342 117978
rect 241398 117922 258970 117978
rect 259026 117922 259094 117978
rect 259150 117922 259218 117978
rect 259274 117922 259342 117978
rect 259398 117922 276970 117978
rect 277026 117922 277094 117978
rect 277150 117922 277218 117978
rect 277274 117922 277342 117978
rect 277398 117922 330970 117978
rect 331026 117922 331094 117978
rect 331150 117922 331218 117978
rect 331274 117922 331342 117978
rect 331398 117922 348970 117978
rect 349026 117922 349094 117978
rect 349150 117922 349218 117978
rect 349274 117922 349342 117978
rect 349398 117922 350740 117978
rect 239468 117916 350740 117922
rect 239468 117860 294022 117916
rect 294078 117860 294146 117916
rect 294202 117860 294270 117916
rect 294326 117860 294394 117916
rect 294450 117860 294518 117916
rect 294574 117860 294642 117916
rect 294698 117860 294766 117916
rect 294822 117860 294890 117916
rect 294946 117860 295014 117916
rect 295070 117860 295138 117916
rect 295194 117860 314022 117916
rect 314078 117860 314146 117916
rect 314202 117860 314270 117916
rect 314326 117860 314394 117916
rect 314450 117860 314518 117916
rect 314574 117860 314642 117916
rect 314698 117860 314766 117916
rect 314822 117860 314890 117916
rect 314946 117860 315014 117916
rect 315070 117860 315138 117916
rect 315194 117860 350740 117916
rect 239468 117826 350740 117860
rect 545484 118350 597980 118446
rect 545484 118294 564970 118350
rect 565026 118294 565094 118350
rect 565150 118294 565218 118350
rect 565274 118294 565342 118350
rect 565398 118294 582970 118350
rect 583026 118294 583094 118350
rect 583150 118294 583218 118350
rect 583274 118294 583342 118350
rect 583398 118294 597456 118350
rect 597512 118294 597580 118350
rect 597636 118294 597704 118350
rect 597760 118294 597828 118350
rect 597884 118294 597980 118350
rect 545484 118226 597980 118294
rect 545484 118170 564970 118226
rect 565026 118170 565094 118226
rect 565150 118170 565218 118226
rect 565274 118170 565342 118226
rect 565398 118170 582970 118226
rect 583026 118170 583094 118226
rect 583150 118170 583218 118226
rect 583274 118170 583342 118226
rect 583398 118170 597456 118226
rect 597512 118170 597580 118226
rect 597636 118170 597704 118226
rect 597760 118170 597828 118226
rect 597884 118170 597980 118226
rect 545484 118102 597980 118170
rect 545484 118046 564970 118102
rect 565026 118046 565094 118102
rect 565150 118046 565218 118102
rect 565274 118046 565342 118102
rect 565398 118046 582970 118102
rect 583026 118046 583094 118102
rect 583150 118046 583218 118102
rect 583274 118046 583342 118102
rect 583398 118046 597456 118102
rect 597512 118046 597580 118102
rect 597636 118046 597704 118102
rect 597760 118046 597828 118102
rect 597884 118046 597980 118102
rect 545484 117978 597980 118046
rect 545484 117922 564970 117978
rect 565026 117922 565094 117978
rect 565150 117922 565218 117978
rect 565274 117922 565342 117978
rect 565398 117922 582970 117978
rect 583026 117922 583094 117978
rect 583150 117922 583218 117978
rect 583274 117922 583342 117978
rect 583398 117922 597456 117978
rect 597512 117922 597580 117978
rect 597636 117922 597704 117978
rect 597760 117922 597828 117978
rect 597884 117922 597980 117978
rect 545484 117826 597980 117922
rect -1916 112350 66564 112446
rect -1916 112294 -860 112350
rect -804 112294 -736 112350
rect -680 112294 -612 112350
rect -556 112294 -488 112350
rect -432 112294 3250 112350
rect 3306 112294 3374 112350
rect 3430 112294 3498 112350
rect 3554 112294 3622 112350
rect 3678 112294 21250 112350
rect 21306 112294 21374 112350
rect 21430 112294 21498 112350
rect 21554 112294 21622 112350
rect 21678 112294 39250 112350
rect 39306 112294 39374 112350
rect 39430 112294 39498 112350
rect 39554 112294 39622 112350
rect 39678 112294 57250 112350
rect 57306 112294 57374 112350
rect 57430 112294 57498 112350
rect 57554 112294 57622 112350
rect 57678 112294 64518 112350
rect 64574 112294 64642 112350
rect 64698 112294 66564 112350
rect -1916 112226 66564 112294
rect -1916 112170 -860 112226
rect -804 112170 -736 112226
rect -680 112170 -612 112226
rect -556 112170 -488 112226
rect -432 112170 3250 112226
rect 3306 112170 3374 112226
rect 3430 112170 3498 112226
rect 3554 112170 3622 112226
rect 3678 112170 21250 112226
rect 21306 112170 21374 112226
rect 21430 112170 21498 112226
rect 21554 112170 21622 112226
rect 21678 112170 39250 112226
rect 39306 112170 39374 112226
rect 39430 112170 39498 112226
rect 39554 112170 39622 112226
rect 39678 112170 57250 112226
rect 57306 112170 57374 112226
rect 57430 112170 57498 112226
rect 57554 112170 57622 112226
rect 57678 112170 64518 112226
rect 64574 112170 64642 112226
rect 64698 112170 66564 112226
rect -1916 112102 66564 112170
rect -1916 112046 -860 112102
rect -804 112046 -736 112102
rect -680 112046 -612 112102
rect -556 112046 -488 112102
rect -432 112046 3250 112102
rect 3306 112046 3374 112102
rect 3430 112046 3498 112102
rect 3554 112046 3622 112102
rect 3678 112046 21250 112102
rect 21306 112046 21374 112102
rect 21430 112046 21498 112102
rect 21554 112046 21622 112102
rect 21678 112046 39250 112102
rect 39306 112046 39374 112102
rect 39430 112046 39498 112102
rect 39554 112046 39622 112102
rect 39678 112046 57250 112102
rect 57306 112046 57374 112102
rect 57430 112046 57498 112102
rect 57554 112046 57622 112102
rect 57678 112046 64518 112102
rect 64574 112046 64642 112102
rect 64698 112046 66564 112102
rect -1916 111978 66564 112046
rect -1916 111922 -860 111978
rect -804 111922 -736 111978
rect -680 111922 -612 111978
rect -556 111922 -488 111978
rect -432 111922 3250 111978
rect 3306 111922 3374 111978
rect 3430 111922 3498 111978
rect 3554 111922 3622 111978
rect 3678 111922 21250 111978
rect 21306 111922 21374 111978
rect 21430 111922 21498 111978
rect 21554 111922 21622 111978
rect 21678 111922 39250 111978
rect 39306 111922 39374 111978
rect 39430 111922 39498 111978
rect 39554 111922 39622 111978
rect 39678 111922 57250 111978
rect 57306 111922 57374 111978
rect 57430 111922 57498 111978
rect 57554 111922 57622 111978
rect 57678 111922 64518 111978
rect 64574 111922 64642 111978
rect 64698 111922 66564 111978
rect -1916 111826 66564 111922
rect 239468 112412 350740 112446
rect 239468 112356 284022 112412
rect 284078 112356 284146 112412
rect 284202 112356 284270 112412
rect 284326 112356 284394 112412
rect 284450 112356 284518 112412
rect 284574 112356 284642 112412
rect 284698 112356 284766 112412
rect 284822 112356 284890 112412
rect 284946 112356 285014 112412
rect 285070 112356 285138 112412
rect 285194 112356 304022 112412
rect 304078 112356 304146 112412
rect 304202 112356 304270 112412
rect 304326 112356 304394 112412
rect 304450 112356 304518 112412
rect 304574 112356 304642 112412
rect 304698 112356 304766 112412
rect 304822 112356 304890 112412
rect 304946 112356 305014 112412
rect 305070 112356 305138 112412
rect 305194 112356 350740 112412
rect 239468 112350 350740 112356
rect 239468 112294 255250 112350
rect 255306 112294 255374 112350
rect 255430 112294 255498 112350
rect 255554 112294 255622 112350
rect 255678 112294 273250 112350
rect 273306 112294 273374 112350
rect 273430 112294 273498 112350
rect 273554 112294 273622 112350
rect 273678 112294 327250 112350
rect 327306 112294 327374 112350
rect 327430 112294 327498 112350
rect 327554 112294 327622 112350
rect 327678 112294 345250 112350
rect 345306 112294 345374 112350
rect 345430 112294 345498 112350
rect 345554 112294 345622 112350
rect 345678 112294 350740 112350
rect 239468 112288 350740 112294
rect 239468 112232 284022 112288
rect 284078 112232 284146 112288
rect 284202 112232 284270 112288
rect 284326 112232 284394 112288
rect 284450 112232 284518 112288
rect 284574 112232 284642 112288
rect 284698 112232 284766 112288
rect 284822 112232 284890 112288
rect 284946 112232 285014 112288
rect 285070 112232 285138 112288
rect 285194 112232 304022 112288
rect 304078 112232 304146 112288
rect 304202 112232 304270 112288
rect 304326 112232 304394 112288
rect 304450 112232 304518 112288
rect 304574 112232 304642 112288
rect 304698 112232 304766 112288
rect 304822 112232 304890 112288
rect 304946 112232 305014 112288
rect 305070 112232 305138 112288
rect 305194 112232 350740 112288
rect 239468 112226 350740 112232
rect 239468 112170 255250 112226
rect 255306 112170 255374 112226
rect 255430 112170 255498 112226
rect 255554 112170 255622 112226
rect 255678 112170 273250 112226
rect 273306 112170 273374 112226
rect 273430 112170 273498 112226
rect 273554 112170 273622 112226
rect 273678 112170 327250 112226
rect 327306 112170 327374 112226
rect 327430 112170 327498 112226
rect 327554 112170 327622 112226
rect 327678 112170 345250 112226
rect 345306 112170 345374 112226
rect 345430 112170 345498 112226
rect 345554 112170 345622 112226
rect 345678 112170 350740 112226
rect 239468 112164 350740 112170
rect 239468 112108 284022 112164
rect 284078 112108 284146 112164
rect 284202 112108 284270 112164
rect 284326 112108 284394 112164
rect 284450 112108 284518 112164
rect 284574 112108 284642 112164
rect 284698 112108 284766 112164
rect 284822 112108 284890 112164
rect 284946 112108 285014 112164
rect 285070 112108 285138 112164
rect 285194 112108 304022 112164
rect 304078 112108 304146 112164
rect 304202 112108 304270 112164
rect 304326 112108 304394 112164
rect 304450 112108 304518 112164
rect 304574 112108 304642 112164
rect 304698 112108 304766 112164
rect 304822 112108 304890 112164
rect 304946 112108 305014 112164
rect 305070 112108 305138 112164
rect 305194 112108 350740 112164
rect 239468 112102 350740 112108
rect 239468 112046 255250 112102
rect 255306 112046 255374 112102
rect 255430 112046 255498 112102
rect 255554 112046 255622 112102
rect 255678 112046 273250 112102
rect 273306 112046 273374 112102
rect 273430 112046 273498 112102
rect 273554 112046 273622 112102
rect 273678 112046 327250 112102
rect 327306 112046 327374 112102
rect 327430 112046 327498 112102
rect 327554 112046 327622 112102
rect 327678 112046 345250 112102
rect 345306 112046 345374 112102
rect 345430 112046 345498 112102
rect 345554 112046 345622 112102
rect 345678 112046 350740 112102
rect 239468 112040 350740 112046
rect 239468 111984 284022 112040
rect 284078 111984 284146 112040
rect 284202 111984 284270 112040
rect 284326 111984 284394 112040
rect 284450 111984 284518 112040
rect 284574 111984 284642 112040
rect 284698 111984 284766 112040
rect 284822 111984 284890 112040
rect 284946 111984 285014 112040
rect 285070 111984 285138 112040
rect 285194 111984 304022 112040
rect 304078 111984 304146 112040
rect 304202 111984 304270 112040
rect 304326 111984 304394 112040
rect 304450 111984 304518 112040
rect 304574 111984 304642 112040
rect 304698 111984 304766 112040
rect 304822 111984 304890 112040
rect 304946 111984 305014 112040
rect 305070 111984 305138 112040
rect 305194 111984 350740 112040
rect 239468 111978 350740 111984
rect 239468 111922 255250 111978
rect 255306 111922 255374 111978
rect 255430 111922 255498 111978
rect 255554 111922 255622 111978
rect 255678 111922 273250 111978
rect 273306 111922 273374 111978
rect 273430 111922 273498 111978
rect 273554 111922 273622 111978
rect 273678 111922 327250 111978
rect 327306 111922 327374 111978
rect 327430 111922 327498 111978
rect 327554 111922 327622 111978
rect 327678 111922 345250 111978
rect 345306 111922 345374 111978
rect 345430 111922 345498 111978
rect 345554 111922 345622 111978
rect 345678 111922 350740 111978
rect 239468 111916 350740 111922
rect 239468 111860 284022 111916
rect 284078 111860 284146 111916
rect 284202 111860 284270 111916
rect 284326 111860 284394 111916
rect 284450 111860 284518 111916
rect 284574 111860 284642 111916
rect 284698 111860 284766 111916
rect 284822 111860 284890 111916
rect 284946 111860 285014 111916
rect 285070 111860 285138 111916
rect 285194 111860 304022 111916
rect 304078 111860 304146 111916
rect 304202 111860 304270 111916
rect 304326 111860 304394 111916
rect 304450 111860 304518 111916
rect 304574 111860 304642 111916
rect 304698 111860 304766 111916
rect 304822 111860 304890 111916
rect 304946 111860 305014 111916
rect 305070 111860 305138 111916
rect 305194 111860 350740 111916
rect 239468 111826 350740 111860
rect 545484 112350 597980 112446
rect 545484 112294 561250 112350
rect 561306 112294 561374 112350
rect 561430 112294 561498 112350
rect 561554 112294 561622 112350
rect 561678 112294 579250 112350
rect 579306 112294 579374 112350
rect 579430 112294 579498 112350
rect 579554 112294 579622 112350
rect 579678 112294 596496 112350
rect 596552 112294 596620 112350
rect 596676 112294 596744 112350
rect 596800 112294 596868 112350
rect 596924 112294 597980 112350
rect 545484 112226 597980 112294
rect 545484 112170 561250 112226
rect 561306 112170 561374 112226
rect 561430 112170 561498 112226
rect 561554 112170 561622 112226
rect 561678 112170 579250 112226
rect 579306 112170 579374 112226
rect 579430 112170 579498 112226
rect 579554 112170 579622 112226
rect 579678 112170 596496 112226
rect 596552 112170 596620 112226
rect 596676 112170 596744 112226
rect 596800 112170 596868 112226
rect 596924 112170 597980 112226
rect 545484 112102 597980 112170
rect 545484 112046 561250 112102
rect 561306 112046 561374 112102
rect 561430 112046 561498 112102
rect 561554 112046 561622 112102
rect 561678 112046 579250 112102
rect 579306 112046 579374 112102
rect 579430 112046 579498 112102
rect 579554 112046 579622 112102
rect 579678 112046 596496 112102
rect 596552 112046 596620 112102
rect 596676 112046 596744 112102
rect 596800 112046 596868 112102
rect 596924 112046 597980 112102
rect 545484 111978 597980 112046
rect 545484 111922 561250 111978
rect 561306 111922 561374 111978
rect 561430 111922 561498 111978
rect 561554 111922 561622 111978
rect 561678 111922 579250 111978
rect 579306 111922 579374 111978
rect 579430 111922 579498 111978
rect 579554 111922 579622 111978
rect 579678 111922 596496 111978
rect 596552 111922 596620 111978
rect 596676 111922 596744 111978
rect 596800 111922 596868 111978
rect 596924 111922 597980 111978
rect 545484 111826 597980 111922
rect -1916 100350 66564 100446
rect -1916 100294 -1820 100350
rect -1764 100294 -1696 100350
rect -1640 100294 -1572 100350
rect -1516 100294 -1448 100350
rect -1392 100294 6970 100350
rect 7026 100294 7094 100350
rect 7150 100294 7218 100350
rect 7274 100294 7342 100350
rect 7398 100294 24970 100350
rect 25026 100294 25094 100350
rect 25150 100294 25218 100350
rect 25274 100294 25342 100350
rect 25398 100294 42970 100350
rect 43026 100294 43094 100350
rect 43150 100294 43218 100350
rect 43274 100294 43342 100350
rect 43398 100294 66564 100350
rect -1916 100226 66564 100294
rect -1916 100170 -1820 100226
rect -1764 100170 -1696 100226
rect -1640 100170 -1572 100226
rect -1516 100170 -1448 100226
rect -1392 100170 6970 100226
rect 7026 100170 7094 100226
rect 7150 100170 7218 100226
rect 7274 100170 7342 100226
rect 7398 100170 24970 100226
rect 25026 100170 25094 100226
rect 25150 100170 25218 100226
rect 25274 100170 25342 100226
rect 25398 100170 42970 100226
rect 43026 100170 43094 100226
rect 43150 100170 43218 100226
rect 43274 100170 43342 100226
rect 43398 100170 66564 100226
rect -1916 100102 66564 100170
rect -1916 100046 -1820 100102
rect -1764 100046 -1696 100102
rect -1640 100046 -1572 100102
rect -1516 100046 -1448 100102
rect -1392 100046 6970 100102
rect 7026 100046 7094 100102
rect 7150 100046 7218 100102
rect 7274 100046 7342 100102
rect 7398 100046 24970 100102
rect 25026 100046 25094 100102
rect 25150 100046 25218 100102
rect 25274 100046 25342 100102
rect 25398 100046 42970 100102
rect 43026 100046 43094 100102
rect 43150 100046 43218 100102
rect 43274 100046 43342 100102
rect 43398 100046 66564 100102
rect -1916 99978 66564 100046
rect -1916 99922 -1820 99978
rect -1764 99922 -1696 99978
rect -1640 99922 -1572 99978
rect -1516 99922 -1448 99978
rect -1392 99922 6970 99978
rect 7026 99922 7094 99978
rect 7150 99922 7218 99978
rect 7274 99922 7342 99978
rect 7398 99922 24970 99978
rect 25026 99922 25094 99978
rect 25150 99922 25218 99978
rect 25274 99922 25342 99978
rect 25398 99922 42970 99978
rect 43026 99922 43094 99978
rect 43150 99922 43218 99978
rect 43274 99922 43342 99978
rect 43398 99922 66564 99978
rect -1916 99826 66564 99922
rect 239468 100412 350740 100446
rect 239468 100356 294022 100412
rect 294078 100356 294146 100412
rect 294202 100356 294270 100412
rect 294326 100356 294394 100412
rect 294450 100356 294518 100412
rect 294574 100356 294642 100412
rect 294698 100356 294766 100412
rect 294822 100356 294890 100412
rect 294946 100356 295014 100412
rect 295070 100356 295138 100412
rect 295194 100356 314022 100412
rect 314078 100356 314146 100412
rect 314202 100356 314270 100412
rect 314326 100356 314394 100412
rect 314450 100356 314518 100412
rect 314574 100356 314642 100412
rect 314698 100356 314766 100412
rect 314822 100356 314890 100412
rect 314946 100356 315014 100412
rect 315070 100356 315138 100412
rect 315194 100356 350740 100412
rect 239468 100350 350740 100356
rect 239468 100294 240970 100350
rect 241026 100294 241094 100350
rect 241150 100294 241218 100350
rect 241274 100294 241342 100350
rect 241398 100294 258970 100350
rect 259026 100294 259094 100350
rect 259150 100294 259218 100350
rect 259274 100294 259342 100350
rect 259398 100294 276970 100350
rect 277026 100294 277094 100350
rect 277150 100294 277218 100350
rect 277274 100294 277342 100350
rect 277398 100294 330970 100350
rect 331026 100294 331094 100350
rect 331150 100294 331218 100350
rect 331274 100294 331342 100350
rect 331398 100294 348970 100350
rect 349026 100294 349094 100350
rect 349150 100294 349218 100350
rect 349274 100294 349342 100350
rect 349398 100294 350740 100350
rect 239468 100288 350740 100294
rect 239468 100232 294022 100288
rect 294078 100232 294146 100288
rect 294202 100232 294270 100288
rect 294326 100232 294394 100288
rect 294450 100232 294518 100288
rect 294574 100232 294642 100288
rect 294698 100232 294766 100288
rect 294822 100232 294890 100288
rect 294946 100232 295014 100288
rect 295070 100232 295138 100288
rect 295194 100232 314022 100288
rect 314078 100232 314146 100288
rect 314202 100232 314270 100288
rect 314326 100232 314394 100288
rect 314450 100232 314518 100288
rect 314574 100232 314642 100288
rect 314698 100232 314766 100288
rect 314822 100232 314890 100288
rect 314946 100232 315014 100288
rect 315070 100232 315138 100288
rect 315194 100232 350740 100288
rect 239468 100226 350740 100232
rect 239468 100170 240970 100226
rect 241026 100170 241094 100226
rect 241150 100170 241218 100226
rect 241274 100170 241342 100226
rect 241398 100170 258970 100226
rect 259026 100170 259094 100226
rect 259150 100170 259218 100226
rect 259274 100170 259342 100226
rect 259398 100170 276970 100226
rect 277026 100170 277094 100226
rect 277150 100170 277218 100226
rect 277274 100170 277342 100226
rect 277398 100170 330970 100226
rect 331026 100170 331094 100226
rect 331150 100170 331218 100226
rect 331274 100170 331342 100226
rect 331398 100170 348970 100226
rect 349026 100170 349094 100226
rect 349150 100170 349218 100226
rect 349274 100170 349342 100226
rect 349398 100170 350740 100226
rect 239468 100164 350740 100170
rect 239468 100108 294022 100164
rect 294078 100108 294146 100164
rect 294202 100108 294270 100164
rect 294326 100108 294394 100164
rect 294450 100108 294518 100164
rect 294574 100108 294642 100164
rect 294698 100108 294766 100164
rect 294822 100108 294890 100164
rect 294946 100108 295014 100164
rect 295070 100108 295138 100164
rect 295194 100108 314022 100164
rect 314078 100108 314146 100164
rect 314202 100108 314270 100164
rect 314326 100108 314394 100164
rect 314450 100108 314518 100164
rect 314574 100108 314642 100164
rect 314698 100108 314766 100164
rect 314822 100108 314890 100164
rect 314946 100108 315014 100164
rect 315070 100108 315138 100164
rect 315194 100108 350740 100164
rect 239468 100102 350740 100108
rect 239468 100046 240970 100102
rect 241026 100046 241094 100102
rect 241150 100046 241218 100102
rect 241274 100046 241342 100102
rect 241398 100046 258970 100102
rect 259026 100046 259094 100102
rect 259150 100046 259218 100102
rect 259274 100046 259342 100102
rect 259398 100046 276970 100102
rect 277026 100046 277094 100102
rect 277150 100046 277218 100102
rect 277274 100046 277342 100102
rect 277398 100046 330970 100102
rect 331026 100046 331094 100102
rect 331150 100046 331218 100102
rect 331274 100046 331342 100102
rect 331398 100046 348970 100102
rect 349026 100046 349094 100102
rect 349150 100046 349218 100102
rect 349274 100046 349342 100102
rect 349398 100046 350740 100102
rect 239468 100040 350740 100046
rect 239468 99984 294022 100040
rect 294078 99984 294146 100040
rect 294202 99984 294270 100040
rect 294326 99984 294394 100040
rect 294450 99984 294518 100040
rect 294574 99984 294642 100040
rect 294698 99984 294766 100040
rect 294822 99984 294890 100040
rect 294946 99984 295014 100040
rect 295070 99984 295138 100040
rect 295194 99984 314022 100040
rect 314078 99984 314146 100040
rect 314202 99984 314270 100040
rect 314326 99984 314394 100040
rect 314450 99984 314518 100040
rect 314574 99984 314642 100040
rect 314698 99984 314766 100040
rect 314822 99984 314890 100040
rect 314946 99984 315014 100040
rect 315070 99984 315138 100040
rect 315194 99984 350740 100040
rect 239468 99978 350740 99984
rect 239468 99922 240970 99978
rect 241026 99922 241094 99978
rect 241150 99922 241218 99978
rect 241274 99922 241342 99978
rect 241398 99922 258970 99978
rect 259026 99922 259094 99978
rect 259150 99922 259218 99978
rect 259274 99922 259342 99978
rect 259398 99922 276970 99978
rect 277026 99922 277094 99978
rect 277150 99922 277218 99978
rect 277274 99922 277342 99978
rect 277398 99922 330970 99978
rect 331026 99922 331094 99978
rect 331150 99922 331218 99978
rect 331274 99922 331342 99978
rect 331398 99922 348970 99978
rect 349026 99922 349094 99978
rect 349150 99922 349218 99978
rect 349274 99922 349342 99978
rect 349398 99922 350740 99978
rect 239468 99916 350740 99922
rect 239468 99860 294022 99916
rect 294078 99860 294146 99916
rect 294202 99860 294270 99916
rect 294326 99860 294394 99916
rect 294450 99860 294518 99916
rect 294574 99860 294642 99916
rect 294698 99860 294766 99916
rect 294822 99860 294890 99916
rect 294946 99860 295014 99916
rect 295070 99860 295138 99916
rect 295194 99860 314022 99916
rect 314078 99860 314146 99916
rect 314202 99860 314270 99916
rect 314326 99860 314394 99916
rect 314450 99860 314518 99916
rect 314574 99860 314642 99916
rect 314698 99860 314766 99916
rect 314822 99860 314890 99916
rect 314946 99860 315014 99916
rect 315070 99860 315138 99916
rect 315194 99860 350740 99916
rect 239468 99826 350740 99860
rect 545484 100350 597980 100446
rect 545484 100294 564970 100350
rect 565026 100294 565094 100350
rect 565150 100294 565218 100350
rect 565274 100294 565342 100350
rect 565398 100294 582970 100350
rect 583026 100294 583094 100350
rect 583150 100294 583218 100350
rect 583274 100294 583342 100350
rect 583398 100294 597456 100350
rect 597512 100294 597580 100350
rect 597636 100294 597704 100350
rect 597760 100294 597828 100350
rect 597884 100294 597980 100350
rect 545484 100226 597980 100294
rect 545484 100170 564970 100226
rect 565026 100170 565094 100226
rect 565150 100170 565218 100226
rect 565274 100170 565342 100226
rect 565398 100170 582970 100226
rect 583026 100170 583094 100226
rect 583150 100170 583218 100226
rect 583274 100170 583342 100226
rect 583398 100170 597456 100226
rect 597512 100170 597580 100226
rect 597636 100170 597704 100226
rect 597760 100170 597828 100226
rect 597884 100170 597980 100226
rect 545484 100102 597980 100170
rect 545484 100046 564970 100102
rect 565026 100046 565094 100102
rect 565150 100046 565218 100102
rect 565274 100046 565342 100102
rect 565398 100046 582970 100102
rect 583026 100046 583094 100102
rect 583150 100046 583218 100102
rect 583274 100046 583342 100102
rect 583398 100046 597456 100102
rect 597512 100046 597580 100102
rect 597636 100046 597704 100102
rect 597760 100046 597828 100102
rect 597884 100046 597980 100102
rect 545484 99978 597980 100046
rect 545484 99922 564970 99978
rect 565026 99922 565094 99978
rect 565150 99922 565218 99978
rect 565274 99922 565342 99978
rect 565398 99922 582970 99978
rect 583026 99922 583094 99978
rect 583150 99922 583218 99978
rect 583274 99922 583342 99978
rect 583398 99922 597456 99978
rect 597512 99922 597580 99978
rect 597636 99922 597704 99978
rect 597760 99922 597828 99978
rect 597884 99922 597980 99978
rect 545484 99826 597980 99922
rect -1916 94350 66564 94446
rect -1916 94294 -860 94350
rect -804 94294 -736 94350
rect -680 94294 -612 94350
rect -556 94294 -488 94350
rect -432 94294 3250 94350
rect 3306 94294 3374 94350
rect 3430 94294 3498 94350
rect 3554 94294 3622 94350
rect 3678 94294 21250 94350
rect 21306 94294 21374 94350
rect 21430 94294 21498 94350
rect 21554 94294 21622 94350
rect 21678 94294 39250 94350
rect 39306 94294 39374 94350
rect 39430 94294 39498 94350
rect 39554 94294 39622 94350
rect 39678 94294 57250 94350
rect 57306 94294 57374 94350
rect 57430 94294 57498 94350
rect 57554 94294 57622 94350
rect 57678 94294 64518 94350
rect 64574 94294 64642 94350
rect 64698 94294 66564 94350
rect -1916 94226 66564 94294
rect -1916 94170 -860 94226
rect -804 94170 -736 94226
rect -680 94170 -612 94226
rect -556 94170 -488 94226
rect -432 94170 3250 94226
rect 3306 94170 3374 94226
rect 3430 94170 3498 94226
rect 3554 94170 3622 94226
rect 3678 94170 21250 94226
rect 21306 94170 21374 94226
rect 21430 94170 21498 94226
rect 21554 94170 21622 94226
rect 21678 94170 39250 94226
rect 39306 94170 39374 94226
rect 39430 94170 39498 94226
rect 39554 94170 39622 94226
rect 39678 94170 57250 94226
rect 57306 94170 57374 94226
rect 57430 94170 57498 94226
rect 57554 94170 57622 94226
rect 57678 94170 64518 94226
rect 64574 94170 64642 94226
rect 64698 94170 66564 94226
rect -1916 94102 66564 94170
rect -1916 94046 -860 94102
rect -804 94046 -736 94102
rect -680 94046 -612 94102
rect -556 94046 -488 94102
rect -432 94046 3250 94102
rect 3306 94046 3374 94102
rect 3430 94046 3498 94102
rect 3554 94046 3622 94102
rect 3678 94046 21250 94102
rect 21306 94046 21374 94102
rect 21430 94046 21498 94102
rect 21554 94046 21622 94102
rect 21678 94046 39250 94102
rect 39306 94046 39374 94102
rect 39430 94046 39498 94102
rect 39554 94046 39622 94102
rect 39678 94046 57250 94102
rect 57306 94046 57374 94102
rect 57430 94046 57498 94102
rect 57554 94046 57622 94102
rect 57678 94046 64518 94102
rect 64574 94046 64642 94102
rect 64698 94046 66564 94102
rect -1916 93978 66564 94046
rect -1916 93922 -860 93978
rect -804 93922 -736 93978
rect -680 93922 -612 93978
rect -556 93922 -488 93978
rect -432 93922 3250 93978
rect 3306 93922 3374 93978
rect 3430 93922 3498 93978
rect 3554 93922 3622 93978
rect 3678 93922 21250 93978
rect 21306 93922 21374 93978
rect 21430 93922 21498 93978
rect 21554 93922 21622 93978
rect 21678 93922 39250 93978
rect 39306 93922 39374 93978
rect 39430 93922 39498 93978
rect 39554 93922 39622 93978
rect 39678 93922 57250 93978
rect 57306 93922 57374 93978
rect 57430 93922 57498 93978
rect 57554 93922 57622 93978
rect 57678 93922 64518 93978
rect 64574 93922 64642 93978
rect 64698 93922 66564 93978
rect -1916 93826 66564 93922
rect 239468 94412 350740 94446
rect 239468 94356 284022 94412
rect 284078 94356 284146 94412
rect 284202 94356 284270 94412
rect 284326 94356 284394 94412
rect 284450 94356 284518 94412
rect 284574 94356 284642 94412
rect 284698 94356 284766 94412
rect 284822 94356 284890 94412
rect 284946 94356 285014 94412
rect 285070 94356 285138 94412
rect 285194 94356 304022 94412
rect 304078 94356 304146 94412
rect 304202 94356 304270 94412
rect 304326 94356 304394 94412
rect 304450 94356 304518 94412
rect 304574 94356 304642 94412
rect 304698 94356 304766 94412
rect 304822 94356 304890 94412
rect 304946 94356 305014 94412
rect 305070 94356 305138 94412
rect 305194 94356 350740 94412
rect 239468 94350 350740 94356
rect 239468 94294 255250 94350
rect 255306 94294 255374 94350
rect 255430 94294 255498 94350
rect 255554 94294 255622 94350
rect 255678 94294 273250 94350
rect 273306 94294 273374 94350
rect 273430 94294 273498 94350
rect 273554 94294 273622 94350
rect 273678 94294 327250 94350
rect 327306 94294 327374 94350
rect 327430 94294 327498 94350
rect 327554 94294 327622 94350
rect 327678 94294 345250 94350
rect 345306 94294 345374 94350
rect 345430 94294 345498 94350
rect 345554 94294 345622 94350
rect 345678 94294 350740 94350
rect 239468 94288 350740 94294
rect 239468 94232 284022 94288
rect 284078 94232 284146 94288
rect 284202 94232 284270 94288
rect 284326 94232 284394 94288
rect 284450 94232 284518 94288
rect 284574 94232 284642 94288
rect 284698 94232 284766 94288
rect 284822 94232 284890 94288
rect 284946 94232 285014 94288
rect 285070 94232 285138 94288
rect 285194 94232 304022 94288
rect 304078 94232 304146 94288
rect 304202 94232 304270 94288
rect 304326 94232 304394 94288
rect 304450 94232 304518 94288
rect 304574 94232 304642 94288
rect 304698 94232 304766 94288
rect 304822 94232 304890 94288
rect 304946 94232 305014 94288
rect 305070 94232 305138 94288
rect 305194 94232 350740 94288
rect 239468 94226 350740 94232
rect 239468 94170 255250 94226
rect 255306 94170 255374 94226
rect 255430 94170 255498 94226
rect 255554 94170 255622 94226
rect 255678 94170 273250 94226
rect 273306 94170 273374 94226
rect 273430 94170 273498 94226
rect 273554 94170 273622 94226
rect 273678 94170 327250 94226
rect 327306 94170 327374 94226
rect 327430 94170 327498 94226
rect 327554 94170 327622 94226
rect 327678 94170 345250 94226
rect 345306 94170 345374 94226
rect 345430 94170 345498 94226
rect 345554 94170 345622 94226
rect 345678 94170 350740 94226
rect 239468 94164 350740 94170
rect 239468 94108 284022 94164
rect 284078 94108 284146 94164
rect 284202 94108 284270 94164
rect 284326 94108 284394 94164
rect 284450 94108 284518 94164
rect 284574 94108 284642 94164
rect 284698 94108 284766 94164
rect 284822 94108 284890 94164
rect 284946 94108 285014 94164
rect 285070 94108 285138 94164
rect 285194 94108 304022 94164
rect 304078 94108 304146 94164
rect 304202 94108 304270 94164
rect 304326 94108 304394 94164
rect 304450 94108 304518 94164
rect 304574 94108 304642 94164
rect 304698 94108 304766 94164
rect 304822 94108 304890 94164
rect 304946 94108 305014 94164
rect 305070 94108 305138 94164
rect 305194 94108 350740 94164
rect 239468 94102 350740 94108
rect 239468 94046 255250 94102
rect 255306 94046 255374 94102
rect 255430 94046 255498 94102
rect 255554 94046 255622 94102
rect 255678 94046 273250 94102
rect 273306 94046 273374 94102
rect 273430 94046 273498 94102
rect 273554 94046 273622 94102
rect 273678 94046 327250 94102
rect 327306 94046 327374 94102
rect 327430 94046 327498 94102
rect 327554 94046 327622 94102
rect 327678 94046 345250 94102
rect 345306 94046 345374 94102
rect 345430 94046 345498 94102
rect 345554 94046 345622 94102
rect 345678 94046 350740 94102
rect 239468 94040 350740 94046
rect 239468 93984 284022 94040
rect 284078 93984 284146 94040
rect 284202 93984 284270 94040
rect 284326 93984 284394 94040
rect 284450 93984 284518 94040
rect 284574 93984 284642 94040
rect 284698 93984 284766 94040
rect 284822 93984 284890 94040
rect 284946 93984 285014 94040
rect 285070 93984 285138 94040
rect 285194 93984 304022 94040
rect 304078 93984 304146 94040
rect 304202 93984 304270 94040
rect 304326 93984 304394 94040
rect 304450 93984 304518 94040
rect 304574 93984 304642 94040
rect 304698 93984 304766 94040
rect 304822 93984 304890 94040
rect 304946 93984 305014 94040
rect 305070 93984 305138 94040
rect 305194 93984 350740 94040
rect 239468 93978 350740 93984
rect 239468 93922 255250 93978
rect 255306 93922 255374 93978
rect 255430 93922 255498 93978
rect 255554 93922 255622 93978
rect 255678 93922 273250 93978
rect 273306 93922 273374 93978
rect 273430 93922 273498 93978
rect 273554 93922 273622 93978
rect 273678 93922 327250 93978
rect 327306 93922 327374 93978
rect 327430 93922 327498 93978
rect 327554 93922 327622 93978
rect 327678 93922 345250 93978
rect 345306 93922 345374 93978
rect 345430 93922 345498 93978
rect 345554 93922 345622 93978
rect 345678 93922 350740 93978
rect 239468 93916 350740 93922
rect 239468 93860 284022 93916
rect 284078 93860 284146 93916
rect 284202 93860 284270 93916
rect 284326 93860 284394 93916
rect 284450 93860 284518 93916
rect 284574 93860 284642 93916
rect 284698 93860 284766 93916
rect 284822 93860 284890 93916
rect 284946 93860 285014 93916
rect 285070 93860 285138 93916
rect 285194 93860 304022 93916
rect 304078 93860 304146 93916
rect 304202 93860 304270 93916
rect 304326 93860 304394 93916
rect 304450 93860 304518 93916
rect 304574 93860 304642 93916
rect 304698 93860 304766 93916
rect 304822 93860 304890 93916
rect 304946 93860 305014 93916
rect 305070 93860 305138 93916
rect 305194 93860 350740 93916
rect 239468 93826 350740 93860
rect 545484 94350 597980 94446
rect 545484 94294 561250 94350
rect 561306 94294 561374 94350
rect 561430 94294 561498 94350
rect 561554 94294 561622 94350
rect 561678 94294 579250 94350
rect 579306 94294 579374 94350
rect 579430 94294 579498 94350
rect 579554 94294 579622 94350
rect 579678 94294 596496 94350
rect 596552 94294 596620 94350
rect 596676 94294 596744 94350
rect 596800 94294 596868 94350
rect 596924 94294 597980 94350
rect 545484 94226 597980 94294
rect 545484 94170 561250 94226
rect 561306 94170 561374 94226
rect 561430 94170 561498 94226
rect 561554 94170 561622 94226
rect 561678 94170 579250 94226
rect 579306 94170 579374 94226
rect 579430 94170 579498 94226
rect 579554 94170 579622 94226
rect 579678 94170 596496 94226
rect 596552 94170 596620 94226
rect 596676 94170 596744 94226
rect 596800 94170 596868 94226
rect 596924 94170 597980 94226
rect 545484 94102 597980 94170
rect 545484 94046 561250 94102
rect 561306 94046 561374 94102
rect 561430 94046 561498 94102
rect 561554 94046 561622 94102
rect 561678 94046 579250 94102
rect 579306 94046 579374 94102
rect 579430 94046 579498 94102
rect 579554 94046 579622 94102
rect 579678 94046 596496 94102
rect 596552 94046 596620 94102
rect 596676 94046 596744 94102
rect 596800 94046 596868 94102
rect 596924 94046 597980 94102
rect 545484 93978 597980 94046
rect 545484 93922 561250 93978
rect 561306 93922 561374 93978
rect 561430 93922 561498 93978
rect 561554 93922 561622 93978
rect 561678 93922 579250 93978
rect 579306 93922 579374 93978
rect 579430 93922 579498 93978
rect 579554 93922 579622 93978
rect 579678 93922 596496 93978
rect 596552 93922 596620 93978
rect 596676 93922 596744 93978
rect 596800 93922 596868 93978
rect 596924 93922 597980 93978
rect 545484 93826 597980 93922
rect -1916 82350 66564 82446
rect -1916 82294 -1820 82350
rect -1764 82294 -1696 82350
rect -1640 82294 -1572 82350
rect -1516 82294 -1448 82350
rect -1392 82294 6970 82350
rect 7026 82294 7094 82350
rect 7150 82294 7218 82350
rect 7274 82294 7342 82350
rect 7398 82294 24970 82350
rect 25026 82294 25094 82350
rect 25150 82294 25218 82350
rect 25274 82294 25342 82350
rect 25398 82294 42970 82350
rect 43026 82294 43094 82350
rect 43150 82294 43218 82350
rect 43274 82294 43342 82350
rect 43398 82294 66564 82350
rect -1916 82226 66564 82294
rect -1916 82170 -1820 82226
rect -1764 82170 -1696 82226
rect -1640 82170 -1572 82226
rect -1516 82170 -1448 82226
rect -1392 82170 6970 82226
rect 7026 82170 7094 82226
rect 7150 82170 7218 82226
rect 7274 82170 7342 82226
rect 7398 82170 24970 82226
rect 25026 82170 25094 82226
rect 25150 82170 25218 82226
rect 25274 82170 25342 82226
rect 25398 82170 42970 82226
rect 43026 82170 43094 82226
rect 43150 82170 43218 82226
rect 43274 82170 43342 82226
rect 43398 82170 66564 82226
rect -1916 82102 66564 82170
rect -1916 82046 -1820 82102
rect -1764 82046 -1696 82102
rect -1640 82046 -1572 82102
rect -1516 82046 -1448 82102
rect -1392 82046 6970 82102
rect 7026 82046 7094 82102
rect 7150 82046 7218 82102
rect 7274 82046 7342 82102
rect 7398 82046 24970 82102
rect 25026 82046 25094 82102
rect 25150 82046 25218 82102
rect 25274 82046 25342 82102
rect 25398 82046 42970 82102
rect 43026 82046 43094 82102
rect 43150 82046 43218 82102
rect 43274 82046 43342 82102
rect 43398 82046 66564 82102
rect -1916 81978 66564 82046
rect -1916 81922 -1820 81978
rect -1764 81922 -1696 81978
rect -1640 81922 -1572 81978
rect -1516 81922 -1448 81978
rect -1392 81922 6970 81978
rect 7026 81922 7094 81978
rect 7150 81922 7218 81978
rect 7274 81922 7342 81978
rect 7398 81922 24970 81978
rect 25026 81922 25094 81978
rect 25150 81922 25218 81978
rect 25274 81922 25342 81978
rect 25398 81922 42970 81978
rect 43026 81922 43094 81978
rect 43150 81922 43218 81978
rect 43274 81922 43342 81978
rect 43398 81922 66564 81978
rect -1916 81826 66564 81922
rect 239468 82412 350740 82446
rect 239468 82356 294022 82412
rect 294078 82356 294146 82412
rect 294202 82356 294270 82412
rect 294326 82356 294394 82412
rect 294450 82356 294518 82412
rect 294574 82356 294642 82412
rect 294698 82356 294766 82412
rect 294822 82356 294890 82412
rect 294946 82356 295014 82412
rect 295070 82356 295138 82412
rect 295194 82356 314022 82412
rect 314078 82356 314146 82412
rect 314202 82356 314270 82412
rect 314326 82356 314394 82412
rect 314450 82356 314518 82412
rect 314574 82356 314642 82412
rect 314698 82356 314766 82412
rect 314822 82356 314890 82412
rect 314946 82356 315014 82412
rect 315070 82356 315138 82412
rect 315194 82356 350740 82412
rect 239468 82350 350740 82356
rect 239468 82294 240970 82350
rect 241026 82294 241094 82350
rect 241150 82294 241218 82350
rect 241274 82294 241342 82350
rect 241398 82294 258970 82350
rect 259026 82294 259094 82350
rect 259150 82294 259218 82350
rect 259274 82294 259342 82350
rect 259398 82294 276970 82350
rect 277026 82294 277094 82350
rect 277150 82294 277218 82350
rect 277274 82294 277342 82350
rect 277398 82294 330970 82350
rect 331026 82294 331094 82350
rect 331150 82294 331218 82350
rect 331274 82294 331342 82350
rect 331398 82294 348970 82350
rect 349026 82294 349094 82350
rect 349150 82294 349218 82350
rect 349274 82294 349342 82350
rect 349398 82294 350740 82350
rect 239468 82288 350740 82294
rect 239468 82232 294022 82288
rect 294078 82232 294146 82288
rect 294202 82232 294270 82288
rect 294326 82232 294394 82288
rect 294450 82232 294518 82288
rect 294574 82232 294642 82288
rect 294698 82232 294766 82288
rect 294822 82232 294890 82288
rect 294946 82232 295014 82288
rect 295070 82232 295138 82288
rect 295194 82232 314022 82288
rect 314078 82232 314146 82288
rect 314202 82232 314270 82288
rect 314326 82232 314394 82288
rect 314450 82232 314518 82288
rect 314574 82232 314642 82288
rect 314698 82232 314766 82288
rect 314822 82232 314890 82288
rect 314946 82232 315014 82288
rect 315070 82232 315138 82288
rect 315194 82232 350740 82288
rect 239468 82226 350740 82232
rect 239468 82170 240970 82226
rect 241026 82170 241094 82226
rect 241150 82170 241218 82226
rect 241274 82170 241342 82226
rect 241398 82170 258970 82226
rect 259026 82170 259094 82226
rect 259150 82170 259218 82226
rect 259274 82170 259342 82226
rect 259398 82170 276970 82226
rect 277026 82170 277094 82226
rect 277150 82170 277218 82226
rect 277274 82170 277342 82226
rect 277398 82170 330970 82226
rect 331026 82170 331094 82226
rect 331150 82170 331218 82226
rect 331274 82170 331342 82226
rect 331398 82170 348970 82226
rect 349026 82170 349094 82226
rect 349150 82170 349218 82226
rect 349274 82170 349342 82226
rect 349398 82170 350740 82226
rect 239468 82164 350740 82170
rect 239468 82108 294022 82164
rect 294078 82108 294146 82164
rect 294202 82108 294270 82164
rect 294326 82108 294394 82164
rect 294450 82108 294518 82164
rect 294574 82108 294642 82164
rect 294698 82108 294766 82164
rect 294822 82108 294890 82164
rect 294946 82108 295014 82164
rect 295070 82108 295138 82164
rect 295194 82108 314022 82164
rect 314078 82108 314146 82164
rect 314202 82108 314270 82164
rect 314326 82108 314394 82164
rect 314450 82108 314518 82164
rect 314574 82108 314642 82164
rect 314698 82108 314766 82164
rect 314822 82108 314890 82164
rect 314946 82108 315014 82164
rect 315070 82108 315138 82164
rect 315194 82108 350740 82164
rect 239468 82102 350740 82108
rect 239468 82046 240970 82102
rect 241026 82046 241094 82102
rect 241150 82046 241218 82102
rect 241274 82046 241342 82102
rect 241398 82046 258970 82102
rect 259026 82046 259094 82102
rect 259150 82046 259218 82102
rect 259274 82046 259342 82102
rect 259398 82046 276970 82102
rect 277026 82046 277094 82102
rect 277150 82046 277218 82102
rect 277274 82046 277342 82102
rect 277398 82046 330970 82102
rect 331026 82046 331094 82102
rect 331150 82046 331218 82102
rect 331274 82046 331342 82102
rect 331398 82046 348970 82102
rect 349026 82046 349094 82102
rect 349150 82046 349218 82102
rect 349274 82046 349342 82102
rect 349398 82046 350740 82102
rect 239468 82040 350740 82046
rect 239468 81984 294022 82040
rect 294078 81984 294146 82040
rect 294202 81984 294270 82040
rect 294326 81984 294394 82040
rect 294450 81984 294518 82040
rect 294574 81984 294642 82040
rect 294698 81984 294766 82040
rect 294822 81984 294890 82040
rect 294946 81984 295014 82040
rect 295070 81984 295138 82040
rect 295194 81984 314022 82040
rect 314078 81984 314146 82040
rect 314202 81984 314270 82040
rect 314326 81984 314394 82040
rect 314450 81984 314518 82040
rect 314574 81984 314642 82040
rect 314698 81984 314766 82040
rect 314822 81984 314890 82040
rect 314946 81984 315014 82040
rect 315070 81984 315138 82040
rect 315194 81984 350740 82040
rect 239468 81978 350740 81984
rect 239468 81922 240970 81978
rect 241026 81922 241094 81978
rect 241150 81922 241218 81978
rect 241274 81922 241342 81978
rect 241398 81922 258970 81978
rect 259026 81922 259094 81978
rect 259150 81922 259218 81978
rect 259274 81922 259342 81978
rect 259398 81922 276970 81978
rect 277026 81922 277094 81978
rect 277150 81922 277218 81978
rect 277274 81922 277342 81978
rect 277398 81922 330970 81978
rect 331026 81922 331094 81978
rect 331150 81922 331218 81978
rect 331274 81922 331342 81978
rect 331398 81922 348970 81978
rect 349026 81922 349094 81978
rect 349150 81922 349218 81978
rect 349274 81922 349342 81978
rect 349398 81922 350740 81978
rect 239468 81916 350740 81922
rect 239468 81860 294022 81916
rect 294078 81860 294146 81916
rect 294202 81860 294270 81916
rect 294326 81860 294394 81916
rect 294450 81860 294518 81916
rect 294574 81860 294642 81916
rect 294698 81860 294766 81916
rect 294822 81860 294890 81916
rect 294946 81860 295014 81916
rect 295070 81860 295138 81916
rect 295194 81860 314022 81916
rect 314078 81860 314146 81916
rect 314202 81860 314270 81916
rect 314326 81860 314394 81916
rect 314450 81860 314518 81916
rect 314574 81860 314642 81916
rect 314698 81860 314766 81916
rect 314822 81860 314890 81916
rect 314946 81860 315014 81916
rect 315070 81860 315138 81916
rect 315194 81860 350740 81916
rect 239468 81826 350740 81860
rect 545484 82350 597980 82446
rect 545484 82294 564970 82350
rect 565026 82294 565094 82350
rect 565150 82294 565218 82350
rect 565274 82294 565342 82350
rect 565398 82294 582970 82350
rect 583026 82294 583094 82350
rect 583150 82294 583218 82350
rect 583274 82294 583342 82350
rect 583398 82294 597456 82350
rect 597512 82294 597580 82350
rect 597636 82294 597704 82350
rect 597760 82294 597828 82350
rect 597884 82294 597980 82350
rect 545484 82226 597980 82294
rect 545484 82170 564970 82226
rect 565026 82170 565094 82226
rect 565150 82170 565218 82226
rect 565274 82170 565342 82226
rect 565398 82170 582970 82226
rect 583026 82170 583094 82226
rect 583150 82170 583218 82226
rect 583274 82170 583342 82226
rect 583398 82170 597456 82226
rect 597512 82170 597580 82226
rect 597636 82170 597704 82226
rect 597760 82170 597828 82226
rect 597884 82170 597980 82226
rect 545484 82102 597980 82170
rect 545484 82046 564970 82102
rect 565026 82046 565094 82102
rect 565150 82046 565218 82102
rect 565274 82046 565342 82102
rect 565398 82046 582970 82102
rect 583026 82046 583094 82102
rect 583150 82046 583218 82102
rect 583274 82046 583342 82102
rect 583398 82046 597456 82102
rect 597512 82046 597580 82102
rect 597636 82046 597704 82102
rect 597760 82046 597828 82102
rect 597884 82046 597980 82102
rect 545484 81978 597980 82046
rect 545484 81922 564970 81978
rect 565026 81922 565094 81978
rect 565150 81922 565218 81978
rect 565274 81922 565342 81978
rect 565398 81922 582970 81978
rect 583026 81922 583094 81978
rect 583150 81922 583218 81978
rect 583274 81922 583342 81978
rect 583398 81922 597456 81978
rect 597512 81922 597580 81978
rect 597636 81922 597704 81978
rect 597760 81922 597828 81978
rect 597884 81922 597980 81978
rect 545484 81826 597980 81922
rect -1916 76350 66564 76446
rect -1916 76294 -860 76350
rect -804 76294 -736 76350
rect -680 76294 -612 76350
rect -556 76294 -488 76350
rect -432 76294 3250 76350
rect 3306 76294 3374 76350
rect 3430 76294 3498 76350
rect 3554 76294 3622 76350
rect 3678 76294 21250 76350
rect 21306 76294 21374 76350
rect 21430 76294 21498 76350
rect 21554 76294 21622 76350
rect 21678 76294 39250 76350
rect 39306 76294 39374 76350
rect 39430 76294 39498 76350
rect 39554 76294 39622 76350
rect 39678 76294 57250 76350
rect 57306 76294 57374 76350
rect 57430 76294 57498 76350
rect 57554 76294 57622 76350
rect 57678 76294 64518 76350
rect 64574 76294 64642 76350
rect 64698 76294 66564 76350
rect -1916 76226 66564 76294
rect -1916 76170 -860 76226
rect -804 76170 -736 76226
rect -680 76170 -612 76226
rect -556 76170 -488 76226
rect -432 76170 3250 76226
rect 3306 76170 3374 76226
rect 3430 76170 3498 76226
rect 3554 76170 3622 76226
rect 3678 76170 21250 76226
rect 21306 76170 21374 76226
rect 21430 76170 21498 76226
rect 21554 76170 21622 76226
rect 21678 76170 39250 76226
rect 39306 76170 39374 76226
rect 39430 76170 39498 76226
rect 39554 76170 39622 76226
rect 39678 76170 57250 76226
rect 57306 76170 57374 76226
rect 57430 76170 57498 76226
rect 57554 76170 57622 76226
rect 57678 76170 64518 76226
rect 64574 76170 64642 76226
rect 64698 76170 66564 76226
rect -1916 76102 66564 76170
rect -1916 76046 -860 76102
rect -804 76046 -736 76102
rect -680 76046 -612 76102
rect -556 76046 -488 76102
rect -432 76046 3250 76102
rect 3306 76046 3374 76102
rect 3430 76046 3498 76102
rect 3554 76046 3622 76102
rect 3678 76046 21250 76102
rect 21306 76046 21374 76102
rect 21430 76046 21498 76102
rect 21554 76046 21622 76102
rect 21678 76046 39250 76102
rect 39306 76046 39374 76102
rect 39430 76046 39498 76102
rect 39554 76046 39622 76102
rect 39678 76046 57250 76102
rect 57306 76046 57374 76102
rect 57430 76046 57498 76102
rect 57554 76046 57622 76102
rect 57678 76046 64518 76102
rect 64574 76046 64642 76102
rect 64698 76046 66564 76102
rect -1916 75978 66564 76046
rect -1916 75922 -860 75978
rect -804 75922 -736 75978
rect -680 75922 -612 75978
rect -556 75922 -488 75978
rect -432 75922 3250 75978
rect 3306 75922 3374 75978
rect 3430 75922 3498 75978
rect 3554 75922 3622 75978
rect 3678 75922 21250 75978
rect 21306 75922 21374 75978
rect 21430 75922 21498 75978
rect 21554 75922 21622 75978
rect 21678 75922 39250 75978
rect 39306 75922 39374 75978
rect 39430 75922 39498 75978
rect 39554 75922 39622 75978
rect 39678 75922 57250 75978
rect 57306 75922 57374 75978
rect 57430 75922 57498 75978
rect 57554 75922 57622 75978
rect 57678 75922 64518 75978
rect 64574 75922 64642 75978
rect 64698 75922 66564 75978
rect -1916 75826 66564 75922
rect 239468 76412 350740 76446
rect 239468 76356 284022 76412
rect 284078 76356 284146 76412
rect 284202 76356 284270 76412
rect 284326 76356 284394 76412
rect 284450 76356 284518 76412
rect 284574 76356 284642 76412
rect 284698 76356 284766 76412
rect 284822 76356 284890 76412
rect 284946 76356 285014 76412
rect 285070 76356 285138 76412
rect 285194 76356 304022 76412
rect 304078 76356 304146 76412
rect 304202 76356 304270 76412
rect 304326 76356 304394 76412
rect 304450 76356 304518 76412
rect 304574 76356 304642 76412
rect 304698 76356 304766 76412
rect 304822 76356 304890 76412
rect 304946 76356 305014 76412
rect 305070 76356 305138 76412
rect 305194 76356 350740 76412
rect 239468 76350 350740 76356
rect 239468 76294 255250 76350
rect 255306 76294 255374 76350
rect 255430 76294 255498 76350
rect 255554 76294 255622 76350
rect 255678 76294 273250 76350
rect 273306 76294 273374 76350
rect 273430 76294 273498 76350
rect 273554 76294 273622 76350
rect 273678 76294 291250 76350
rect 291306 76294 291374 76350
rect 291430 76294 291498 76350
rect 291554 76294 291622 76350
rect 291678 76294 309250 76350
rect 309306 76294 309374 76350
rect 309430 76294 309498 76350
rect 309554 76294 309622 76350
rect 309678 76294 327250 76350
rect 327306 76294 327374 76350
rect 327430 76294 327498 76350
rect 327554 76294 327622 76350
rect 327678 76294 345250 76350
rect 345306 76294 345374 76350
rect 345430 76294 345498 76350
rect 345554 76294 345622 76350
rect 345678 76294 350740 76350
rect 239468 76288 350740 76294
rect 239468 76232 284022 76288
rect 284078 76232 284146 76288
rect 284202 76232 284270 76288
rect 284326 76232 284394 76288
rect 284450 76232 284518 76288
rect 284574 76232 284642 76288
rect 284698 76232 284766 76288
rect 284822 76232 284890 76288
rect 284946 76232 285014 76288
rect 285070 76232 285138 76288
rect 285194 76232 304022 76288
rect 304078 76232 304146 76288
rect 304202 76232 304270 76288
rect 304326 76232 304394 76288
rect 304450 76232 304518 76288
rect 304574 76232 304642 76288
rect 304698 76232 304766 76288
rect 304822 76232 304890 76288
rect 304946 76232 305014 76288
rect 305070 76232 305138 76288
rect 305194 76232 350740 76288
rect 239468 76226 350740 76232
rect 239468 76170 255250 76226
rect 255306 76170 255374 76226
rect 255430 76170 255498 76226
rect 255554 76170 255622 76226
rect 255678 76170 273250 76226
rect 273306 76170 273374 76226
rect 273430 76170 273498 76226
rect 273554 76170 273622 76226
rect 273678 76170 291250 76226
rect 291306 76170 291374 76226
rect 291430 76170 291498 76226
rect 291554 76170 291622 76226
rect 291678 76170 309250 76226
rect 309306 76170 309374 76226
rect 309430 76170 309498 76226
rect 309554 76170 309622 76226
rect 309678 76170 327250 76226
rect 327306 76170 327374 76226
rect 327430 76170 327498 76226
rect 327554 76170 327622 76226
rect 327678 76170 345250 76226
rect 345306 76170 345374 76226
rect 345430 76170 345498 76226
rect 345554 76170 345622 76226
rect 345678 76170 350740 76226
rect 239468 76164 350740 76170
rect 239468 76108 284022 76164
rect 284078 76108 284146 76164
rect 284202 76108 284270 76164
rect 284326 76108 284394 76164
rect 284450 76108 284518 76164
rect 284574 76108 284642 76164
rect 284698 76108 284766 76164
rect 284822 76108 284890 76164
rect 284946 76108 285014 76164
rect 285070 76108 285138 76164
rect 285194 76108 304022 76164
rect 304078 76108 304146 76164
rect 304202 76108 304270 76164
rect 304326 76108 304394 76164
rect 304450 76108 304518 76164
rect 304574 76108 304642 76164
rect 304698 76108 304766 76164
rect 304822 76108 304890 76164
rect 304946 76108 305014 76164
rect 305070 76108 305138 76164
rect 305194 76108 350740 76164
rect 239468 76102 350740 76108
rect 239468 76046 255250 76102
rect 255306 76046 255374 76102
rect 255430 76046 255498 76102
rect 255554 76046 255622 76102
rect 255678 76046 273250 76102
rect 273306 76046 273374 76102
rect 273430 76046 273498 76102
rect 273554 76046 273622 76102
rect 273678 76046 291250 76102
rect 291306 76046 291374 76102
rect 291430 76046 291498 76102
rect 291554 76046 291622 76102
rect 291678 76046 309250 76102
rect 309306 76046 309374 76102
rect 309430 76046 309498 76102
rect 309554 76046 309622 76102
rect 309678 76046 327250 76102
rect 327306 76046 327374 76102
rect 327430 76046 327498 76102
rect 327554 76046 327622 76102
rect 327678 76046 345250 76102
rect 345306 76046 345374 76102
rect 345430 76046 345498 76102
rect 345554 76046 345622 76102
rect 345678 76046 350740 76102
rect 239468 76040 350740 76046
rect 239468 75984 284022 76040
rect 284078 75984 284146 76040
rect 284202 75984 284270 76040
rect 284326 75984 284394 76040
rect 284450 75984 284518 76040
rect 284574 75984 284642 76040
rect 284698 75984 284766 76040
rect 284822 75984 284890 76040
rect 284946 75984 285014 76040
rect 285070 75984 285138 76040
rect 285194 75984 304022 76040
rect 304078 75984 304146 76040
rect 304202 75984 304270 76040
rect 304326 75984 304394 76040
rect 304450 75984 304518 76040
rect 304574 75984 304642 76040
rect 304698 75984 304766 76040
rect 304822 75984 304890 76040
rect 304946 75984 305014 76040
rect 305070 75984 305138 76040
rect 305194 75984 350740 76040
rect 239468 75978 350740 75984
rect 239468 75922 255250 75978
rect 255306 75922 255374 75978
rect 255430 75922 255498 75978
rect 255554 75922 255622 75978
rect 255678 75922 273250 75978
rect 273306 75922 273374 75978
rect 273430 75922 273498 75978
rect 273554 75922 273622 75978
rect 273678 75922 291250 75978
rect 291306 75922 291374 75978
rect 291430 75922 291498 75978
rect 291554 75922 291622 75978
rect 291678 75922 309250 75978
rect 309306 75922 309374 75978
rect 309430 75922 309498 75978
rect 309554 75922 309622 75978
rect 309678 75922 327250 75978
rect 327306 75922 327374 75978
rect 327430 75922 327498 75978
rect 327554 75922 327622 75978
rect 327678 75922 345250 75978
rect 345306 75922 345374 75978
rect 345430 75922 345498 75978
rect 345554 75922 345622 75978
rect 345678 75922 350740 75978
rect 239468 75916 350740 75922
rect 239468 75860 284022 75916
rect 284078 75860 284146 75916
rect 284202 75860 284270 75916
rect 284326 75860 284394 75916
rect 284450 75860 284518 75916
rect 284574 75860 284642 75916
rect 284698 75860 284766 75916
rect 284822 75860 284890 75916
rect 284946 75860 285014 75916
rect 285070 75860 285138 75916
rect 285194 75860 304022 75916
rect 304078 75860 304146 75916
rect 304202 75860 304270 75916
rect 304326 75860 304394 75916
rect 304450 75860 304518 75916
rect 304574 75860 304642 75916
rect 304698 75860 304766 75916
rect 304822 75860 304890 75916
rect 304946 75860 305014 75916
rect 305070 75860 305138 75916
rect 305194 75860 350740 75916
rect 239468 75826 350740 75860
rect 545484 76350 597980 76446
rect 545484 76294 561250 76350
rect 561306 76294 561374 76350
rect 561430 76294 561498 76350
rect 561554 76294 561622 76350
rect 561678 76294 579250 76350
rect 579306 76294 579374 76350
rect 579430 76294 579498 76350
rect 579554 76294 579622 76350
rect 579678 76294 596496 76350
rect 596552 76294 596620 76350
rect 596676 76294 596744 76350
rect 596800 76294 596868 76350
rect 596924 76294 597980 76350
rect 545484 76226 597980 76294
rect 545484 76170 561250 76226
rect 561306 76170 561374 76226
rect 561430 76170 561498 76226
rect 561554 76170 561622 76226
rect 561678 76170 579250 76226
rect 579306 76170 579374 76226
rect 579430 76170 579498 76226
rect 579554 76170 579622 76226
rect 579678 76170 596496 76226
rect 596552 76170 596620 76226
rect 596676 76170 596744 76226
rect 596800 76170 596868 76226
rect 596924 76170 597980 76226
rect 545484 76102 597980 76170
rect 545484 76046 561250 76102
rect 561306 76046 561374 76102
rect 561430 76046 561498 76102
rect 561554 76046 561622 76102
rect 561678 76046 579250 76102
rect 579306 76046 579374 76102
rect 579430 76046 579498 76102
rect 579554 76046 579622 76102
rect 579678 76046 596496 76102
rect 596552 76046 596620 76102
rect 596676 76046 596744 76102
rect 596800 76046 596868 76102
rect 596924 76046 597980 76102
rect 545484 75978 597980 76046
rect 545484 75922 561250 75978
rect 561306 75922 561374 75978
rect 561430 75922 561498 75978
rect 561554 75922 561622 75978
rect 561678 75922 579250 75978
rect 579306 75922 579374 75978
rect 579430 75922 579498 75978
rect 579554 75922 579622 75978
rect 579678 75922 596496 75978
rect 596552 75922 596620 75978
rect 596676 75922 596744 75978
rect 596800 75922 596868 75978
rect 596924 75922 597980 75978
rect 545484 75826 597980 75922
rect -1916 64350 66564 64446
rect -1916 64294 -1820 64350
rect -1764 64294 -1696 64350
rect -1640 64294 -1572 64350
rect -1516 64294 -1448 64350
rect -1392 64294 6970 64350
rect 7026 64294 7094 64350
rect 7150 64294 7218 64350
rect 7274 64294 7342 64350
rect 7398 64294 24970 64350
rect 25026 64294 25094 64350
rect 25150 64294 25218 64350
rect 25274 64294 25342 64350
rect 25398 64294 42970 64350
rect 43026 64294 43094 64350
rect 43150 64294 43218 64350
rect 43274 64294 43342 64350
rect 43398 64294 66564 64350
rect -1916 64226 66564 64294
rect -1916 64170 -1820 64226
rect -1764 64170 -1696 64226
rect -1640 64170 -1572 64226
rect -1516 64170 -1448 64226
rect -1392 64170 6970 64226
rect 7026 64170 7094 64226
rect 7150 64170 7218 64226
rect 7274 64170 7342 64226
rect 7398 64170 24970 64226
rect 25026 64170 25094 64226
rect 25150 64170 25218 64226
rect 25274 64170 25342 64226
rect 25398 64170 42970 64226
rect 43026 64170 43094 64226
rect 43150 64170 43218 64226
rect 43274 64170 43342 64226
rect 43398 64170 66564 64226
rect -1916 64102 66564 64170
rect -1916 64046 -1820 64102
rect -1764 64046 -1696 64102
rect -1640 64046 -1572 64102
rect -1516 64046 -1448 64102
rect -1392 64046 6970 64102
rect 7026 64046 7094 64102
rect 7150 64046 7218 64102
rect 7274 64046 7342 64102
rect 7398 64046 24970 64102
rect 25026 64046 25094 64102
rect 25150 64046 25218 64102
rect 25274 64046 25342 64102
rect 25398 64046 42970 64102
rect 43026 64046 43094 64102
rect 43150 64046 43218 64102
rect 43274 64046 43342 64102
rect 43398 64046 66564 64102
rect -1916 63978 66564 64046
rect -1916 63922 -1820 63978
rect -1764 63922 -1696 63978
rect -1640 63922 -1572 63978
rect -1516 63922 -1448 63978
rect -1392 63922 6970 63978
rect 7026 63922 7094 63978
rect 7150 63922 7218 63978
rect 7274 63922 7342 63978
rect 7398 63922 24970 63978
rect 25026 63922 25094 63978
rect 25150 63922 25218 63978
rect 25274 63922 25342 63978
rect 25398 63922 42970 63978
rect 43026 63922 43094 63978
rect 43150 63922 43218 63978
rect 43274 63922 43342 63978
rect 43398 63922 66564 63978
rect -1916 63826 66564 63922
rect 239468 64350 350740 64446
rect 239468 64294 240970 64350
rect 241026 64294 241094 64350
rect 241150 64294 241218 64350
rect 241274 64294 241342 64350
rect 241398 64294 258970 64350
rect 259026 64294 259094 64350
rect 259150 64294 259218 64350
rect 259274 64294 259342 64350
rect 259398 64294 276970 64350
rect 277026 64294 277094 64350
rect 277150 64294 277218 64350
rect 277274 64294 277342 64350
rect 277398 64294 294970 64350
rect 295026 64294 295094 64350
rect 295150 64294 295218 64350
rect 295274 64294 295342 64350
rect 295398 64294 312970 64350
rect 313026 64294 313094 64350
rect 313150 64294 313218 64350
rect 313274 64294 313342 64350
rect 313398 64294 330970 64350
rect 331026 64294 331094 64350
rect 331150 64294 331218 64350
rect 331274 64294 331342 64350
rect 331398 64294 348970 64350
rect 349026 64294 349094 64350
rect 349150 64294 349218 64350
rect 349274 64294 349342 64350
rect 349398 64294 350740 64350
rect 239468 64226 350740 64294
rect 239468 64170 240970 64226
rect 241026 64170 241094 64226
rect 241150 64170 241218 64226
rect 241274 64170 241342 64226
rect 241398 64170 258970 64226
rect 259026 64170 259094 64226
rect 259150 64170 259218 64226
rect 259274 64170 259342 64226
rect 259398 64170 276970 64226
rect 277026 64170 277094 64226
rect 277150 64170 277218 64226
rect 277274 64170 277342 64226
rect 277398 64170 294970 64226
rect 295026 64170 295094 64226
rect 295150 64170 295218 64226
rect 295274 64170 295342 64226
rect 295398 64170 312970 64226
rect 313026 64170 313094 64226
rect 313150 64170 313218 64226
rect 313274 64170 313342 64226
rect 313398 64170 330970 64226
rect 331026 64170 331094 64226
rect 331150 64170 331218 64226
rect 331274 64170 331342 64226
rect 331398 64170 348970 64226
rect 349026 64170 349094 64226
rect 349150 64170 349218 64226
rect 349274 64170 349342 64226
rect 349398 64170 350740 64226
rect 239468 64102 350740 64170
rect 239468 64046 240970 64102
rect 241026 64046 241094 64102
rect 241150 64046 241218 64102
rect 241274 64046 241342 64102
rect 241398 64046 258970 64102
rect 259026 64046 259094 64102
rect 259150 64046 259218 64102
rect 259274 64046 259342 64102
rect 259398 64046 276970 64102
rect 277026 64046 277094 64102
rect 277150 64046 277218 64102
rect 277274 64046 277342 64102
rect 277398 64046 294970 64102
rect 295026 64046 295094 64102
rect 295150 64046 295218 64102
rect 295274 64046 295342 64102
rect 295398 64046 312970 64102
rect 313026 64046 313094 64102
rect 313150 64046 313218 64102
rect 313274 64046 313342 64102
rect 313398 64046 330970 64102
rect 331026 64046 331094 64102
rect 331150 64046 331218 64102
rect 331274 64046 331342 64102
rect 331398 64046 348970 64102
rect 349026 64046 349094 64102
rect 349150 64046 349218 64102
rect 349274 64046 349342 64102
rect 349398 64046 350740 64102
rect 239468 63978 350740 64046
rect 239468 63922 240970 63978
rect 241026 63922 241094 63978
rect 241150 63922 241218 63978
rect 241274 63922 241342 63978
rect 241398 63922 258970 63978
rect 259026 63922 259094 63978
rect 259150 63922 259218 63978
rect 259274 63922 259342 63978
rect 259398 63922 276970 63978
rect 277026 63922 277094 63978
rect 277150 63922 277218 63978
rect 277274 63922 277342 63978
rect 277398 63922 294970 63978
rect 295026 63922 295094 63978
rect 295150 63922 295218 63978
rect 295274 63922 295342 63978
rect 295398 63922 312970 63978
rect 313026 63922 313094 63978
rect 313150 63922 313218 63978
rect 313274 63922 313342 63978
rect 313398 63922 330970 63978
rect 331026 63922 331094 63978
rect 331150 63922 331218 63978
rect 331274 63922 331342 63978
rect 331398 63922 348970 63978
rect 349026 63922 349094 63978
rect 349150 63922 349218 63978
rect 349274 63922 349342 63978
rect 349398 63922 350740 63978
rect 239468 63826 350740 63922
rect 545484 64350 597980 64446
rect 545484 64294 564970 64350
rect 565026 64294 565094 64350
rect 565150 64294 565218 64350
rect 565274 64294 565342 64350
rect 565398 64294 582970 64350
rect 583026 64294 583094 64350
rect 583150 64294 583218 64350
rect 583274 64294 583342 64350
rect 583398 64294 597456 64350
rect 597512 64294 597580 64350
rect 597636 64294 597704 64350
rect 597760 64294 597828 64350
rect 597884 64294 597980 64350
rect 545484 64226 597980 64294
rect 545484 64170 564970 64226
rect 565026 64170 565094 64226
rect 565150 64170 565218 64226
rect 565274 64170 565342 64226
rect 565398 64170 582970 64226
rect 583026 64170 583094 64226
rect 583150 64170 583218 64226
rect 583274 64170 583342 64226
rect 583398 64170 597456 64226
rect 597512 64170 597580 64226
rect 597636 64170 597704 64226
rect 597760 64170 597828 64226
rect 597884 64170 597980 64226
rect 545484 64102 597980 64170
rect 545484 64046 564970 64102
rect 565026 64046 565094 64102
rect 565150 64046 565218 64102
rect 565274 64046 565342 64102
rect 565398 64046 582970 64102
rect 583026 64046 583094 64102
rect 583150 64046 583218 64102
rect 583274 64046 583342 64102
rect 583398 64046 597456 64102
rect 597512 64046 597580 64102
rect 597636 64046 597704 64102
rect 597760 64046 597828 64102
rect 597884 64046 597980 64102
rect 545484 63978 597980 64046
rect 545484 63922 564970 63978
rect 565026 63922 565094 63978
rect 565150 63922 565218 63978
rect 565274 63922 565342 63978
rect 565398 63922 582970 63978
rect 583026 63922 583094 63978
rect 583150 63922 583218 63978
rect 583274 63922 583342 63978
rect 583398 63922 597456 63978
rect 597512 63922 597580 63978
rect 597636 63922 597704 63978
rect 597760 63922 597828 63978
rect 597884 63922 597980 63978
rect 545484 63826 597980 63922
rect 548924 59878 550132 59894
rect 548924 59822 548940 59878
rect 548996 59822 550060 59878
rect 550116 59822 550132 59878
rect 548924 59806 550132 59822
rect -1916 58350 66564 58446
rect -1916 58294 -860 58350
rect -804 58294 -736 58350
rect -680 58294 -612 58350
rect -556 58294 -488 58350
rect -432 58294 3250 58350
rect 3306 58294 3374 58350
rect 3430 58294 3498 58350
rect 3554 58294 3622 58350
rect 3678 58294 21250 58350
rect 21306 58294 21374 58350
rect 21430 58294 21498 58350
rect 21554 58294 21622 58350
rect 21678 58294 39250 58350
rect 39306 58294 39374 58350
rect 39430 58294 39498 58350
rect 39554 58294 39622 58350
rect 39678 58294 57250 58350
rect 57306 58294 57374 58350
rect 57430 58294 57498 58350
rect 57554 58294 57622 58350
rect 57678 58294 64518 58350
rect 64574 58294 64642 58350
rect 64698 58294 66564 58350
rect -1916 58226 66564 58294
rect -1916 58170 -860 58226
rect -804 58170 -736 58226
rect -680 58170 -612 58226
rect -556 58170 -488 58226
rect -432 58170 3250 58226
rect 3306 58170 3374 58226
rect 3430 58170 3498 58226
rect 3554 58170 3622 58226
rect 3678 58170 21250 58226
rect 21306 58170 21374 58226
rect 21430 58170 21498 58226
rect 21554 58170 21622 58226
rect 21678 58170 39250 58226
rect 39306 58170 39374 58226
rect 39430 58170 39498 58226
rect 39554 58170 39622 58226
rect 39678 58170 57250 58226
rect 57306 58170 57374 58226
rect 57430 58170 57498 58226
rect 57554 58170 57622 58226
rect 57678 58170 64518 58226
rect 64574 58170 64642 58226
rect 64698 58170 66564 58226
rect -1916 58102 66564 58170
rect -1916 58046 -860 58102
rect -804 58046 -736 58102
rect -680 58046 -612 58102
rect -556 58046 -488 58102
rect -432 58046 3250 58102
rect 3306 58046 3374 58102
rect 3430 58046 3498 58102
rect 3554 58046 3622 58102
rect 3678 58046 21250 58102
rect 21306 58046 21374 58102
rect 21430 58046 21498 58102
rect 21554 58046 21622 58102
rect 21678 58046 39250 58102
rect 39306 58046 39374 58102
rect 39430 58046 39498 58102
rect 39554 58046 39622 58102
rect 39678 58046 57250 58102
rect 57306 58046 57374 58102
rect 57430 58046 57498 58102
rect 57554 58046 57622 58102
rect 57678 58046 64518 58102
rect 64574 58046 64642 58102
rect 64698 58046 66564 58102
rect -1916 57978 66564 58046
rect -1916 57922 -860 57978
rect -804 57922 -736 57978
rect -680 57922 -612 57978
rect -556 57922 -488 57978
rect -432 57922 3250 57978
rect 3306 57922 3374 57978
rect 3430 57922 3498 57978
rect 3554 57922 3622 57978
rect 3678 57922 21250 57978
rect 21306 57922 21374 57978
rect 21430 57922 21498 57978
rect 21554 57922 21622 57978
rect 21678 57922 39250 57978
rect 39306 57922 39374 57978
rect 39430 57922 39498 57978
rect 39554 57922 39622 57978
rect 39678 57922 57250 57978
rect 57306 57922 57374 57978
rect 57430 57922 57498 57978
rect 57554 57922 57622 57978
rect 57678 57922 64518 57978
rect 64574 57922 64642 57978
rect 64698 57922 66564 57978
rect -1916 57826 66564 57922
rect 239468 58350 350740 58446
rect 239468 58294 255250 58350
rect 255306 58294 255374 58350
rect 255430 58294 255498 58350
rect 255554 58294 255622 58350
rect 255678 58294 273250 58350
rect 273306 58294 273374 58350
rect 273430 58294 273498 58350
rect 273554 58294 273622 58350
rect 273678 58294 291250 58350
rect 291306 58294 291374 58350
rect 291430 58294 291498 58350
rect 291554 58294 291622 58350
rect 291678 58294 309250 58350
rect 309306 58294 309374 58350
rect 309430 58294 309498 58350
rect 309554 58294 309622 58350
rect 309678 58294 327250 58350
rect 327306 58294 327374 58350
rect 327430 58294 327498 58350
rect 327554 58294 327622 58350
rect 327678 58294 345250 58350
rect 345306 58294 345374 58350
rect 345430 58294 345498 58350
rect 345554 58294 345622 58350
rect 345678 58294 350740 58350
rect 239468 58226 350740 58294
rect 239468 58170 255250 58226
rect 255306 58170 255374 58226
rect 255430 58170 255498 58226
rect 255554 58170 255622 58226
rect 255678 58170 273250 58226
rect 273306 58170 273374 58226
rect 273430 58170 273498 58226
rect 273554 58170 273622 58226
rect 273678 58170 291250 58226
rect 291306 58170 291374 58226
rect 291430 58170 291498 58226
rect 291554 58170 291622 58226
rect 291678 58170 309250 58226
rect 309306 58170 309374 58226
rect 309430 58170 309498 58226
rect 309554 58170 309622 58226
rect 309678 58170 327250 58226
rect 327306 58170 327374 58226
rect 327430 58170 327498 58226
rect 327554 58170 327622 58226
rect 327678 58170 345250 58226
rect 345306 58170 345374 58226
rect 345430 58170 345498 58226
rect 345554 58170 345622 58226
rect 345678 58170 350740 58226
rect 239468 58102 350740 58170
rect 239468 58046 255250 58102
rect 255306 58046 255374 58102
rect 255430 58046 255498 58102
rect 255554 58046 255622 58102
rect 255678 58046 273250 58102
rect 273306 58046 273374 58102
rect 273430 58046 273498 58102
rect 273554 58046 273622 58102
rect 273678 58046 291250 58102
rect 291306 58046 291374 58102
rect 291430 58046 291498 58102
rect 291554 58046 291622 58102
rect 291678 58046 309250 58102
rect 309306 58046 309374 58102
rect 309430 58046 309498 58102
rect 309554 58046 309622 58102
rect 309678 58046 327250 58102
rect 327306 58046 327374 58102
rect 327430 58046 327498 58102
rect 327554 58046 327622 58102
rect 327678 58046 345250 58102
rect 345306 58046 345374 58102
rect 345430 58046 345498 58102
rect 345554 58046 345622 58102
rect 345678 58046 350740 58102
rect 239468 57978 350740 58046
rect 239468 57922 255250 57978
rect 255306 57922 255374 57978
rect 255430 57922 255498 57978
rect 255554 57922 255622 57978
rect 255678 57922 273250 57978
rect 273306 57922 273374 57978
rect 273430 57922 273498 57978
rect 273554 57922 273622 57978
rect 273678 57922 291250 57978
rect 291306 57922 291374 57978
rect 291430 57922 291498 57978
rect 291554 57922 291622 57978
rect 291678 57922 309250 57978
rect 309306 57922 309374 57978
rect 309430 57922 309498 57978
rect 309554 57922 309622 57978
rect 309678 57922 327250 57978
rect 327306 57922 327374 57978
rect 327430 57922 327498 57978
rect 327554 57922 327622 57978
rect 327678 57922 345250 57978
rect 345306 57922 345374 57978
rect 345430 57922 345498 57978
rect 345554 57922 345622 57978
rect 345678 57922 350740 57978
rect 239468 57826 350740 57922
rect 545484 58350 597980 58446
rect 545484 58294 561250 58350
rect 561306 58294 561374 58350
rect 561430 58294 561498 58350
rect 561554 58294 561622 58350
rect 561678 58294 596496 58350
rect 596552 58294 596620 58350
rect 596676 58294 596744 58350
rect 596800 58294 596868 58350
rect 596924 58294 597980 58350
rect 545484 58226 597980 58294
rect 545484 58170 561250 58226
rect 561306 58170 561374 58226
rect 561430 58170 561498 58226
rect 561554 58170 561622 58226
rect 561678 58170 596496 58226
rect 596552 58170 596620 58226
rect 596676 58170 596744 58226
rect 596800 58170 596868 58226
rect 596924 58170 597980 58226
rect 545484 58102 597980 58170
rect 545484 58046 561250 58102
rect 561306 58046 561374 58102
rect 561430 58046 561498 58102
rect 561554 58046 561622 58102
rect 561678 58046 596496 58102
rect 596552 58046 596620 58102
rect 596676 58046 596744 58102
rect 596800 58046 596868 58102
rect 596924 58046 597980 58102
rect 545484 57978 597980 58046
rect 545484 57922 561250 57978
rect 561306 57922 561374 57978
rect 561430 57922 561498 57978
rect 561554 57922 561622 57978
rect 561678 57922 596496 57978
rect 596552 57922 596620 57978
rect 596676 57922 596744 57978
rect 596800 57922 596868 57978
rect 596924 57922 597980 57978
rect 545484 57826 597980 57922
rect 548700 54658 549460 54674
rect 548700 54602 548716 54658
rect 548772 54602 549388 54658
rect 549444 54602 549460 54658
rect 548700 54586 549460 54602
rect 548700 51598 549460 51614
rect 548700 51542 548716 51598
rect 548772 51542 549388 51598
rect 549444 51542 549460 51598
rect 548700 51526 549460 51542
rect 548588 49798 549460 49814
rect 548588 49742 548604 49798
rect 548660 49742 549388 49798
rect 549444 49742 549460 49798
rect 548588 49726 549460 49742
rect 557324 47818 584964 47834
rect 557324 47762 557340 47818
rect 557396 47762 584892 47818
rect 584948 47762 584964 47818
rect 557324 47746 584964 47762
rect -1916 46350 66564 46446
rect -1916 46294 -1820 46350
rect -1764 46294 -1696 46350
rect -1640 46294 -1572 46350
rect -1516 46294 -1448 46350
rect -1392 46294 6970 46350
rect 7026 46294 7094 46350
rect 7150 46294 7218 46350
rect 7274 46294 7342 46350
rect 7398 46294 24970 46350
rect 25026 46294 25094 46350
rect 25150 46294 25218 46350
rect 25274 46294 25342 46350
rect 25398 46294 42970 46350
rect 43026 46294 43094 46350
rect 43150 46294 43218 46350
rect 43274 46294 43342 46350
rect 43398 46294 66564 46350
rect -1916 46226 66564 46294
rect -1916 46170 -1820 46226
rect -1764 46170 -1696 46226
rect -1640 46170 -1572 46226
rect -1516 46170 -1448 46226
rect -1392 46170 6970 46226
rect 7026 46170 7094 46226
rect 7150 46170 7218 46226
rect 7274 46170 7342 46226
rect 7398 46170 24970 46226
rect 25026 46170 25094 46226
rect 25150 46170 25218 46226
rect 25274 46170 25342 46226
rect 25398 46170 42970 46226
rect 43026 46170 43094 46226
rect 43150 46170 43218 46226
rect 43274 46170 43342 46226
rect 43398 46170 66564 46226
rect -1916 46102 66564 46170
rect -1916 46046 -1820 46102
rect -1764 46046 -1696 46102
rect -1640 46046 -1572 46102
rect -1516 46046 -1448 46102
rect -1392 46046 6970 46102
rect 7026 46046 7094 46102
rect 7150 46046 7218 46102
rect 7274 46046 7342 46102
rect 7398 46046 24970 46102
rect 25026 46046 25094 46102
rect 25150 46046 25218 46102
rect 25274 46046 25342 46102
rect 25398 46046 42970 46102
rect 43026 46046 43094 46102
rect 43150 46046 43218 46102
rect 43274 46046 43342 46102
rect 43398 46046 66564 46102
rect -1916 45978 66564 46046
rect -1916 45922 -1820 45978
rect -1764 45922 -1696 45978
rect -1640 45922 -1572 45978
rect -1516 45922 -1448 45978
rect -1392 45922 6970 45978
rect 7026 45922 7094 45978
rect 7150 45922 7218 45978
rect 7274 45922 7342 45978
rect 7398 45922 24970 45978
rect 25026 45922 25094 45978
rect 25150 45922 25218 45978
rect 25274 45922 25342 45978
rect 25398 45922 42970 45978
rect 43026 45922 43094 45978
rect 43150 45922 43218 45978
rect 43274 45922 43342 45978
rect 43398 45922 66564 45978
rect -1916 45826 66564 45922
rect 239468 46350 350740 46446
rect 239468 46294 240970 46350
rect 241026 46294 241094 46350
rect 241150 46294 241218 46350
rect 241274 46294 241342 46350
rect 241398 46294 258970 46350
rect 259026 46294 259094 46350
rect 259150 46294 259218 46350
rect 259274 46294 259342 46350
rect 259398 46294 276970 46350
rect 277026 46294 277094 46350
rect 277150 46294 277218 46350
rect 277274 46294 277342 46350
rect 277398 46294 294970 46350
rect 295026 46294 295094 46350
rect 295150 46294 295218 46350
rect 295274 46294 295342 46350
rect 295398 46294 312970 46350
rect 313026 46294 313094 46350
rect 313150 46294 313218 46350
rect 313274 46294 313342 46350
rect 313398 46294 330970 46350
rect 331026 46294 331094 46350
rect 331150 46294 331218 46350
rect 331274 46294 331342 46350
rect 331398 46294 348970 46350
rect 349026 46294 349094 46350
rect 349150 46294 349218 46350
rect 349274 46294 349342 46350
rect 349398 46294 350740 46350
rect 239468 46226 350740 46294
rect 239468 46170 240970 46226
rect 241026 46170 241094 46226
rect 241150 46170 241218 46226
rect 241274 46170 241342 46226
rect 241398 46170 258970 46226
rect 259026 46170 259094 46226
rect 259150 46170 259218 46226
rect 259274 46170 259342 46226
rect 259398 46170 276970 46226
rect 277026 46170 277094 46226
rect 277150 46170 277218 46226
rect 277274 46170 277342 46226
rect 277398 46170 294970 46226
rect 295026 46170 295094 46226
rect 295150 46170 295218 46226
rect 295274 46170 295342 46226
rect 295398 46170 312970 46226
rect 313026 46170 313094 46226
rect 313150 46170 313218 46226
rect 313274 46170 313342 46226
rect 313398 46170 330970 46226
rect 331026 46170 331094 46226
rect 331150 46170 331218 46226
rect 331274 46170 331342 46226
rect 331398 46170 348970 46226
rect 349026 46170 349094 46226
rect 349150 46170 349218 46226
rect 349274 46170 349342 46226
rect 349398 46170 350740 46226
rect 239468 46102 350740 46170
rect 239468 46046 240970 46102
rect 241026 46046 241094 46102
rect 241150 46046 241218 46102
rect 241274 46046 241342 46102
rect 241398 46046 258970 46102
rect 259026 46046 259094 46102
rect 259150 46046 259218 46102
rect 259274 46046 259342 46102
rect 259398 46046 276970 46102
rect 277026 46046 277094 46102
rect 277150 46046 277218 46102
rect 277274 46046 277342 46102
rect 277398 46046 294970 46102
rect 295026 46046 295094 46102
rect 295150 46046 295218 46102
rect 295274 46046 295342 46102
rect 295398 46046 312970 46102
rect 313026 46046 313094 46102
rect 313150 46046 313218 46102
rect 313274 46046 313342 46102
rect 313398 46046 330970 46102
rect 331026 46046 331094 46102
rect 331150 46046 331218 46102
rect 331274 46046 331342 46102
rect 331398 46046 348970 46102
rect 349026 46046 349094 46102
rect 349150 46046 349218 46102
rect 349274 46046 349342 46102
rect 349398 46046 350740 46102
rect 239468 45978 350740 46046
rect 239468 45922 240970 45978
rect 241026 45922 241094 45978
rect 241150 45922 241218 45978
rect 241274 45922 241342 45978
rect 241398 45922 258970 45978
rect 259026 45922 259094 45978
rect 259150 45922 259218 45978
rect 259274 45922 259342 45978
rect 259398 45922 276970 45978
rect 277026 45922 277094 45978
rect 277150 45922 277218 45978
rect 277274 45922 277342 45978
rect 277398 45922 294970 45978
rect 295026 45922 295094 45978
rect 295150 45922 295218 45978
rect 295274 45922 295342 45978
rect 295398 45922 312970 45978
rect 313026 45922 313094 45978
rect 313150 45922 313218 45978
rect 313274 45922 313342 45978
rect 313398 45922 330970 45978
rect 331026 45922 331094 45978
rect 331150 45922 331218 45978
rect 331274 45922 331342 45978
rect 331398 45922 348970 45978
rect 349026 45922 349094 45978
rect 349150 45922 349218 45978
rect 349274 45922 349342 45978
rect 349398 45922 350740 45978
rect 239468 45826 350740 45922
rect 545484 46412 597980 46446
rect 545484 46356 568022 46412
rect 568078 46356 568146 46412
rect 568202 46356 568270 46412
rect 568326 46356 568394 46412
rect 568450 46356 568518 46412
rect 568574 46356 568642 46412
rect 568698 46356 568766 46412
rect 568822 46356 568890 46412
rect 568946 46356 569014 46412
rect 569070 46356 569138 46412
rect 569194 46356 588022 46412
rect 588078 46356 588146 46412
rect 588202 46356 588270 46412
rect 588326 46356 588394 46412
rect 588450 46356 588518 46412
rect 588574 46356 588642 46412
rect 588698 46356 588766 46412
rect 588822 46356 588890 46412
rect 588946 46356 589014 46412
rect 589070 46356 589138 46412
rect 589194 46356 597980 46412
rect 545484 46350 597980 46356
rect 545484 46294 564970 46350
rect 565026 46294 565094 46350
rect 565150 46294 565218 46350
rect 565274 46294 565342 46350
rect 565398 46294 582970 46350
rect 583026 46294 583094 46350
rect 583150 46294 583218 46350
rect 583274 46294 583342 46350
rect 583398 46294 597456 46350
rect 597512 46294 597580 46350
rect 597636 46294 597704 46350
rect 597760 46294 597828 46350
rect 597884 46294 597980 46350
rect 545484 46288 597980 46294
rect 545484 46232 568022 46288
rect 568078 46232 568146 46288
rect 568202 46232 568270 46288
rect 568326 46232 568394 46288
rect 568450 46232 568518 46288
rect 568574 46232 568642 46288
rect 568698 46232 568766 46288
rect 568822 46232 568890 46288
rect 568946 46232 569014 46288
rect 569070 46232 569138 46288
rect 569194 46232 588022 46288
rect 588078 46232 588146 46288
rect 588202 46232 588270 46288
rect 588326 46232 588394 46288
rect 588450 46232 588518 46288
rect 588574 46232 588642 46288
rect 588698 46232 588766 46288
rect 588822 46232 588890 46288
rect 588946 46232 589014 46288
rect 589070 46232 589138 46288
rect 589194 46232 597980 46288
rect 545484 46226 597980 46232
rect 545484 46170 564970 46226
rect 565026 46170 565094 46226
rect 565150 46170 565218 46226
rect 565274 46170 565342 46226
rect 565398 46170 582970 46226
rect 583026 46170 583094 46226
rect 583150 46170 583218 46226
rect 583274 46170 583342 46226
rect 583398 46170 597456 46226
rect 597512 46170 597580 46226
rect 597636 46170 597704 46226
rect 597760 46170 597828 46226
rect 597884 46170 597980 46226
rect 545484 46164 597980 46170
rect 545484 46108 568022 46164
rect 568078 46108 568146 46164
rect 568202 46108 568270 46164
rect 568326 46108 568394 46164
rect 568450 46108 568518 46164
rect 568574 46108 568642 46164
rect 568698 46108 568766 46164
rect 568822 46108 568890 46164
rect 568946 46108 569014 46164
rect 569070 46108 569138 46164
rect 569194 46108 588022 46164
rect 588078 46108 588146 46164
rect 588202 46108 588270 46164
rect 588326 46108 588394 46164
rect 588450 46108 588518 46164
rect 588574 46108 588642 46164
rect 588698 46108 588766 46164
rect 588822 46108 588890 46164
rect 588946 46108 589014 46164
rect 589070 46108 589138 46164
rect 589194 46108 597980 46164
rect 545484 46102 597980 46108
rect 545484 46046 564970 46102
rect 565026 46046 565094 46102
rect 565150 46046 565218 46102
rect 565274 46046 565342 46102
rect 565398 46046 582970 46102
rect 583026 46046 583094 46102
rect 583150 46046 583218 46102
rect 583274 46046 583342 46102
rect 583398 46046 597456 46102
rect 597512 46046 597580 46102
rect 597636 46046 597704 46102
rect 597760 46046 597828 46102
rect 597884 46046 597980 46102
rect 545484 46040 597980 46046
rect 545484 45984 568022 46040
rect 568078 45984 568146 46040
rect 568202 45984 568270 46040
rect 568326 45984 568394 46040
rect 568450 45984 568518 46040
rect 568574 45984 568642 46040
rect 568698 45984 568766 46040
rect 568822 45984 568890 46040
rect 568946 45984 569014 46040
rect 569070 45984 569138 46040
rect 569194 45984 588022 46040
rect 588078 45984 588146 46040
rect 588202 45984 588270 46040
rect 588326 45984 588394 46040
rect 588450 45984 588518 46040
rect 588574 45984 588642 46040
rect 588698 45984 588766 46040
rect 588822 45984 588890 46040
rect 588946 45984 589014 46040
rect 589070 45984 589138 46040
rect 589194 45984 597980 46040
rect 545484 45978 597980 45984
rect 545484 45922 564970 45978
rect 565026 45922 565094 45978
rect 565150 45922 565218 45978
rect 565274 45922 565342 45978
rect 565398 45922 582970 45978
rect 583026 45922 583094 45978
rect 583150 45922 583218 45978
rect 583274 45922 583342 45978
rect 583398 45922 597456 45978
rect 597512 45922 597580 45978
rect 597636 45922 597704 45978
rect 597760 45922 597828 45978
rect 597884 45922 597980 45978
rect 545484 45916 597980 45922
rect 545484 45860 568022 45916
rect 568078 45860 568146 45916
rect 568202 45860 568270 45916
rect 568326 45860 568394 45916
rect 568450 45860 568518 45916
rect 568574 45860 568642 45916
rect 568698 45860 568766 45916
rect 568822 45860 568890 45916
rect 568946 45860 569014 45916
rect 569070 45860 569138 45916
rect 569194 45860 588022 45916
rect 588078 45860 588146 45916
rect 588202 45860 588270 45916
rect 588326 45860 588394 45916
rect 588450 45860 588518 45916
rect 588574 45860 588642 45916
rect 588698 45860 588766 45916
rect 588822 45860 588890 45916
rect 588946 45860 589014 45916
rect 589070 45860 589138 45916
rect 589194 45860 597980 45916
rect 545484 45826 597980 45860
rect 560236 44578 582164 44594
rect 560236 44522 560252 44578
rect 560308 44522 582092 44578
rect 582148 44522 582164 44578
rect 560236 44506 582164 44522
rect 553964 44218 555396 44234
rect 553964 44162 553980 44218
rect 554036 44162 555324 44218
rect 555380 44162 555396 44218
rect 553964 44146 555396 44162
rect 525292 43138 559428 43154
rect 525292 43082 525308 43138
rect 525364 43082 559356 43138
rect 559412 43082 559428 43138
rect 525292 43066 559428 43082
rect 516444 42958 556964 42974
rect 516444 42902 516460 42958
rect 516516 42902 556892 42958
rect 556948 42902 556964 42958
rect 516444 42886 556964 42902
rect 567740 42958 577124 42974
rect 567740 42902 567756 42958
rect 567812 42902 577052 42958
rect 577108 42902 577124 42958
rect 567740 42886 577124 42902
rect 346764 42778 551140 42794
rect 346764 42722 346780 42778
rect 346836 42722 551068 42778
rect 551124 42722 551140 42778
rect 346764 42706 551140 42722
rect 561916 42778 586532 42794
rect 561916 42722 561932 42778
rect 561988 42722 586460 42778
rect 586516 42722 586532 42778
rect 561916 42706 586532 42722
rect 532684 41518 550356 41534
rect 532684 41462 532700 41518
rect 532756 41462 550284 41518
rect 550340 41462 550356 41518
rect 532684 41446 550356 41462
rect 436252 41338 554612 41354
rect 436252 41282 436268 41338
rect 436324 41282 554540 41338
rect 554596 41282 554612 41338
rect 436252 41266 554612 41282
rect 431772 41158 559988 41174
rect 431772 41102 431788 41158
rect 431844 41102 559916 41158
rect 559972 41102 559988 41158
rect 431772 41086 559988 41102
rect 560124 41158 584852 41174
rect 560124 41102 560140 41158
rect 560196 41102 584780 41158
rect 584836 41102 584852 41158
rect 560124 41086 584852 41102
rect -1916 40350 66564 40446
rect -1916 40294 -860 40350
rect -804 40294 -736 40350
rect -680 40294 -612 40350
rect -556 40294 -488 40350
rect -432 40294 3250 40350
rect 3306 40294 3374 40350
rect 3430 40294 3498 40350
rect 3554 40294 3622 40350
rect 3678 40294 21250 40350
rect 21306 40294 21374 40350
rect 21430 40294 21498 40350
rect 21554 40294 21622 40350
rect 21678 40294 39250 40350
rect 39306 40294 39374 40350
rect 39430 40294 39498 40350
rect 39554 40294 39622 40350
rect 39678 40294 57250 40350
rect 57306 40294 57374 40350
rect 57430 40294 57498 40350
rect 57554 40294 57622 40350
rect 57678 40294 64518 40350
rect 64574 40294 64642 40350
rect 64698 40294 66564 40350
rect -1916 40226 66564 40294
rect -1916 40170 -860 40226
rect -804 40170 -736 40226
rect -680 40170 -612 40226
rect -556 40170 -488 40226
rect -432 40170 3250 40226
rect 3306 40170 3374 40226
rect 3430 40170 3498 40226
rect 3554 40170 3622 40226
rect 3678 40170 21250 40226
rect 21306 40170 21374 40226
rect 21430 40170 21498 40226
rect 21554 40170 21622 40226
rect 21678 40170 39250 40226
rect 39306 40170 39374 40226
rect 39430 40170 39498 40226
rect 39554 40170 39622 40226
rect 39678 40170 57250 40226
rect 57306 40170 57374 40226
rect 57430 40170 57498 40226
rect 57554 40170 57622 40226
rect 57678 40170 64518 40226
rect 64574 40170 64642 40226
rect 64698 40170 66564 40226
rect -1916 40102 66564 40170
rect -1916 40046 -860 40102
rect -804 40046 -736 40102
rect -680 40046 -612 40102
rect -556 40046 -488 40102
rect -432 40046 3250 40102
rect 3306 40046 3374 40102
rect 3430 40046 3498 40102
rect 3554 40046 3622 40102
rect 3678 40046 21250 40102
rect 21306 40046 21374 40102
rect 21430 40046 21498 40102
rect 21554 40046 21622 40102
rect 21678 40046 39250 40102
rect 39306 40046 39374 40102
rect 39430 40046 39498 40102
rect 39554 40046 39622 40102
rect 39678 40046 57250 40102
rect 57306 40046 57374 40102
rect 57430 40046 57498 40102
rect 57554 40046 57622 40102
rect 57678 40046 64518 40102
rect 64574 40046 64642 40102
rect 64698 40046 66564 40102
rect -1916 39978 66564 40046
rect -1916 39922 -860 39978
rect -804 39922 -736 39978
rect -680 39922 -612 39978
rect -556 39922 -488 39978
rect -432 39922 3250 39978
rect 3306 39922 3374 39978
rect 3430 39922 3498 39978
rect 3554 39922 3622 39978
rect 3678 39922 21250 39978
rect 21306 39922 21374 39978
rect 21430 39922 21498 39978
rect 21554 39922 21622 39978
rect 21678 39922 39250 39978
rect 39306 39922 39374 39978
rect 39430 39922 39498 39978
rect 39554 39922 39622 39978
rect 39678 39922 57250 39978
rect 57306 39922 57374 39978
rect 57430 39922 57498 39978
rect 57554 39922 57622 39978
rect 57678 39922 64518 39978
rect 64574 39922 64642 39978
rect 64698 39922 66564 39978
rect -1916 39826 66564 39922
rect 239468 40412 597980 40446
rect 239468 40356 558022 40412
rect 558078 40356 558146 40412
rect 558202 40356 558270 40412
rect 558326 40356 558394 40412
rect 558450 40356 558518 40412
rect 558574 40356 558642 40412
rect 558698 40356 558766 40412
rect 558822 40356 558890 40412
rect 558946 40356 559014 40412
rect 559070 40356 559138 40412
rect 559194 40356 578022 40412
rect 578078 40356 578146 40412
rect 578202 40356 578270 40412
rect 578326 40356 578394 40412
rect 578450 40356 578518 40412
rect 578574 40356 578642 40412
rect 578698 40356 578766 40412
rect 578822 40356 578890 40412
rect 578946 40356 579014 40412
rect 579070 40356 579138 40412
rect 579194 40356 597980 40412
rect 239468 40350 597980 40356
rect 239468 40294 255250 40350
rect 255306 40294 255374 40350
rect 255430 40294 255498 40350
rect 255554 40294 255622 40350
rect 255678 40294 273250 40350
rect 273306 40294 273374 40350
rect 273430 40294 273498 40350
rect 273554 40294 273622 40350
rect 273678 40294 291250 40350
rect 291306 40294 291374 40350
rect 291430 40294 291498 40350
rect 291554 40294 291622 40350
rect 291678 40294 309250 40350
rect 309306 40294 309374 40350
rect 309430 40294 309498 40350
rect 309554 40294 309622 40350
rect 309678 40294 327250 40350
rect 327306 40294 327374 40350
rect 327430 40294 327498 40350
rect 327554 40294 327622 40350
rect 327678 40294 345250 40350
rect 345306 40294 345374 40350
rect 345430 40294 345498 40350
rect 345554 40294 345622 40350
rect 345678 40294 363250 40350
rect 363306 40294 363374 40350
rect 363430 40294 363498 40350
rect 363554 40294 363622 40350
rect 363678 40294 381250 40350
rect 381306 40294 381374 40350
rect 381430 40294 381498 40350
rect 381554 40294 381622 40350
rect 381678 40294 399250 40350
rect 399306 40294 399374 40350
rect 399430 40294 399498 40350
rect 399554 40294 399622 40350
rect 399678 40294 417250 40350
rect 417306 40294 417374 40350
rect 417430 40294 417498 40350
rect 417554 40294 417622 40350
rect 417678 40294 435250 40350
rect 435306 40294 435374 40350
rect 435430 40294 435498 40350
rect 435554 40294 435622 40350
rect 435678 40294 453250 40350
rect 453306 40294 453374 40350
rect 453430 40294 453498 40350
rect 453554 40294 453622 40350
rect 453678 40294 471250 40350
rect 471306 40294 471374 40350
rect 471430 40294 471498 40350
rect 471554 40294 471622 40350
rect 471678 40294 489250 40350
rect 489306 40294 489374 40350
rect 489430 40294 489498 40350
rect 489554 40294 489622 40350
rect 489678 40294 507250 40350
rect 507306 40294 507374 40350
rect 507430 40294 507498 40350
rect 507554 40294 507622 40350
rect 507678 40294 525250 40350
rect 525306 40294 525374 40350
rect 525430 40294 525498 40350
rect 525554 40294 525622 40350
rect 525678 40294 543250 40350
rect 543306 40294 543374 40350
rect 543430 40294 543498 40350
rect 543554 40294 543622 40350
rect 543678 40294 561250 40350
rect 561306 40294 561374 40350
rect 561430 40294 561498 40350
rect 561554 40294 561622 40350
rect 561678 40294 596496 40350
rect 596552 40294 596620 40350
rect 596676 40294 596744 40350
rect 596800 40294 596868 40350
rect 596924 40294 597980 40350
rect 239468 40288 597980 40294
rect 239468 40232 558022 40288
rect 558078 40232 558146 40288
rect 558202 40232 558270 40288
rect 558326 40232 558394 40288
rect 558450 40232 558518 40288
rect 558574 40232 558642 40288
rect 558698 40232 558766 40288
rect 558822 40232 558890 40288
rect 558946 40232 559014 40288
rect 559070 40232 559138 40288
rect 559194 40232 578022 40288
rect 578078 40232 578146 40288
rect 578202 40232 578270 40288
rect 578326 40232 578394 40288
rect 578450 40232 578518 40288
rect 578574 40232 578642 40288
rect 578698 40232 578766 40288
rect 578822 40232 578890 40288
rect 578946 40232 579014 40288
rect 579070 40232 579138 40288
rect 579194 40232 597980 40288
rect 239468 40226 597980 40232
rect 239468 40170 255250 40226
rect 255306 40170 255374 40226
rect 255430 40170 255498 40226
rect 255554 40170 255622 40226
rect 255678 40170 273250 40226
rect 273306 40170 273374 40226
rect 273430 40170 273498 40226
rect 273554 40170 273622 40226
rect 273678 40170 291250 40226
rect 291306 40170 291374 40226
rect 291430 40170 291498 40226
rect 291554 40170 291622 40226
rect 291678 40170 309250 40226
rect 309306 40170 309374 40226
rect 309430 40170 309498 40226
rect 309554 40170 309622 40226
rect 309678 40170 327250 40226
rect 327306 40170 327374 40226
rect 327430 40170 327498 40226
rect 327554 40170 327622 40226
rect 327678 40170 345250 40226
rect 345306 40170 345374 40226
rect 345430 40170 345498 40226
rect 345554 40170 345622 40226
rect 345678 40170 363250 40226
rect 363306 40170 363374 40226
rect 363430 40170 363498 40226
rect 363554 40170 363622 40226
rect 363678 40170 381250 40226
rect 381306 40170 381374 40226
rect 381430 40170 381498 40226
rect 381554 40170 381622 40226
rect 381678 40170 399250 40226
rect 399306 40170 399374 40226
rect 399430 40170 399498 40226
rect 399554 40170 399622 40226
rect 399678 40170 417250 40226
rect 417306 40170 417374 40226
rect 417430 40170 417498 40226
rect 417554 40170 417622 40226
rect 417678 40170 435250 40226
rect 435306 40170 435374 40226
rect 435430 40170 435498 40226
rect 435554 40170 435622 40226
rect 435678 40170 453250 40226
rect 453306 40170 453374 40226
rect 453430 40170 453498 40226
rect 453554 40170 453622 40226
rect 453678 40170 471250 40226
rect 471306 40170 471374 40226
rect 471430 40170 471498 40226
rect 471554 40170 471622 40226
rect 471678 40170 489250 40226
rect 489306 40170 489374 40226
rect 489430 40170 489498 40226
rect 489554 40170 489622 40226
rect 489678 40170 507250 40226
rect 507306 40170 507374 40226
rect 507430 40170 507498 40226
rect 507554 40170 507622 40226
rect 507678 40170 525250 40226
rect 525306 40170 525374 40226
rect 525430 40170 525498 40226
rect 525554 40170 525622 40226
rect 525678 40170 543250 40226
rect 543306 40170 543374 40226
rect 543430 40170 543498 40226
rect 543554 40170 543622 40226
rect 543678 40170 561250 40226
rect 561306 40170 561374 40226
rect 561430 40170 561498 40226
rect 561554 40170 561622 40226
rect 561678 40170 596496 40226
rect 596552 40170 596620 40226
rect 596676 40170 596744 40226
rect 596800 40170 596868 40226
rect 596924 40170 597980 40226
rect 239468 40164 597980 40170
rect 239468 40108 558022 40164
rect 558078 40108 558146 40164
rect 558202 40108 558270 40164
rect 558326 40108 558394 40164
rect 558450 40108 558518 40164
rect 558574 40108 558642 40164
rect 558698 40108 558766 40164
rect 558822 40108 558890 40164
rect 558946 40108 559014 40164
rect 559070 40108 559138 40164
rect 559194 40108 578022 40164
rect 578078 40108 578146 40164
rect 578202 40108 578270 40164
rect 578326 40108 578394 40164
rect 578450 40108 578518 40164
rect 578574 40108 578642 40164
rect 578698 40108 578766 40164
rect 578822 40108 578890 40164
rect 578946 40108 579014 40164
rect 579070 40108 579138 40164
rect 579194 40108 597980 40164
rect 239468 40102 597980 40108
rect 239468 40046 255250 40102
rect 255306 40046 255374 40102
rect 255430 40046 255498 40102
rect 255554 40046 255622 40102
rect 255678 40046 273250 40102
rect 273306 40046 273374 40102
rect 273430 40046 273498 40102
rect 273554 40046 273622 40102
rect 273678 40046 291250 40102
rect 291306 40046 291374 40102
rect 291430 40046 291498 40102
rect 291554 40046 291622 40102
rect 291678 40046 309250 40102
rect 309306 40046 309374 40102
rect 309430 40046 309498 40102
rect 309554 40046 309622 40102
rect 309678 40046 327250 40102
rect 327306 40046 327374 40102
rect 327430 40046 327498 40102
rect 327554 40046 327622 40102
rect 327678 40046 345250 40102
rect 345306 40046 345374 40102
rect 345430 40046 345498 40102
rect 345554 40046 345622 40102
rect 345678 40046 363250 40102
rect 363306 40046 363374 40102
rect 363430 40046 363498 40102
rect 363554 40046 363622 40102
rect 363678 40046 381250 40102
rect 381306 40046 381374 40102
rect 381430 40046 381498 40102
rect 381554 40046 381622 40102
rect 381678 40046 399250 40102
rect 399306 40046 399374 40102
rect 399430 40046 399498 40102
rect 399554 40046 399622 40102
rect 399678 40046 417250 40102
rect 417306 40046 417374 40102
rect 417430 40046 417498 40102
rect 417554 40046 417622 40102
rect 417678 40046 435250 40102
rect 435306 40046 435374 40102
rect 435430 40046 435498 40102
rect 435554 40046 435622 40102
rect 435678 40046 453250 40102
rect 453306 40046 453374 40102
rect 453430 40046 453498 40102
rect 453554 40046 453622 40102
rect 453678 40046 471250 40102
rect 471306 40046 471374 40102
rect 471430 40046 471498 40102
rect 471554 40046 471622 40102
rect 471678 40046 489250 40102
rect 489306 40046 489374 40102
rect 489430 40046 489498 40102
rect 489554 40046 489622 40102
rect 489678 40046 507250 40102
rect 507306 40046 507374 40102
rect 507430 40046 507498 40102
rect 507554 40046 507622 40102
rect 507678 40046 525250 40102
rect 525306 40046 525374 40102
rect 525430 40046 525498 40102
rect 525554 40046 525622 40102
rect 525678 40046 543250 40102
rect 543306 40046 543374 40102
rect 543430 40046 543498 40102
rect 543554 40046 543622 40102
rect 543678 40046 561250 40102
rect 561306 40046 561374 40102
rect 561430 40046 561498 40102
rect 561554 40046 561622 40102
rect 561678 40046 596496 40102
rect 596552 40046 596620 40102
rect 596676 40046 596744 40102
rect 596800 40046 596868 40102
rect 596924 40046 597980 40102
rect 239468 40040 597980 40046
rect 239468 39984 558022 40040
rect 558078 39984 558146 40040
rect 558202 39984 558270 40040
rect 558326 39984 558394 40040
rect 558450 39984 558518 40040
rect 558574 39984 558642 40040
rect 558698 39984 558766 40040
rect 558822 39984 558890 40040
rect 558946 39984 559014 40040
rect 559070 39984 559138 40040
rect 559194 39984 578022 40040
rect 578078 39984 578146 40040
rect 578202 39984 578270 40040
rect 578326 39984 578394 40040
rect 578450 39984 578518 40040
rect 578574 39984 578642 40040
rect 578698 39984 578766 40040
rect 578822 39984 578890 40040
rect 578946 39984 579014 40040
rect 579070 39984 579138 40040
rect 579194 39984 597980 40040
rect 239468 39978 597980 39984
rect 239468 39922 255250 39978
rect 255306 39922 255374 39978
rect 255430 39922 255498 39978
rect 255554 39922 255622 39978
rect 255678 39922 273250 39978
rect 273306 39922 273374 39978
rect 273430 39922 273498 39978
rect 273554 39922 273622 39978
rect 273678 39922 291250 39978
rect 291306 39922 291374 39978
rect 291430 39922 291498 39978
rect 291554 39922 291622 39978
rect 291678 39922 309250 39978
rect 309306 39922 309374 39978
rect 309430 39922 309498 39978
rect 309554 39922 309622 39978
rect 309678 39922 327250 39978
rect 327306 39922 327374 39978
rect 327430 39922 327498 39978
rect 327554 39922 327622 39978
rect 327678 39922 345250 39978
rect 345306 39922 345374 39978
rect 345430 39922 345498 39978
rect 345554 39922 345622 39978
rect 345678 39922 363250 39978
rect 363306 39922 363374 39978
rect 363430 39922 363498 39978
rect 363554 39922 363622 39978
rect 363678 39922 381250 39978
rect 381306 39922 381374 39978
rect 381430 39922 381498 39978
rect 381554 39922 381622 39978
rect 381678 39922 399250 39978
rect 399306 39922 399374 39978
rect 399430 39922 399498 39978
rect 399554 39922 399622 39978
rect 399678 39922 417250 39978
rect 417306 39922 417374 39978
rect 417430 39922 417498 39978
rect 417554 39922 417622 39978
rect 417678 39922 435250 39978
rect 435306 39922 435374 39978
rect 435430 39922 435498 39978
rect 435554 39922 435622 39978
rect 435678 39922 453250 39978
rect 453306 39922 453374 39978
rect 453430 39922 453498 39978
rect 453554 39922 453622 39978
rect 453678 39922 471250 39978
rect 471306 39922 471374 39978
rect 471430 39922 471498 39978
rect 471554 39922 471622 39978
rect 471678 39922 489250 39978
rect 489306 39922 489374 39978
rect 489430 39922 489498 39978
rect 489554 39922 489622 39978
rect 489678 39922 507250 39978
rect 507306 39922 507374 39978
rect 507430 39922 507498 39978
rect 507554 39922 507622 39978
rect 507678 39922 525250 39978
rect 525306 39922 525374 39978
rect 525430 39922 525498 39978
rect 525554 39922 525622 39978
rect 525678 39922 543250 39978
rect 543306 39922 543374 39978
rect 543430 39922 543498 39978
rect 543554 39922 543622 39978
rect 543678 39922 561250 39978
rect 561306 39922 561374 39978
rect 561430 39922 561498 39978
rect 561554 39922 561622 39978
rect 561678 39922 596496 39978
rect 596552 39922 596620 39978
rect 596676 39922 596744 39978
rect 596800 39922 596868 39978
rect 596924 39922 597980 39978
rect 239468 39916 597980 39922
rect 239468 39860 558022 39916
rect 558078 39860 558146 39916
rect 558202 39860 558270 39916
rect 558326 39860 558394 39916
rect 558450 39860 558518 39916
rect 558574 39860 558642 39916
rect 558698 39860 558766 39916
rect 558822 39860 558890 39916
rect 558946 39860 559014 39916
rect 559070 39860 559138 39916
rect 559194 39860 578022 39916
rect 578078 39860 578146 39916
rect 578202 39860 578270 39916
rect 578326 39860 578394 39916
rect 578450 39860 578518 39916
rect 578574 39860 578642 39916
rect 578698 39860 578766 39916
rect 578822 39860 578890 39916
rect 578946 39860 579014 39916
rect 579070 39860 579138 39916
rect 579194 39860 597980 39916
rect 239468 39826 597980 39860
rect 418332 39718 560100 39734
rect 418332 39662 418348 39718
rect 418404 39662 419692 39718
rect 419748 39662 560028 39718
rect 560084 39662 560100 39718
rect 418332 39646 560100 39662
rect 451932 39538 559876 39554
rect 451932 39482 451948 39538
rect 452004 39482 559804 39538
rect 559860 39482 559876 39538
rect 451932 39466 559876 39482
rect 459996 39358 559764 39374
rect 459996 39302 460012 39358
rect 460068 39302 559692 39358
rect 559748 39302 559764 39358
rect 459996 39286 559764 39302
rect 565724 38638 573764 38654
rect 565724 38582 565740 38638
rect 565796 38582 573692 38638
rect 573748 38582 573764 38638
rect 565724 38566 573764 38582
rect 550828 38098 557300 38114
rect 550828 38042 550844 38098
rect 550900 38042 557228 38098
rect 557284 38042 557300 38098
rect 550828 38026 557300 38042
rect 546012 37918 554388 37934
rect 546012 37862 546028 37918
rect 546084 37862 554388 37918
rect 546012 37846 554388 37862
rect 554524 37918 560212 37934
rect 554524 37862 554540 37918
rect 554596 37862 560140 37918
rect 560196 37862 560212 37918
rect 554524 37846 560212 37862
rect 554300 37754 554388 37846
rect 354492 37738 549404 37754
rect 354492 37682 354508 37738
rect 354564 37682 549404 37738
rect 354492 37666 549404 37682
rect 554300 37738 557076 37754
rect 554300 37682 557004 37738
rect 557060 37682 557076 37738
rect 554300 37666 557076 37682
rect 557324 37738 557412 37754
rect 557324 37682 557340 37738
rect 557396 37682 557412 37738
rect 549316 37574 549404 37666
rect 557324 37574 557412 37682
rect 565612 37738 581492 37754
rect 565612 37682 565628 37738
rect 565684 37682 581420 37738
rect 581476 37682 581492 37738
rect 565612 37666 581492 37682
rect 549316 37486 557412 37574
rect 362892 37018 577236 37034
rect 362892 36962 362908 37018
rect 362964 36962 572908 37018
rect 572964 36962 577164 37018
rect 577220 36962 577236 37018
rect 362892 36946 577236 36962
rect 554300 36838 567044 36854
rect 554300 36782 554316 36838
rect 554372 36782 566972 36838
rect 567028 36782 567044 36838
rect 554300 36766 567044 36782
rect 423372 35218 549348 35234
rect 423372 35162 423388 35218
rect 423444 35162 549276 35218
rect 549332 35162 549348 35218
rect 423372 35146 549348 35162
rect 238460 34498 418420 34514
rect 238460 34442 238476 34498
rect 238532 34442 418348 34498
rect 418404 34442 418420 34498
rect 238460 34426 418420 34442
rect 153452 33238 512500 33254
rect 153452 33182 153468 33238
rect 153524 33182 512428 33238
rect 512484 33182 512500 33238
rect 153452 33166 512500 33182
rect 158828 33058 524596 33074
rect 158828 33002 158844 33058
rect 158900 33002 524524 33058
rect 524580 33002 524596 33058
rect 158828 32986 524596 33002
rect 160620 32878 528628 32894
rect 160620 32822 160636 32878
rect 160692 32822 528556 32878
rect 528612 32822 528628 32878
rect 160620 32806 528628 32822
rect 162412 32698 532660 32714
rect 162412 32642 162428 32698
rect 162484 32642 532588 32698
rect 532644 32642 532660 32698
rect 162412 32626 532660 32642
rect 140796 31798 463780 31814
rect 140796 31742 140812 31798
rect 140868 31742 463708 31798
rect 463764 31742 463780 31798
rect 140796 31726 463780 31742
rect 139116 31618 478900 31634
rect 139116 31562 139132 31618
rect 139188 31562 478828 31618
rect 478884 31562 478900 31618
rect 139116 31546 478900 31562
rect 140908 31438 483940 31454
rect 140908 31382 140924 31438
rect 140980 31382 483868 31438
rect 483924 31382 483940 31438
rect 140908 31366 483940 31382
rect 142700 31258 487300 31274
rect 142700 31202 142716 31258
rect 142772 31202 487228 31258
rect 487284 31202 487300 31258
rect 142700 31186 487300 31202
rect 149868 31078 504884 31094
rect 149868 31022 149884 31078
rect 149940 31022 504812 31078
rect 504868 31022 504884 31078
rect 149868 31006 504884 31022
rect 157036 30178 519220 30194
rect 157036 30122 157052 30178
rect 157108 30122 519148 30178
rect 519204 30122 519220 30178
rect 157036 30106 519220 30122
rect 591260 30178 593364 30194
rect 591260 30122 591276 30178
rect 591332 30122 593292 30178
rect 593348 30122 593364 30178
rect 591260 30106 593364 30122
rect 155244 29998 516532 30014
rect 155244 29942 155260 29998
rect 155316 29942 516460 29998
rect 516516 29942 516532 29998
rect 155244 29926 516532 29942
rect 147852 29818 500404 29834
rect 147852 29762 147868 29818
rect 147924 29762 500332 29818
rect 500388 29762 500404 29818
rect 147852 29746 500404 29762
rect 221548 29638 244484 29654
rect 221548 29582 221564 29638
rect 221620 29582 244412 29638
rect 244468 29582 244484 29638
rect 221548 29566 244484 29582
rect 394812 29638 557860 29654
rect 394812 29582 394828 29638
rect 394884 29582 557788 29638
rect 557844 29582 557860 29638
rect 394812 29566 557860 29582
rect 186492 29458 431860 29474
rect 186492 29402 186508 29458
rect 186564 29402 431788 29458
rect 431844 29402 431860 29458
rect 186492 29386 431860 29402
rect 554524 29458 565812 29474
rect 554524 29402 554540 29458
rect 554596 29402 556892 29458
rect 556948 29402 565740 29458
rect 565796 29402 565812 29458
rect 554524 29386 565812 29402
rect -1916 28412 597980 28446
rect -1916 28356 568022 28412
rect 568078 28356 568146 28412
rect 568202 28356 568270 28412
rect 568326 28356 568394 28412
rect 568450 28356 568518 28412
rect 568574 28356 568642 28412
rect 568698 28356 568766 28412
rect 568822 28356 568890 28412
rect 568946 28356 569014 28412
rect 569070 28356 569138 28412
rect 569194 28356 588022 28412
rect 588078 28356 588146 28412
rect 588202 28356 588270 28412
rect 588326 28356 588394 28412
rect 588450 28356 588518 28412
rect 588574 28356 588642 28412
rect 588698 28356 588766 28412
rect 588822 28356 588890 28412
rect 588946 28356 589014 28412
rect 589070 28356 589138 28412
rect 589194 28356 597980 28412
rect -1916 28350 597980 28356
rect -1916 28294 -1820 28350
rect -1764 28294 -1696 28350
rect -1640 28294 -1572 28350
rect -1516 28294 -1448 28350
rect -1392 28294 6970 28350
rect 7026 28294 7094 28350
rect 7150 28294 7218 28350
rect 7274 28294 7342 28350
rect 7398 28294 24970 28350
rect 25026 28294 25094 28350
rect 25150 28294 25218 28350
rect 25274 28294 25342 28350
rect 25398 28294 42970 28350
rect 43026 28294 43094 28350
rect 43150 28294 43218 28350
rect 43274 28294 43342 28350
rect 43398 28294 60970 28350
rect 61026 28294 61094 28350
rect 61150 28294 61218 28350
rect 61274 28294 61342 28350
rect 61398 28294 78970 28350
rect 79026 28294 79094 28350
rect 79150 28294 79218 28350
rect 79274 28294 79342 28350
rect 79398 28294 96970 28350
rect 97026 28294 97094 28350
rect 97150 28294 97218 28350
rect 97274 28294 97342 28350
rect 97398 28294 114970 28350
rect 115026 28294 115094 28350
rect 115150 28294 115218 28350
rect 115274 28294 115342 28350
rect 115398 28294 132970 28350
rect 133026 28294 133094 28350
rect 133150 28294 133218 28350
rect 133274 28294 133342 28350
rect 133398 28294 150970 28350
rect 151026 28294 151094 28350
rect 151150 28294 151218 28350
rect 151274 28294 151342 28350
rect 151398 28294 168970 28350
rect 169026 28294 169094 28350
rect 169150 28294 169218 28350
rect 169274 28294 169342 28350
rect 169398 28294 186970 28350
rect 187026 28294 187094 28350
rect 187150 28294 187218 28350
rect 187274 28294 187342 28350
rect 187398 28294 204970 28350
rect 205026 28294 205094 28350
rect 205150 28294 205218 28350
rect 205274 28294 205342 28350
rect 205398 28294 222970 28350
rect 223026 28294 223094 28350
rect 223150 28294 223218 28350
rect 223274 28294 223342 28350
rect 223398 28294 240970 28350
rect 241026 28294 241094 28350
rect 241150 28294 241218 28350
rect 241274 28294 241342 28350
rect 241398 28294 258970 28350
rect 259026 28294 259094 28350
rect 259150 28294 259218 28350
rect 259274 28294 259342 28350
rect 259398 28294 276970 28350
rect 277026 28294 277094 28350
rect 277150 28294 277218 28350
rect 277274 28294 277342 28350
rect 277398 28294 294970 28350
rect 295026 28294 295094 28350
rect 295150 28294 295218 28350
rect 295274 28294 295342 28350
rect 295398 28294 312970 28350
rect 313026 28294 313094 28350
rect 313150 28294 313218 28350
rect 313274 28294 313342 28350
rect 313398 28294 330970 28350
rect 331026 28294 331094 28350
rect 331150 28294 331218 28350
rect 331274 28294 331342 28350
rect 331398 28294 348970 28350
rect 349026 28294 349094 28350
rect 349150 28294 349218 28350
rect 349274 28294 349342 28350
rect 349398 28294 366970 28350
rect 367026 28294 367094 28350
rect 367150 28294 367218 28350
rect 367274 28294 367342 28350
rect 367398 28294 384970 28350
rect 385026 28294 385094 28350
rect 385150 28294 385218 28350
rect 385274 28294 385342 28350
rect 385398 28294 402970 28350
rect 403026 28294 403094 28350
rect 403150 28294 403218 28350
rect 403274 28294 403342 28350
rect 403398 28294 420970 28350
rect 421026 28294 421094 28350
rect 421150 28294 421218 28350
rect 421274 28294 421342 28350
rect 421398 28294 438970 28350
rect 439026 28294 439094 28350
rect 439150 28294 439218 28350
rect 439274 28294 439342 28350
rect 439398 28294 456970 28350
rect 457026 28294 457094 28350
rect 457150 28294 457218 28350
rect 457274 28294 457342 28350
rect 457398 28294 474970 28350
rect 475026 28294 475094 28350
rect 475150 28294 475218 28350
rect 475274 28294 475342 28350
rect 475398 28294 492970 28350
rect 493026 28294 493094 28350
rect 493150 28294 493218 28350
rect 493274 28294 493342 28350
rect 493398 28294 510970 28350
rect 511026 28294 511094 28350
rect 511150 28294 511218 28350
rect 511274 28294 511342 28350
rect 511398 28294 528970 28350
rect 529026 28294 529094 28350
rect 529150 28294 529218 28350
rect 529274 28294 529342 28350
rect 529398 28294 546970 28350
rect 547026 28294 547094 28350
rect 547150 28294 547218 28350
rect 547274 28294 547342 28350
rect 547398 28294 564970 28350
rect 565026 28294 565094 28350
rect 565150 28294 565218 28350
rect 565274 28294 565342 28350
rect 565398 28294 582970 28350
rect 583026 28294 583094 28350
rect 583150 28294 583218 28350
rect 583274 28294 583342 28350
rect 583398 28294 597456 28350
rect 597512 28294 597580 28350
rect 597636 28294 597704 28350
rect 597760 28294 597828 28350
rect 597884 28294 597980 28350
rect -1916 28288 597980 28294
rect -1916 28232 568022 28288
rect 568078 28232 568146 28288
rect 568202 28232 568270 28288
rect 568326 28232 568394 28288
rect 568450 28232 568518 28288
rect 568574 28232 568642 28288
rect 568698 28232 568766 28288
rect 568822 28232 568890 28288
rect 568946 28232 569014 28288
rect 569070 28232 569138 28288
rect 569194 28232 588022 28288
rect 588078 28232 588146 28288
rect 588202 28232 588270 28288
rect 588326 28232 588394 28288
rect 588450 28232 588518 28288
rect 588574 28232 588642 28288
rect 588698 28232 588766 28288
rect 588822 28232 588890 28288
rect 588946 28232 589014 28288
rect 589070 28232 589138 28288
rect 589194 28232 597980 28288
rect -1916 28226 597980 28232
rect -1916 28170 -1820 28226
rect -1764 28170 -1696 28226
rect -1640 28170 -1572 28226
rect -1516 28170 -1448 28226
rect -1392 28170 6970 28226
rect 7026 28170 7094 28226
rect 7150 28170 7218 28226
rect 7274 28170 7342 28226
rect 7398 28170 24970 28226
rect 25026 28170 25094 28226
rect 25150 28170 25218 28226
rect 25274 28170 25342 28226
rect 25398 28170 42970 28226
rect 43026 28170 43094 28226
rect 43150 28170 43218 28226
rect 43274 28170 43342 28226
rect 43398 28170 60970 28226
rect 61026 28170 61094 28226
rect 61150 28170 61218 28226
rect 61274 28170 61342 28226
rect 61398 28170 78970 28226
rect 79026 28170 79094 28226
rect 79150 28170 79218 28226
rect 79274 28170 79342 28226
rect 79398 28170 96970 28226
rect 97026 28170 97094 28226
rect 97150 28170 97218 28226
rect 97274 28170 97342 28226
rect 97398 28170 114970 28226
rect 115026 28170 115094 28226
rect 115150 28170 115218 28226
rect 115274 28170 115342 28226
rect 115398 28170 132970 28226
rect 133026 28170 133094 28226
rect 133150 28170 133218 28226
rect 133274 28170 133342 28226
rect 133398 28170 150970 28226
rect 151026 28170 151094 28226
rect 151150 28170 151218 28226
rect 151274 28170 151342 28226
rect 151398 28170 168970 28226
rect 169026 28170 169094 28226
rect 169150 28170 169218 28226
rect 169274 28170 169342 28226
rect 169398 28170 186970 28226
rect 187026 28170 187094 28226
rect 187150 28170 187218 28226
rect 187274 28170 187342 28226
rect 187398 28170 204970 28226
rect 205026 28170 205094 28226
rect 205150 28170 205218 28226
rect 205274 28170 205342 28226
rect 205398 28170 222970 28226
rect 223026 28170 223094 28226
rect 223150 28170 223218 28226
rect 223274 28170 223342 28226
rect 223398 28170 240970 28226
rect 241026 28170 241094 28226
rect 241150 28170 241218 28226
rect 241274 28170 241342 28226
rect 241398 28170 258970 28226
rect 259026 28170 259094 28226
rect 259150 28170 259218 28226
rect 259274 28170 259342 28226
rect 259398 28170 276970 28226
rect 277026 28170 277094 28226
rect 277150 28170 277218 28226
rect 277274 28170 277342 28226
rect 277398 28170 294970 28226
rect 295026 28170 295094 28226
rect 295150 28170 295218 28226
rect 295274 28170 295342 28226
rect 295398 28170 312970 28226
rect 313026 28170 313094 28226
rect 313150 28170 313218 28226
rect 313274 28170 313342 28226
rect 313398 28170 330970 28226
rect 331026 28170 331094 28226
rect 331150 28170 331218 28226
rect 331274 28170 331342 28226
rect 331398 28170 348970 28226
rect 349026 28170 349094 28226
rect 349150 28170 349218 28226
rect 349274 28170 349342 28226
rect 349398 28170 366970 28226
rect 367026 28170 367094 28226
rect 367150 28170 367218 28226
rect 367274 28170 367342 28226
rect 367398 28170 384970 28226
rect 385026 28170 385094 28226
rect 385150 28170 385218 28226
rect 385274 28170 385342 28226
rect 385398 28170 402970 28226
rect 403026 28170 403094 28226
rect 403150 28170 403218 28226
rect 403274 28170 403342 28226
rect 403398 28170 420970 28226
rect 421026 28170 421094 28226
rect 421150 28170 421218 28226
rect 421274 28170 421342 28226
rect 421398 28170 438970 28226
rect 439026 28170 439094 28226
rect 439150 28170 439218 28226
rect 439274 28170 439342 28226
rect 439398 28170 456970 28226
rect 457026 28170 457094 28226
rect 457150 28170 457218 28226
rect 457274 28170 457342 28226
rect 457398 28170 474970 28226
rect 475026 28170 475094 28226
rect 475150 28170 475218 28226
rect 475274 28170 475342 28226
rect 475398 28170 492970 28226
rect 493026 28170 493094 28226
rect 493150 28170 493218 28226
rect 493274 28170 493342 28226
rect 493398 28170 510970 28226
rect 511026 28170 511094 28226
rect 511150 28170 511218 28226
rect 511274 28170 511342 28226
rect 511398 28170 528970 28226
rect 529026 28170 529094 28226
rect 529150 28170 529218 28226
rect 529274 28170 529342 28226
rect 529398 28170 546970 28226
rect 547026 28170 547094 28226
rect 547150 28170 547218 28226
rect 547274 28170 547342 28226
rect 547398 28170 564970 28226
rect 565026 28170 565094 28226
rect 565150 28170 565218 28226
rect 565274 28170 565342 28226
rect 565398 28170 582970 28226
rect 583026 28170 583094 28226
rect 583150 28170 583218 28226
rect 583274 28170 583342 28226
rect 583398 28170 597456 28226
rect 597512 28170 597580 28226
rect 597636 28170 597704 28226
rect 597760 28170 597828 28226
rect 597884 28170 597980 28226
rect -1916 28164 597980 28170
rect -1916 28108 568022 28164
rect 568078 28108 568146 28164
rect 568202 28108 568270 28164
rect 568326 28108 568394 28164
rect 568450 28108 568518 28164
rect 568574 28108 568642 28164
rect 568698 28108 568766 28164
rect 568822 28108 568890 28164
rect 568946 28108 569014 28164
rect 569070 28108 569138 28164
rect 569194 28108 588022 28164
rect 588078 28108 588146 28164
rect 588202 28108 588270 28164
rect 588326 28108 588394 28164
rect 588450 28108 588518 28164
rect 588574 28108 588642 28164
rect 588698 28108 588766 28164
rect 588822 28108 588890 28164
rect 588946 28108 589014 28164
rect 589070 28108 589138 28164
rect 589194 28108 597980 28164
rect -1916 28102 597980 28108
rect -1916 28046 -1820 28102
rect -1764 28046 -1696 28102
rect -1640 28046 -1572 28102
rect -1516 28046 -1448 28102
rect -1392 28046 6970 28102
rect 7026 28046 7094 28102
rect 7150 28046 7218 28102
rect 7274 28046 7342 28102
rect 7398 28046 24970 28102
rect 25026 28046 25094 28102
rect 25150 28046 25218 28102
rect 25274 28046 25342 28102
rect 25398 28046 42970 28102
rect 43026 28046 43094 28102
rect 43150 28046 43218 28102
rect 43274 28046 43342 28102
rect 43398 28046 60970 28102
rect 61026 28046 61094 28102
rect 61150 28046 61218 28102
rect 61274 28046 61342 28102
rect 61398 28046 78970 28102
rect 79026 28046 79094 28102
rect 79150 28046 79218 28102
rect 79274 28046 79342 28102
rect 79398 28046 96970 28102
rect 97026 28046 97094 28102
rect 97150 28046 97218 28102
rect 97274 28046 97342 28102
rect 97398 28046 114970 28102
rect 115026 28046 115094 28102
rect 115150 28046 115218 28102
rect 115274 28046 115342 28102
rect 115398 28046 132970 28102
rect 133026 28046 133094 28102
rect 133150 28046 133218 28102
rect 133274 28046 133342 28102
rect 133398 28046 150970 28102
rect 151026 28046 151094 28102
rect 151150 28046 151218 28102
rect 151274 28046 151342 28102
rect 151398 28046 168970 28102
rect 169026 28046 169094 28102
rect 169150 28046 169218 28102
rect 169274 28046 169342 28102
rect 169398 28046 186970 28102
rect 187026 28046 187094 28102
rect 187150 28046 187218 28102
rect 187274 28046 187342 28102
rect 187398 28046 204970 28102
rect 205026 28046 205094 28102
rect 205150 28046 205218 28102
rect 205274 28046 205342 28102
rect 205398 28046 222970 28102
rect 223026 28046 223094 28102
rect 223150 28046 223218 28102
rect 223274 28046 223342 28102
rect 223398 28046 240970 28102
rect 241026 28046 241094 28102
rect 241150 28046 241218 28102
rect 241274 28046 241342 28102
rect 241398 28046 258970 28102
rect 259026 28046 259094 28102
rect 259150 28046 259218 28102
rect 259274 28046 259342 28102
rect 259398 28046 276970 28102
rect 277026 28046 277094 28102
rect 277150 28046 277218 28102
rect 277274 28046 277342 28102
rect 277398 28046 294970 28102
rect 295026 28046 295094 28102
rect 295150 28046 295218 28102
rect 295274 28046 295342 28102
rect 295398 28046 312970 28102
rect 313026 28046 313094 28102
rect 313150 28046 313218 28102
rect 313274 28046 313342 28102
rect 313398 28046 330970 28102
rect 331026 28046 331094 28102
rect 331150 28046 331218 28102
rect 331274 28046 331342 28102
rect 331398 28046 348970 28102
rect 349026 28046 349094 28102
rect 349150 28046 349218 28102
rect 349274 28046 349342 28102
rect 349398 28046 366970 28102
rect 367026 28046 367094 28102
rect 367150 28046 367218 28102
rect 367274 28046 367342 28102
rect 367398 28046 384970 28102
rect 385026 28046 385094 28102
rect 385150 28046 385218 28102
rect 385274 28046 385342 28102
rect 385398 28046 402970 28102
rect 403026 28046 403094 28102
rect 403150 28046 403218 28102
rect 403274 28046 403342 28102
rect 403398 28046 420970 28102
rect 421026 28046 421094 28102
rect 421150 28046 421218 28102
rect 421274 28046 421342 28102
rect 421398 28046 438970 28102
rect 439026 28046 439094 28102
rect 439150 28046 439218 28102
rect 439274 28046 439342 28102
rect 439398 28046 456970 28102
rect 457026 28046 457094 28102
rect 457150 28046 457218 28102
rect 457274 28046 457342 28102
rect 457398 28046 474970 28102
rect 475026 28046 475094 28102
rect 475150 28046 475218 28102
rect 475274 28046 475342 28102
rect 475398 28046 492970 28102
rect 493026 28046 493094 28102
rect 493150 28046 493218 28102
rect 493274 28046 493342 28102
rect 493398 28046 510970 28102
rect 511026 28046 511094 28102
rect 511150 28046 511218 28102
rect 511274 28046 511342 28102
rect 511398 28046 528970 28102
rect 529026 28046 529094 28102
rect 529150 28046 529218 28102
rect 529274 28046 529342 28102
rect 529398 28046 546970 28102
rect 547026 28046 547094 28102
rect 547150 28046 547218 28102
rect 547274 28046 547342 28102
rect 547398 28046 564970 28102
rect 565026 28046 565094 28102
rect 565150 28046 565218 28102
rect 565274 28046 565342 28102
rect 565398 28046 582970 28102
rect 583026 28046 583094 28102
rect 583150 28046 583218 28102
rect 583274 28046 583342 28102
rect 583398 28046 597456 28102
rect 597512 28046 597580 28102
rect 597636 28046 597704 28102
rect 597760 28046 597828 28102
rect 597884 28046 597980 28102
rect -1916 28040 597980 28046
rect -1916 27984 568022 28040
rect 568078 27984 568146 28040
rect 568202 27984 568270 28040
rect 568326 27984 568394 28040
rect 568450 27984 568518 28040
rect 568574 27984 568642 28040
rect 568698 27984 568766 28040
rect 568822 27984 568890 28040
rect 568946 27984 569014 28040
rect 569070 27984 569138 28040
rect 569194 27984 588022 28040
rect 588078 27984 588146 28040
rect 588202 27984 588270 28040
rect 588326 27984 588394 28040
rect 588450 27984 588518 28040
rect 588574 27984 588642 28040
rect 588698 27984 588766 28040
rect 588822 27984 588890 28040
rect 588946 27984 589014 28040
rect 589070 27984 589138 28040
rect 589194 27984 597980 28040
rect -1916 27978 597980 27984
rect -1916 27922 -1820 27978
rect -1764 27922 -1696 27978
rect -1640 27922 -1572 27978
rect -1516 27922 -1448 27978
rect -1392 27922 6970 27978
rect 7026 27922 7094 27978
rect 7150 27922 7218 27978
rect 7274 27922 7342 27978
rect 7398 27922 24970 27978
rect 25026 27922 25094 27978
rect 25150 27922 25218 27978
rect 25274 27922 25342 27978
rect 25398 27922 42970 27978
rect 43026 27922 43094 27978
rect 43150 27922 43218 27978
rect 43274 27922 43342 27978
rect 43398 27922 60970 27978
rect 61026 27922 61094 27978
rect 61150 27922 61218 27978
rect 61274 27922 61342 27978
rect 61398 27922 78970 27978
rect 79026 27922 79094 27978
rect 79150 27922 79218 27978
rect 79274 27922 79342 27978
rect 79398 27922 96970 27978
rect 97026 27922 97094 27978
rect 97150 27922 97218 27978
rect 97274 27922 97342 27978
rect 97398 27922 114970 27978
rect 115026 27922 115094 27978
rect 115150 27922 115218 27978
rect 115274 27922 115342 27978
rect 115398 27922 132970 27978
rect 133026 27922 133094 27978
rect 133150 27922 133218 27978
rect 133274 27922 133342 27978
rect 133398 27922 150970 27978
rect 151026 27922 151094 27978
rect 151150 27922 151218 27978
rect 151274 27922 151342 27978
rect 151398 27922 168970 27978
rect 169026 27922 169094 27978
rect 169150 27922 169218 27978
rect 169274 27922 169342 27978
rect 169398 27922 186970 27978
rect 187026 27922 187094 27978
rect 187150 27922 187218 27978
rect 187274 27922 187342 27978
rect 187398 27922 204970 27978
rect 205026 27922 205094 27978
rect 205150 27922 205218 27978
rect 205274 27922 205342 27978
rect 205398 27922 222970 27978
rect 223026 27922 223094 27978
rect 223150 27922 223218 27978
rect 223274 27922 223342 27978
rect 223398 27922 240970 27978
rect 241026 27922 241094 27978
rect 241150 27922 241218 27978
rect 241274 27922 241342 27978
rect 241398 27922 258970 27978
rect 259026 27922 259094 27978
rect 259150 27922 259218 27978
rect 259274 27922 259342 27978
rect 259398 27922 276970 27978
rect 277026 27922 277094 27978
rect 277150 27922 277218 27978
rect 277274 27922 277342 27978
rect 277398 27922 294970 27978
rect 295026 27922 295094 27978
rect 295150 27922 295218 27978
rect 295274 27922 295342 27978
rect 295398 27922 312970 27978
rect 313026 27922 313094 27978
rect 313150 27922 313218 27978
rect 313274 27922 313342 27978
rect 313398 27922 330970 27978
rect 331026 27922 331094 27978
rect 331150 27922 331218 27978
rect 331274 27922 331342 27978
rect 331398 27922 348970 27978
rect 349026 27922 349094 27978
rect 349150 27922 349218 27978
rect 349274 27922 349342 27978
rect 349398 27922 366970 27978
rect 367026 27922 367094 27978
rect 367150 27922 367218 27978
rect 367274 27922 367342 27978
rect 367398 27922 384970 27978
rect 385026 27922 385094 27978
rect 385150 27922 385218 27978
rect 385274 27922 385342 27978
rect 385398 27922 402970 27978
rect 403026 27922 403094 27978
rect 403150 27922 403218 27978
rect 403274 27922 403342 27978
rect 403398 27922 420970 27978
rect 421026 27922 421094 27978
rect 421150 27922 421218 27978
rect 421274 27922 421342 27978
rect 421398 27922 438970 27978
rect 439026 27922 439094 27978
rect 439150 27922 439218 27978
rect 439274 27922 439342 27978
rect 439398 27922 456970 27978
rect 457026 27922 457094 27978
rect 457150 27922 457218 27978
rect 457274 27922 457342 27978
rect 457398 27922 474970 27978
rect 475026 27922 475094 27978
rect 475150 27922 475218 27978
rect 475274 27922 475342 27978
rect 475398 27922 492970 27978
rect 493026 27922 493094 27978
rect 493150 27922 493218 27978
rect 493274 27922 493342 27978
rect 493398 27922 510970 27978
rect 511026 27922 511094 27978
rect 511150 27922 511218 27978
rect 511274 27922 511342 27978
rect 511398 27922 528970 27978
rect 529026 27922 529094 27978
rect 529150 27922 529218 27978
rect 529274 27922 529342 27978
rect 529398 27922 546970 27978
rect 547026 27922 547094 27978
rect 547150 27922 547218 27978
rect 547274 27922 547342 27978
rect 547398 27922 564970 27978
rect 565026 27922 565094 27978
rect 565150 27922 565218 27978
rect 565274 27922 565342 27978
rect 565398 27922 582970 27978
rect 583026 27922 583094 27978
rect 583150 27922 583218 27978
rect 583274 27922 583342 27978
rect 583398 27922 597456 27978
rect 597512 27922 597580 27978
rect 597636 27922 597704 27978
rect 597760 27922 597828 27978
rect 597884 27922 597980 27978
rect -1916 27916 597980 27922
rect -1916 27860 568022 27916
rect 568078 27860 568146 27916
rect 568202 27860 568270 27916
rect 568326 27860 568394 27916
rect 568450 27860 568518 27916
rect 568574 27860 568642 27916
rect 568698 27860 568766 27916
rect 568822 27860 568890 27916
rect 568946 27860 569014 27916
rect 569070 27860 569138 27916
rect 569194 27860 588022 27916
rect 588078 27860 588146 27916
rect 588202 27860 588270 27916
rect 588326 27860 588394 27916
rect 588450 27860 588518 27916
rect 588574 27860 588642 27916
rect 588698 27860 588766 27916
rect 588822 27860 588890 27916
rect 588946 27860 589014 27916
rect 589070 27860 589138 27916
rect 589194 27860 597980 27916
rect -1916 27826 597980 27860
rect 112236 27658 203380 27674
rect 112236 27602 112252 27658
rect 112308 27602 203308 27658
rect 203364 27602 203380 27658
rect 112236 27586 203380 27602
rect 215836 27658 551588 27674
rect 215836 27602 215852 27658
rect 215908 27602 551516 27658
rect 551572 27602 551588 27658
rect 215836 27586 551588 27602
rect 218412 27478 551364 27494
rect 218412 27422 218428 27478
rect 218484 27422 219884 27478
rect 219940 27422 551292 27478
rect 551348 27422 551364 27478
rect 218412 27406 551364 27422
rect 110444 26938 209428 26954
rect 110444 26882 110460 26938
rect 110516 26882 209356 26938
rect 209412 26882 209428 26938
rect 110444 26866 209428 26882
rect 554412 26578 562004 26594
rect 554412 26522 554428 26578
rect 554484 26522 557116 26578
rect 557172 26522 561932 26578
rect 561988 26522 562004 26578
rect 554412 26506 562004 26522
rect 554524 26038 565700 26054
rect 554524 25982 554540 26038
rect 554596 25982 559356 26038
rect 559412 25982 565628 26038
rect 565684 25982 565700 26038
rect 554524 25966 565700 25982
rect 554524 25858 560324 25874
rect 554524 25802 554540 25858
rect 554596 25802 557564 25858
rect 557620 25802 560252 25858
rect 560308 25802 560324 25858
rect 554524 25786 560324 25802
rect 563708 25318 577124 25334
rect 563708 25262 563724 25318
rect 563780 25262 577052 25318
rect 577108 25262 577124 25318
rect 563708 25246 577124 25262
rect 350236 25138 591460 25154
rect 350236 25082 350252 25138
rect 350308 25082 591388 25138
rect 591444 25082 591460 25138
rect 350236 25066 591460 25082
rect 371292 24958 570180 24974
rect 371292 24902 371308 24958
rect 371364 24902 567756 24958
rect 567812 24902 570108 24958
rect 570164 24902 570180 24958
rect 371292 24886 570180 24902
rect 561076 24778 563684 24794
rect 561076 24722 563612 24778
rect 563668 24722 563684 24778
rect 561076 24706 563684 24722
rect 561076 24434 561164 24706
rect 383836 24418 561164 24434
rect 383836 24362 383852 24418
rect 383908 24362 557676 24418
rect 557732 24362 561164 24418
rect 383836 24346 561164 24362
rect -1916 22412 597980 22446
rect -1916 22356 558022 22412
rect 558078 22356 558146 22412
rect 558202 22356 558270 22412
rect 558326 22356 558394 22412
rect 558450 22356 558518 22412
rect 558574 22356 558642 22412
rect 558698 22356 558766 22412
rect 558822 22356 558890 22412
rect 558946 22356 559014 22412
rect 559070 22356 559138 22412
rect 559194 22356 578022 22412
rect 578078 22356 578146 22412
rect 578202 22356 578270 22412
rect 578326 22356 578394 22412
rect 578450 22356 578518 22412
rect 578574 22356 578642 22412
rect 578698 22356 578766 22412
rect 578822 22356 578890 22412
rect 578946 22356 579014 22412
rect 579070 22356 579138 22412
rect 579194 22356 597980 22412
rect -1916 22350 597980 22356
rect -1916 22294 -860 22350
rect -804 22294 -736 22350
rect -680 22294 -612 22350
rect -556 22294 -488 22350
rect -432 22294 3250 22350
rect 3306 22294 3374 22350
rect 3430 22294 3498 22350
rect 3554 22294 3622 22350
rect 3678 22294 21250 22350
rect 21306 22294 21374 22350
rect 21430 22294 21498 22350
rect 21554 22294 21622 22350
rect 21678 22294 39250 22350
rect 39306 22294 39374 22350
rect 39430 22294 39498 22350
rect 39554 22294 39622 22350
rect 39678 22294 57250 22350
rect 57306 22294 57374 22350
rect 57430 22294 57498 22350
rect 57554 22294 57622 22350
rect 57678 22294 75250 22350
rect 75306 22294 75374 22350
rect 75430 22294 75498 22350
rect 75554 22294 75622 22350
rect 75678 22294 93250 22350
rect 93306 22294 93374 22350
rect 93430 22294 93498 22350
rect 93554 22294 93622 22350
rect 93678 22294 111250 22350
rect 111306 22294 111374 22350
rect 111430 22294 111498 22350
rect 111554 22294 111622 22350
rect 111678 22294 129250 22350
rect 129306 22294 129374 22350
rect 129430 22294 129498 22350
rect 129554 22294 129622 22350
rect 129678 22294 147250 22350
rect 147306 22294 147374 22350
rect 147430 22294 147498 22350
rect 147554 22294 147622 22350
rect 147678 22294 165250 22350
rect 165306 22294 165374 22350
rect 165430 22294 165498 22350
rect 165554 22294 165622 22350
rect 165678 22294 183250 22350
rect 183306 22294 183374 22350
rect 183430 22294 183498 22350
rect 183554 22294 183622 22350
rect 183678 22294 201250 22350
rect 201306 22294 201374 22350
rect 201430 22294 201498 22350
rect 201554 22294 201622 22350
rect 201678 22294 219250 22350
rect 219306 22294 219374 22350
rect 219430 22294 219498 22350
rect 219554 22294 219622 22350
rect 219678 22294 237250 22350
rect 237306 22294 237374 22350
rect 237430 22294 237498 22350
rect 237554 22294 237622 22350
rect 237678 22294 255250 22350
rect 255306 22294 255374 22350
rect 255430 22294 255498 22350
rect 255554 22294 255622 22350
rect 255678 22294 273250 22350
rect 273306 22294 273374 22350
rect 273430 22294 273498 22350
rect 273554 22294 273622 22350
rect 273678 22294 291250 22350
rect 291306 22294 291374 22350
rect 291430 22294 291498 22350
rect 291554 22294 291622 22350
rect 291678 22294 309250 22350
rect 309306 22294 309374 22350
rect 309430 22294 309498 22350
rect 309554 22294 309622 22350
rect 309678 22294 327250 22350
rect 327306 22294 327374 22350
rect 327430 22294 327498 22350
rect 327554 22294 327622 22350
rect 327678 22294 345250 22350
rect 345306 22294 345374 22350
rect 345430 22294 345498 22350
rect 345554 22294 345622 22350
rect 345678 22294 363250 22350
rect 363306 22294 363374 22350
rect 363430 22294 363498 22350
rect 363554 22294 363622 22350
rect 363678 22294 381250 22350
rect 381306 22294 381374 22350
rect 381430 22294 381498 22350
rect 381554 22294 381622 22350
rect 381678 22294 399250 22350
rect 399306 22294 399374 22350
rect 399430 22294 399498 22350
rect 399554 22294 399622 22350
rect 399678 22294 417250 22350
rect 417306 22294 417374 22350
rect 417430 22294 417498 22350
rect 417554 22294 417622 22350
rect 417678 22294 435250 22350
rect 435306 22294 435374 22350
rect 435430 22294 435498 22350
rect 435554 22294 435622 22350
rect 435678 22294 453250 22350
rect 453306 22294 453374 22350
rect 453430 22294 453498 22350
rect 453554 22294 453622 22350
rect 453678 22294 471250 22350
rect 471306 22294 471374 22350
rect 471430 22294 471498 22350
rect 471554 22294 471622 22350
rect 471678 22294 489250 22350
rect 489306 22294 489374 22350
rect 489430 22294 489498 22350
rect 489554 22294 489622 22350
rect 489678 22294 507250 22350
rect 507306 22294 507374 22350
rect 507430 22294 507498 22350
rect 507554 22294 507622 22350
rect 507678 22294 525250 22350
rect 525306 22294 525374 22350
rect 525430 22294 525498 22350
rect 525554 22294 525622 22350
rect 525678 22294 543250 22350
rect 543306 22294 543374 22350
rect 543430 22294 543498 22350
rect 543554 22294 543622 22350
rect 543678 22294 561250 22350
rect 561306 22294 561374 22350
rect 561430 22294 561498 22350
rect 561554 22294 561622 22350
rect 561678 22294 596496 22350
rect 596552 22294 596620 22350
rect 596676 22294 596744 22350
rect 596800 22294 596868 22350
rect 596924 22294 597980 22350
rect -1916 22288 597980 22294
rect -1916 22232 558022 22288
rect 558078 22232 558146 22288
rect 558202 22232 558270 22288
rect 558326 22232 558394 22288
rect 558450 22232 558518 22288
rect 558574 22232 558642 22288
rect 558698 22232 558766 22288
rect 558822 22232 558890 22288
rect 558946 22232 559014 22288
rect 559070 22232 559138 22288
rect 559194 22232 578022 22288
rect 578078 22232 578146 22288
rect 578202 22232 578270 22288
rect 578326 22232 578394 22288
rect 578450 22232 578518 22288
rect 578574 22232 578642 22288
rect 578698 22232 578766 22288
rect 578822 22232 578890 22288
rect 578946 22232 579014 22288
rect 579070 22232 579138 22288
rect 579194 22232 597980 22288
rect -1916 22226 597980 22232
rect -1916 22170 -860 22226
rect -804 22170 -736 22226
rect -680 22170 -612 22226
rect -556 22170 -488 22226
rect -432 22170 3250 22226
rect 3306 22170 3374 22226
rect 3430 22170 3498 22226
rect 3554 22170 3622 22226
rect 3678 22170 21250 22226
rect 21306 22170 21374 22226
rect 21430 22170 21498 22226
rect 21554 22170 21622 22226
rect 21678 22170 39250 22226
rect 39306 22170 39374 22226
rect 39430 22170 39498 22226
rect 39554 22170 39622 22226
rect 39678 22170 57250 22226
rect 57306 22170 57374 22226
rect 57430 22170 57498 22226
rect 57554 22170 57622 22226
rect 57678 22170 75250 22226
rect 75306 22170 75374 22226
rect 75430 22170 75498 22226
rect 75554 22170 75622 22226
rect 75678 22170 93250 22226
rect 93306 22170 93374 22226
rect 93430 22170 93498 22226
rect 93554 22170 93622 22226
rect 93678 22170 111250 22226
rect 111306 22170 111374 22226
rect 111430 22170 111498 22226
rect 111554 22170 111622 22226
rect 111678 22170 129250 22226
rect 129306 22170 129374 22226
rect 129430 22170 129498 22226
rect 129554 22170 129622 22226
rect 129678 22170 147250 22226
rect 147306 22170 147374 22226
rect 147430 22170 147498 22226
rect 147554 22170 147622 22226
rect 147678 22170 165250 22226
rect 165306 22170 165374 22226
rect 165430 22170 165498 22226
rect 165554 22170 165622 22226
rect 165678 22170 183250 22226
rect 183306 22170 183374 22226
rect 183430 22170 183498 22226
rect 183554 22170 183622 22226
rect 183678 22170 201250 22226
rect 201306 22170 201374 22226
rect 201430 22170 201498 22226
rect 201554 22170 201622 22226
rect 201678 22170 219250 22226
rect 219306 22170 219374 22226
rect 219430 22170 219498 22226
rect 219554 22170 219622 22226
rect 219678 22170 237250 22226
rect 237306 22170 237374 22226
rect 237430 22170 237498 22226
rect 237554 22170 237622 22226
rect 237678 22170 255250 22226
rect 255306 22170 255374 22226
rect 255430 22170 255498 22226
rect 255554 22170 255622 22226
rect 255678 22170 273250 22226
rect 273306 22170 273374 22226
rect 273430 22170 273498 22226
rect 273554 22170 273622 22226
rect 273678 22170 291250 22226
rect 291306 22170 291374 22226
rect 291430 22170 291498 22226
rect 291554 22170 291622 22226
rect 291678 22170 309250 22226
rect 309306 22170 309374 22226
rect 309430 22170 309498 22226
rect 309554 22170 309622 22226
rect 309678 22170 327250 22226
rect 327306 22170 327374 22226
rect 327430 22170 327498 22226
rect 327554 22170 327622 22226
rect 327678 22170 345250 22226
rect 345306 22170 345374 22226
rect 345430 22170 345498 22226
rect 345554 22170 345622 22226
rect 345678 22170 363250 22226
rect 363306 22170 363374 22226
rect 363430 22170 363498 22226
rect 363554 22170 363622 22226
rect 363678 22170 381250 22226
rect 381306 22170 381374 22226
rect 381430 22170 381498 22226
rect 381554 22170 381622 22226
rect 381678 22170 399250 22226
rect 399306 22170 399374 22226
rect 399430 22170 399498 22226
rect 399554 22170 399622 22226
rect 399678 22170 417250 22226
rect 417306 22170 417374 22226
rect 417430 22170 417498 22226
rect 417554 22170 417622 22226
rect 417678 22170 435250 22226
rect 435306 22170 435374 22226
rect 435430 22170 435498 22226
rect 435554 22170 435622 22226
rect 435678 22170 453250 22226
rect 453306 22170 453374 22226
rect 453430 22170 453498 22226
rect 453554 22170 453622 22226
rect 453678 22170 471250 22226
rect 471306 22170 471374 22226
rect 471430 22170 471498 22226
rect 471554 22170 471622 22226
rect 471678 22170 489250 22226
rect 489306 22170 489374 22226
rect 489430 22170 489498 22226
rect 489554 22170 489622 22226
rect 489678 22170 507250 22226
rect 507306 22170 507374 22226
rect 507430 22170 507498 22226
rect 507554 22170 507622 22226
rect 507678 22170 525250 22226
rect 525306 22170 525374 22226
rect 525430 22170 525498 22226
rect 525554 22170 525622 22226
rect 525678 22170 543250 22226
rect 543306 22170 543374 22226
rect 543430 22170 543498 22226
rect 543554 22170 543622 22226
rect 543678 22170 561250 22226
rect 561306 22170 561374 22226
rect 561430 22170 561498 22226
rect 561554 22170 561622 22226
rect 561678 22170 596496 22226
rect 596552 22170 596620 22226
rect 596676 22170 596744 22226
rect 596800 22170 596868 22226
rect 596924 22170 597980 22226
rect -1916 22164 597980 22170
rect -1916 22108 558022 22164
rect 558078 22108 558146 22164
rect 558202 22108 558270 22164
rect 558326 22108 558394 22164
rect 558450 22108 558518 22164
rect 558574 22108 558642 22164
rect 558698 22108 558766 22164
rect 558822 22108 558890 22164
rect 558946 22108 559014 22164
rect 559070 22108 559138 22164
rect 559194 22108 578022 22164
rect 578078 22108 578146 22164
rect 578202 22108 578270 22164
rect 578326 22108 578394 22164
rect 578450 22108 578518 22164
rect 578574 22108 578642 22164
rect 578698 22108 578766 22164
rect 578822 22108 578890 22164
rect 578946 22108 579014 22164
rect 579070 22108 579138 22164
rect 579194 22108 597980 22164
rect -1916 22102 597980 22108
rect -1916 22046 -860 22102
rect -804 22046 -736 22102
rect -680 22046 -612 22102
rect -556 22046 -488 22102
rect -432 22046 3250 22102
rect 3306 22046 3374 22102
rect 3430 22046 3498 22102
rect 3554 22046 3622 22102
rect 3678 22046 21250 22102
rect 21306 22046 21374 22102
rect 21430 22046 21498 22102
rect 21554 22046 21622 22102
rect 21678 22046 39250 22102
rect 39306 22046 39374 22102
rect 39430 22046 39498 22102
rect 39554 22046 39622 22102
rect 39678 22046 57250 22102
rect 57306 22046 57374 22102
rect 57430 22046 57498 22102
rect 57554 22046 57622 22102
rect 57678 22046 75250 22102
rect 75306 22046 75374 22102
rect 75430 22046 75498 22102
rect 75554 22046 75622 22102
rect 75678 22046 93250 22102
rect 93306 22046 93374 22102
rect 93430 22046 93498 22102
rect 93554 22046 93622 22102
rect 93678 22046 111250 22102
rect 111306 22046 111374 22102
rect 111430 22046 111498 22102
rect 111554 22046 111622 22102
rect 111678 22046 129250 22102
rect 129306 22046 129374 22102
rect 129430 22046 129498 22102
rect 129554 22046 129622 22102
rect 129678 22046 147250 22102
rect 147306 22046 147374 22102
rect 147430 22046 147498 22102
rect 147554 22046 147622 22102
rect 147678 22046 165250 22102
rect 165306 22046 165374 22102
rect 165430 22046 165498 22102
rect 165554 22046 165622 22102
rect 165678 22046 183250 22102
rect 183306 22046 183374 22102
rect 183430 22046 183498 22102
rect 183554 22046 183622 22102
rect 183678 22046 201250 22102
rect 201306 22046 201374 22102
rect 201430 22046 201498 22102
rect 201554 22046 201622 22102
rect 201678 22046 219250 22102
rect 219306 22046 219374 22102
rect 219430 22046 219498 22102
rect 219554 22046 219622 22102
rect 219678 22046 237250 22102
rect 237306 22046 237374 22102
rect 237430 22046 237498 22102
rect 237554 22046 237622 22102
rect 237678 22046 255250 22102
rect 255306 22046 255374 22102
rect 255430 22046 255498 22102
rect 255554 22046 255622 22102
rect 255678 22046 273250 22102
rect 273306 22046 273374 22102
rect 273430 22046 273498 22102
rect 273554 22046 273622 22102
rect 273678 22046 291250 22102
rect 291306 22046 291374 22102
rect 291430 22046 291498 22102
rect 291554 22046 291622 22102
rect 291678 22046 309250 22102
rect 309306 22046 309374 22102
rect 309430 22046 309498 22102
rect 309554 22046 309622 22102
rect 309678 22046 327250 22102
rect 327306 22046 327374 22102
rect 327430 22046 327498 22102
rect 327554 22046 327622 22102
rect 327678 22046 345250 22102
rect 345306 22046 345374 22102
rect 345430 22046 345498 22102
rect 345554 22046 345622 22102
rect 345678 22046 363250 22102
rect 363306 22046 363374 22102
rect 363430 22046 363498 22102
rect 363554 22046 363622 22102
rect 363678 22046 381250 22102
rect 381306 22046 381374 22102
rect 381430 22046 381498 22102
rect 381554 22046 381622 22102
rect 381678 22046 399250 22102
rect 399306 22046 399374 22102
rect 399430 22046 399498 22102
rect 399554 22046 399622 22102
rect 399678 22046 417250 22102
rect 417306 22046 417374 22102
rect 417430 22046 417498 22102
rect 417554 22046 417622 22102
rect 417678 22046 435250 22102
rect 435306 22046 435374 22102
rect 435430 22046 435498 22102
rect 435554 22046 435622 22102
rect 435678 22046 453250 22102
rect 453306 22046 453374 22102
rect 453430 22046 453498 22102
rect 453554 22046 453622 22102
rect 453678 22046 471250 22102
rect 471306 22046 471374 22102
rect 471430 22046 471498 22102
rect 471554 22046 471622 22102
rect 471678 22046 489250 22102
rect 489306 22046 489374 22102
rect 489430 22046 489498 22102
rect 489554 22046 489622 22102
rect 489678 22046 507250 22102
rect 507306 22046 507374 22102
rect 507430 22046 507498 22102
rect 507554 22046 507622 22102
rect 507678 22046 525250 22102
rect 525306 22046 525374 22102
rect 525430 22046 525498 22102
rect 525554 22046 525622 22102
rect 525678 22046 543250 22102
rect 543306 22046 543374 22102
rect 543430 22046 543498 22102
rect 543554 22046 543622 22102
rect 543678 22046 561250 22102
rect 561306 22046 561374 22102
rect 561430 22046 561498 22102
rect 561554 22046 561622 22102
rect 561678 22046 596496 22102
rect 596552 22046 596620 22102
rect 596676 22046 596744 22102
rect 596800 22046 596868 22102
rect 596924 22046 597980 22102
rect -1916 22040 597980 22046
rect -1916 21984 558022 22040
rect 558078 21984 558146 22040
rect 558202 21984 558270 22040
rect 558326 21984 558394 22040
rect 558450 21984 558518 22040
rect 558574 21984 558642 22040
rect 558698 21984 558766 22040
rect 558822 21984 558890 22040
rect 558946 21984 559014 22040
rect 559070 21984 559138 22040
rect 559194 21984 578022 22040
rect 578078 21984 578146 22040
rect 578202 21984 578270 22040
rect 578326 21984 578394 22040
rect 578450 21984 578518 22040
rect 578574 21984 578642 22040
rect 578698 21984 578766 22040
rect 578822 21984 578890 22040
rect 578946 21984 579014 22040
rect 579070 21984 579138 22040
rect 579194 21984 597980 22040
rect -1916 21978 597980 21984
rect -1916 21922 -860 21978
rect -804 21922 -736 21978
rect -680 21922 -612 21978
rect -556 21922 -488 21978
rect -432 21922 3250 21978
rect 3306 21922 3374 21978
rect 3430 21922 3498 21978
rect 3554 21922 3622 21978
rect 3678 21922 21250 21978
rect 21306 21922 21374 21978
rect 21430 21922 21498 21978
rect 21554 21922 21622 21978
rect 21678 21922 39250 21978
rect 39306 21922 39374 21978
rect 39430 21922 39498 21978
rect 39554 21922 39622 21978
rect 39678 21922 57250 21978
rect 57306 21922 57374 21978
rect 57430 21922 57498 21978
rect 57554 21922 57622 21978
rect 57678 21922 75250 21978
rect 75306 21922 75374 21978
rect 75430 21922 75498 21978
rect 75554 21922 75622 21978
rect 75678 21922 93250 21978
rect 93306 21922 93374 21978
rect 93430 21922 93498 21978
rect 93554 21922 93622 21978
rect 93678 21922 111250 21978
rect 111306 21922 111374 21978
rect 111430 21922 111498 21978
rect 111554 21922 111622 21978
rect 111678 21922 129250 21978
rect 129306 21922 129374 21978
rect 129430 21922 129498 21978
rect 129554 21922 129622 21978
rect 129678 21922 147250 21978
rect 147306 21922 147374 21978
rect 147430 21922 147498 21978
rect 147554 21922 147622 21978
rect 147678 21922 165250 21978
rect 165306 21922 165374 21978
rect 165430 21922 165498 21978
rect 165554 21922 165622 21978
rect 165678 21922 183250 21978
rect 183306 21922 183374 21978
rect 183430 21922 183498 21978
rect 183554 21922 183622 21978
rect 183678 21922 201250 21978
rect 201306 21922 201374 21978
rect 201430 21922 201498 21978
rect 201554 21922 201622 21978
rect 201678 21922 219250 21978
rect 219306 21922 219374 21978
rect 219430 21922 219498 21978
rect 219554 21922 219622 21978
rect 219678 21922 237250 21978
rect 237306 21922 237374 21978
rect 237430 21922 237498 21978
rect 237554 21922 237622 21978
rect 237678 21922 255250 21978
rect 255306 21922 255374 21978
rect 255430 21922 255498 21978
rect 255554 21922 255622 21978
rect 255678 21922 273250 21978
rect 273306 21922 273374 21978
rect 273430 21922 273498 21978
rect 273554 21922 273622 21978
rect 273678 21922 291250 21978
rect 291306 21922 291374 21978
rect 291430 21922 291498 21978
rect 291554 21922 291622 21978
rect 291678 21922 309250 21978
rect 309306 21922 309374 21978
rect 309430 21922 309498 21978
rect 309554 21922 309622 21978
rect 309678 21922 327250 21978
rect 327306 21922 327374 21978
rect 327430 21922 327498 21978
rect 327554 21922 327622 21978
rect 327678 21922 345250 21978
rect 345306 21922 345374 21978
rect 345430 21922 345498 21978
rect 345554 21922 345622 21978
rect 345678 21922 363250 21978
rect 363306 21922 363374 21978
rect 363430 21922 363498 21978
rect 363554 21922 363622 21978
rect 363678 21922 381250 21978
rect 381306 21922 381374 21978
rect 381430 21922 381498 21978
rect 381554 21922 381622 21978
rect 381678 21922 399250 21978
rect 399306 21922 399374 21978
rect 399430 21922 399498 21978
rect 399554 21922 399622 21978
rect 399678 21922 417250 21978
rect 417306 21922 417374 21978
rect 417430 21922 417498 21978
rect 417554 21922 417622 21978
rect 417678 21922 435250 21978
rect 435306 21922 435374 21978
rect 435430 21922 435498 21978
rect 435554 21922 435622 21978
rect 435678 21922 453250 21978
rect 453306 21922 453374 21978
rect 453430 21922 453498 21978
rect 453554 21922 453622 21978
rect 453678 21922 471250 21978
rect 471306 21922 471374 21978
rect 471430 21922 471498 21978
rect 471554 21922 471622 21978
rect 471678 21922 489250 21978
rect 489306 21922 489374 21978
rect 489430 21922 489498 21978
rect 489554 21922 489622 21978
rect 489678 21922 507250 21978
rect 507306 21922 507374 21978
rect 507430 21922 507498 21978
rect 507554 21922 507622 21978
rect 507678 21922 525250 21978
rect 525306 21922 525374 21978
rect 525430 21922 525498 21978
rect 525554 21922 525622 21978
rect 525678 21922 543250 21978
rect 543306 21922 543374 21978
rect 543430 21922 543498 21978
rect 543554 21922 543622 21978
rect 543678 21922 561250 21978
rect 561306 21922 561374 21978
rect 561430 21922 561498 21978
rect 561554 21922 561622 21978
rect 561678 21922 596496 21978
rect 596552 21922 596620 21978
rect 596676 21922 596744 21978
rect 596800 21922 596868 21978
rect 596924 21922 597980 21978
rect -1916 21916 597980 21922
rect -1916 21860 558022 21916
rect 558078 21860 558146 21916
rect 558202 21860 558270 21916
rect 558326 21860 558394 21916
rect 558450 21860 558518 21916
rect 558574 21860 558642 21916
rect 558698 21860 558766 21916
rect 558822 21860 558890 21916
rect 558946 21860 559014 21916
rect 559070 21860 559138 21916
rect 559194 21860 578022 21916
rect 578078 21860 578146 21916
rect 578202 21860 578270 21916
rect 578326 21860 578394 21916
rect 578450 21860 578518 21916
rect 578574 21860 578642 21916
rect 578698 21860 578766 21916
rect 578822 21860 578890 21916
rect 578946 21860 579014 21916
rect 579070 21860 579138 21916
rect 579194 21860 597980 21916
rect -1916 21826 597980 21860
rect 73820 20098 563796 20114
rect 73820 20042 73836 20098
rect 73892 20042 563724 20098
rect 563780 20042 563796 20098
rect 73820 20026 563796 20042
rect 557212 13078 560100 13094
rect 557212 13022 557228 13078
rect 557284 13022 560028 13078
rect 560084 13022 560100 13078
rect 557212 13006 560100 13022
rect 551052 11638 552708 11654
rect 551052 11582 551068 11638
rect 551124 11582 552636 11638
rect 552692 11582 552708 11638
rect 551052 11566 552708 11582
rect 552620 10738 586084 10754
rect 552620 10682 552636 10738
rect 552692 10682 586012 10738
rect 586068 10682 586084 10738
rect 552620 10666 586084 10682
rect -1916 10350 597980 10446
rect -1916 10294 -1820 10350
rect -1764 10294 -1696 10350
rect -1640 10294 -1572 10350
rect -1516 10294 -1448 10350
rect -1392 10294 6970 10350
rect 7026 10294 7094 10350
rect 7150 10294 7218 10350
rect 7274 10294 7342 10350
rect 7398 10294 24970 10350
rect 25026 10294 25094 10350
rect 25150 10294 25218 10350
rect 25274 10294 25342 10350
rect 25398 10294 42970 10350
rect 43026 10294 43094 10350
rect 43150 10294 43218 10350
rect 43274 10294 43342 10350
rect 43398 10294 60970 10350
rect 61026 10294 61094 10350
rect 61150 10294 61218 10350
rect 61274 10294 61342 10350
rect 61398 10294 78970 10350
rect 79026 10294 79094 10350
rect 79150 10294 79218 10350
rect 79274 10294 79342 10350
rect 79398 10294 96970 10350
rect 97026 10294 97094 10350
rect 97150 10294 97218 10350
rect 97274 10294 97342 10350
rect 97398 10294 114970 10350
rect 115026 10294 115094 10350
rect 115150 10294 115218 10350
rect 115274 10294 115342 10350
rect 115398 10294 132970 10350
rect 133026 10294 133094 10350
rect 133150 10294 133218 10350
rect 133274 10294 133342 10350
rect 133398 10294 150970 10350
rect 151026 10294 151094 10350
rect 151150 10294 151218 10350
rect 151274 10294 151342 10350
rect 151398 10294 168970 10350
rect 169026 10294 169094 10350
rect 169150 10294 169218 10350
rect 169274 10294 169342 10350
rect 169398 10294 186970 10350
rect 187026 10294 187094 10350
rect 187150 10294 187218 10350
rect 187274 10294 187342 10350
rect 187398 10294 204970 10350
rect 205026 10294 205094 10350
rect 205150 10294 205218 10350
rect 205274 10294 205342 10350
rect 205398 10294 222970 10350
rect 223026 10294 223094 10350
rect 223150 10294 223218 10350
rect 223274 10294 223342 10350
rect 223398 10294 240970 10350
rect 241026 10294 241094 10350
rect 241150 10294 241218 10350
rect 241274 10294 241342 10350
rect 241398 10294 258970 10350
rect 259026 10294 259094 10350
rect 259150 10294 259218 10350
rect 259274 10294 259342 10350
rect 259398 10294 276970 10350
rect 277026 10294 277094 10350
rect 277150 10294 277218 10350
rect 277274 10294 277342 10350
rect 277398 10294 294970 10350
rect 295026 10294 295094 10350
rect 295150 10294 295218 10350
rect 295274 10294 295342 10350
rect 295398 10294 312970 10350
rect 313026 10294 313094 10350
rect 313150 10294 313218 10350
rect 313274 10294 313342 10350
rect 313398 10294 330970 10350
rect 331026 10294 331094 10350
rect 331150 10294 331218 10350
rect 331274 10294 331342 10350
rect 331398 10294 348970 10350
rect 349026 10294 349094 10350
rect 349150 10294 349218 10350
rect 349274 10294 349342 10350
rect 349398 10294 366970 10350
rect 367026 10294 367094 10350
rect 367150 10294 367218 10350
rect 367274 10294 367342 10350
rect 367398 10294 384970 10350
rect 385026 10294 385094 10350
rect 385150 10294 385218 10350
rect 385274 10294 385342 10350
rect 385398 10294 402970 10350
rect 403026 10294 403094 10350
rect 403150 10294 403218 10350
rect 403274 10294 403342 10350
rect 403398 10294 420970 10350
rect 421026 10294 421094 10350
rect 421150 10294 421218 10350
rect 421274 10294 421342 10350
rect 421398 10294 438970 10350
rect 439026 10294 439094 10350
rect 439150 10294 439218 10350
rect 439274 10294 439342 10350
rect 439398 10294 456970 10350
rect 457026 10294 457094 10350
rect 457150 10294 457218 10350
rect 457274 10294 457342 10350
rect 457398 10294 474970 10350
rect 475026 10294 475094 10350
rect 475150 10294 475218 10350
rect 475274 10294 475342 10350
rect 475398 10294 492970 10350
rect 493026 10294 493094 10350
rect 493150 10294 493218 10350
rect 493274 10294 493342 10350
rect 493398 10294 510970 10350
rect 511026 10294 511094 10350
rect 511150 10294 511218 10350
rect 511274 10294 511342 10350
rect 511398 10294 528970 10350
rect 529026 10294 529094 10350
rect 529150 10294 529218 10350
rect 529274 10294 529342 10350
rect 529398 10294 546970 10350
rect 547026 10294 547094 10350
rect 547150 10294 547218 10350
rect 547274 10294 547342 10350
rect 547398 10294 564970 10350
rect 565026 10294 565094 10350
rect 565150 10294 565218 10350
rect 565274 10294 565342 10350
rect 565398 10294 582970 10350
rect 583026 10294 583094 10350
rect 583150 10294 583218 10350
rect 583274 10294 583342 10350
rect 583398 10294 597456 10350
rect 597512 10294 597580 10350
rect 597636 10294 597704 10350
rect 597760 10294 597828 10350
rect 597884 10294 597980 10350
rect -1916 10226 597980 10294
rect -1916 10170 -1820 10226
rect -1764 10170 -1696 10226
rect -1640 10170 -1572 10226
rect -1516 10170 -1448 10226
rect -1392 10170 6970 10226
rect 7026 10170 7094 10226
rect 7150 10170 7218 10226
rect 7274 10170 7342 10226
rect 7398 10170 24970 10226
rect 25026 10170 25094 10226
rect 25150 10170 25218 10226
rect 25274 10170 25342 10226
rect 25398 10170 42970 10226
rect 43026 10170 43094 10226
rect 43150 10170 43218 10226
rect 43274 10170 43342 10226
rect 43398 10170 60970 10226
rect 61026 10170 61094 10226
rect 61150 10170 61218 10226
rect 61274 10170 61342 10226
rect 61398 10170 78970 10226
rect 79026 10170 79094 10226
rect 79150 10170 79218 10226
rect 79274 10170 79342 10226
rect 79398 10170 96970 10226
rect 97026 10170 97094 10226
rect 97150 10170 97218 10226
rect 97274 10170 97342 10226
rect 97398 10170 114970 10226
rect 115026 10170 115094 10226
rect 115150 10170 115218 10226
rect 115274 10170 115342 10226
rect 115398 10170 132970 10226
rect 133026 10170 133094 10226
rect 133150 10170 133218 10226
rect 133274 10170 133342 10226
rect 133398 10170 150970 10226
rect 151026 10170 151094 10226
rect 151150 10170 151218 10226
rect 151274 10170 151342 10226
rect 151398 10170 168970 10226
rect 169026 10170 169094 10226
rect 169150 10170 169218 10226
rect 169274 10170 169342 10226
rect 169398 10170 186970 10226
rect 187026 10170 187094 10226
rect 187150 10170 187218 10226
rect 187274 10170 187342 10226
rect 187398 10170 204970 10226
rect 205026 10170 205094 10226
rect 205150 10170 205218 10226
rect 205274 10170 205342 10226
rect 205398 10170 222970 10226
rect 223026 10170 223094 10226
rect 223150 10170 223218 10226
rect 223274 10170 223342 10226
rect 223398 10170 240970 10226
rect 241026 10170 241094 10226
rect 241150 10170 241218 10226
rect 241274 10170 241342 10226
rect 241398 10170 258970 10226
rect 259026 10170 259094 10226
rect 259150 10170 259218 10226
rect 259274 10170 259342 10226
rect 259398 10170 276970 10226
rect 277026 10170 277094 10226
rect 277150 10170 277218 10226
rect 277274 10170 277342 10226
rect 277398 10170 294970 10226
rect 295026 10170 295094 10226
rect 295150 10170 295218 10226
rect 295274 10170 295342 10226
rect 295398 10170 312970 10226
rect 313026 10170 313094 10226
rect 313150 10170 313218 10226
rect 313274 10170 313342 10226
rect 313398 10170 330970 10226
rect 331026 10170 331094 10226
rect 331150 10170 331218 10226
rect 331274 10170 331342 10226
rect 331398 10170 348970 10226
rect 349026 10170 349094 10226
rect 349150 10170 349218 10226
rect 349274 10170 349342 10226
rect 349398 10170 366970 10226
rect 367026 10170 367094 10226
rect 367150 10170 367218 10226
rect 367274 10170 367342 10226
rect 367398 10170 384970 10226
rect 385026 10170 385094 10226
rect 385150 10170 385218 10226
rect 385274 10170 385342 10226
rect 385398 10170 402970 10226
rect 403026 10170 403094 10226
rect 403150 10170 403218 10226
rect 403274 10170 403342 10226
rect 403398 10170 420970 10226
rect 421026 10170 421094 10226
rect 421150 10170 421218 10226
rect 421274 10170 421342 10226
rect 421398 10170 438970 10226
rect 439026 10170 439094 10226
rect 439150 10170 439218 10226
rect 439274 10170 439342 10226
rect 439398 10170 456970 10226
rect 457026 10170 457094 10226
rect 457150 10170 457218 10226
rect 457274 10170 457342 10226
rect 457398 10170 474970 10226
rect 475026 10170 475094 10226
rect 475150 10170 475218 10226
rect 475274 10170 475342 10226
rect 475398 10170 492970 10226
rect 493026 10170 493094 10226
rect 493150 10170 493218 10226
rect 493274 10170 493342 10226
rect 493398 10170 510970 10226
rect 511026 10170 511094 10226
rect 511150 10170 511218 10226
rect 511274 10170 511342 10226
rect 511398 10170 528970 10226
rect 529026 10170 529094 10226
rect 529150 10170 529218 10226
rect 529274 10170 529342 10226
rect 529398 10170 546970 10226
rect 547026 10170 547094 10226
rect 547150 10170 547218 10226
rect 547274 10170 547342 10226
rect 547398 10170 564970 10226
rect 565026 10170 565094 10226
rect 565150 10170 565218 10226
rect 565274 10170 565342 10226
rect 565398 10170 582970 10226
rect 583026 10170 583094 10226
rect 583150 10170 583218 10226
rect 583274 10170 583342 10226
rect 583398 10170 597456 10226
rect 597512 10170 597580 10226
rect 597636 10170 597704 10226
rect 597760 10170 597828 10226
rect 597884 10170 597980 10226
rect -1916 10102 597980 10170
rect -1916 10046 -1820 10102
rect -1764 10046 -1696 10102
rect -1640 10046 -1572 10102
rect -1516 10046 -1448 10102
rect -1392 10046 6970 10102
rect 7026 10046 7094 10102
rect 7150 10046 7218 10102
rect 7274 10046 7342 10102
rect 7398 10046 24970 10102
rect 25026 10046 25094 10102
rect 25150 10046 25218 10102
rect 25274 10046 25342 10102
rect 25398 10046 42970 10102
rect 43026 10046 43094 10102
rect 43150 10046 43218 10102
rect 43274 10046 43342 10102
rect 43398 10046 60970 10102
rect 61026 10046 61094 10102
rect 61150 10046 61218 10102
rect 61274 10046 61342 10102
rect 61398 10046 78970 10102
rect 79026 10046 79094 10102
rect 79150 10046 79218 10102
rect 79274 10046 79342 10102
rect 79398 10046 96970 10102
rect 97026 10046 97094 10102
rect 97150 10046 97218 10102
rect 97274 10046 97342 10102
rect 97398 10046 114970 10102
rect 115026 10046 115094 10102
rect 115150 10046 115218 10102
rect 115274 10046 115342 10102
rect 115398 10046 132970 10102
rect 133026 10046 133094 10102
rect 133150 10046 133218 10102
rect 133274 10046 133342 10102
rect 133398 10046 150970 10102
rect 151026 10046 151094 10102
rect 151150 10046 151218 10102
rect 151274 10046 151342 10102
rect 151398 10046 168970 10102
rect 169026 10046 169094 10102
rect 169150 10046 169218 10102
rect 169274 10046 169342 10102
rect 169398 10046 186970 10102
rect 187026 10046 187094 10102
rect 187150 10046 187218 10102
rect 187274 10046 187342 10102
rect 187398 10046 204970 10102
rect 205026 10046 205094 10102
rect 205150 10046 205218 10102
rect 205274 10046 205342 10102
rect 205398 10046 222970 10102
rect 223026 10046 223094 10102
rect 223150 10046 223218 10102
rect 223274 10046 223342 10102
rect 223398 10046 240970 10102
rect 241026 10046 241094 10102
rect 241150 10046 241218 10102
rect 241274 10046 241342 10102
rect 241398 10046 258970 10102
rect 259026 10046 259094 10102
rect 259150 10046 259218 10102
rect 259274 10046 259342 10102
rect 259398 10046 276970 10102
rect 277026 10046 277094 10102
rect 277150 10046 277218 10102
rect 277274 10046 277342 10102
rect 277398 10046 294970 10102
rect 295026 10046 295094 10102
rect 295150 10046 295218 10102
rect 295274 10046 295342 10102
rect 295398 10046 312970 10102
rect 313026 10046 313094 10102
rect 313150 10046 313218 10102
rect 313274 10046 313342 10102
rect 313398 10046 330970 10102
rect 331026 10046 331094 10102
rect 331150 10046 331218 10102
rect 331274 10046 331342 10102
rect 331398 10046 348970 10102
rect 349026 10046 349094 10102
rect 349150 10046 349218 10102
rect 349274 10046 349342 10102
rect 349398 10046 366970 10102
rect 367026 10046 367094 10102
rect 367150 10046 367218 10102
rect 367274 10046 367342 10102
rect 367398 10046 384970 10102
rect 385026 10046 385094 10102
rect 385150 10046 385218 10102
rect 385274 10046 385342 10102
rect 385398 10046 402970 10102
rect 403026 10046 403094 10102
rect 403150 10046 403218 10102
rect 403274 10046 403342 10102
rect 403398 10046 420970 10102
rect 421026 10046 421094 10102
rect 421150 10046 421218 10102
rect 421274 10046 421342 10102
rect 421398 10046 438970 10102
rect 439026 10046 439094 10102
rect 439150 10046 439218 10102
rect 439274 10046 439342 10102
rect 439398 10046 456970 10102
rect 457026 10046 457094 10102
rect 457150 10046 457218 10102
rect 457274 10046 457342 10102
rect 457398 10046 474970 10102
rect 475026 10046 475094 10102
rect 475150 10046 475218 10102
rect 475274 10046 475342 10102
rect 475398 10046 492970 10102
rect 493026 10046 493094 10102
rect 493150 10046 493218 10102
rect 493274 10046 493342 10102
rect 493398 10046 510970 10102
rect 511026 10046 511094 10102
rect 511150 10046 511218 10102
rect 511274 10046 511342 10102
rect 511398 10046 528970 10102
rect 529026 10046 529094 10102
rect 529150 10046 529218 10102
rect 529274 10046 529342 10102
rect 529398 10046 546970 10102
rect 547026 10046 547094 10102
rect 547150 10046 547218 10102
rect 547274 10046 547342 10102
rect 547398 10046 564970 10102
rect 565026 10046 565094 10102
rect 565150 10046 565218 10102
rect 565274 10046 565342 10102
rect 565398 10046 582970 10102
rect 583026 10046 583094 10102
rect 583150 10046 583218 10102
rect 583274 10046 583342 10102
rect 583398 10046 597456 10102
rect 597512 10046 597580 10102
rect 597636 10046 597704 10102
rect 597760 10046 597828 10102
rect 597884 10046 597980 10102
rect -1916 9978 597980 10046
rect -1916 9922 -1820 9978
rect -1764 9922 -1696 9978
rect -1640 9922 -1572 9978
rect -1516 9922 -1448 9978
rect -1392 9922 6970 9978
rect 7026 9922 7094 9978
rect 7150 9922 7218 9978
rect 7274 9922 7342 9978
rect 7398 9922 24970 9978
rect 25026 9922 25094 9978
rect 25150 9922 25218 9978
rect 25274 9922 25342 9978
rect 25398 9922 42970 9978
rect 43026 9922 43094 9978
rect 43150 9922 43218 9978
rect 43274 9922 43342 9978
rect 43398 9922 60970 9978
rect 61026 9922 61094 9978
rect 61150 9922 61218 9978
rect 61274 9922 61342 9978
rect 61398 9922 78970 9978
rect 79026 9922 79094 9978
rect 79150 9922 79218 9978
rect 79274 9922 79342 9978
rect 79398 9922 96970 9978
rect 97026 9922 97094 9978
rect 97150 9922 97218 9978
rect 97274 9922 97342 9978
rect 97398 9922 114970 9978
rect 115026 9922 115094 9978
rect 115150 9922 115218 9978
rect 115274 9922 115342 9978
rect 115398 9922 132970 9978
rect 133026 9922 133094 9978
rect 133150 9922 133218 9978
rect 133274 9922 133342 9978
rect 133398 9922 150970 9978
rect 151026 9922 151094 9978
rect 151150 9922 151218 9978
rect 151274 9922 151342 9978
rect 151398 9922 168970 9978
rect 169026 9922 169094 9978
rect 169150 9922 169218 9978
rect 169274 9922 169342 9978
rect 169398 9922 186970 9978
rect 187026 9922 187094 9978
rect 187150 9922 187218 9978
rect 187274 9922 187342 9978
rect 187398 9922 204970 9978
rect 205026 9922 205094 9978
rect 205150 9922 205218 9978
rect 205274 9922 205342 9978
rect 205398 9922 222970 9978
rect 223026 9922 223094 9978
rect 223150 9922 223218 9978
rect 223274 9922 223342 9978
rect 223398 9922 240970 9978
rect 241026 9922 241094 9978
rect 241150 9922 241218 9978
rect 241274 9922 241342 9978
rect 241398 9922 258970 9978
rect 259026 9922 259094 9978
rect 259150 9922 259218 9978
rect 259274 9922 259342 9978
rect 259398 9922 276970 9978
rect 277026 9922 277094 9978
rect 277150 9922 277218 9978
rect 277274 9922 277342 9978
rect 277398 9922 294970 9978
rect 295026 9922 295094 9978
rect 295150 9922 295218 9978
rect 295274 9922 295342 9978
rect 295398 9922 312970 9978
rect 313026 9922 313094 9978
rect 313150 9922 313218 9978
rect 313274 9922 313342 9978
rect 313398 9922 330970 9978
rect 331026 9922 331094 9978
rect 331150 9922 331218 9978
rect 331274 9922 331342 9978
rect 331398 9922 348970 9978
rect 349026 9922 349094 9978
rect 349150 9922 349218 9978
rect 349274 9922 349342 9978
rect 349398 9922 366970 9978
rect 367026 9922 367094 9978
rect 367150 9922 367218 9978
rect 367274 9922 367342 9978
rect 367398 9922 384970 9978
rect 385026 9922 385094 9978
rect 385150 9922 385218 9978
rect 385274 9922 385342 9978
rect 385398 9922 402970 9978
rect 403026 9922 403094 9978
rect 403150 9922 403218 9978
rect 403274 9922 403342 9978
rect 403398 9922 420970 9978
rect 421026 9922 421094 9978
rect 421150 9922 421218 9978
rect 421274 9922 421342 9978
rect 421398 9922 438970 9978
rect 439026 9922 439094 9978
rect 439150 9922 439218 9978
rect 439274 9922 439342 9978
rect 439398 9922 456970 9978
rect 457026 9922 457094 9978
rect 457150 9922 457218 9978
rect 457274 9922 457342 9978
rect 457398 9922 474970 9978
rect 475026 9922 475094 9978
rect 475150 9922 475218 9978
rect 475274 9922 475342 9978
rect 475398 9922 492970 9978
rect 493026 9922 493094 9978
rect 493150 9922 493218 9978
rect 493274 9922 493342 9978
rect 493398 9922 510970 9978
rect 511026 9922 511094 9978
rect 511150 9922 511218 9978
rect 511274 9922 511342 9978
rect 511398 9922 528970 9978
rect 529026 9922 529094 9978
rect 529150 9922 529218 9978
rect 529274 9922 529342 9978
rect 529398 9922 546970 9978
rect 547026 9922 547094 9978
rect 547150 9922 547218 9978
rect 547274 9922 547342 9978
rect 547398 9922 564970 9978
rect 565026 9922 565094 9978
rect 565150 9922 565218 9978
rect 565274 9922 565342 9978
rect 565398 9922 582970 9978
rect 583026 9922 583094 9978
rect 583150 9922 583218 9978
rect 583274 9922 583342 9978
rect 583398 9922 597456 9978
rect 597512 9922 597580 9978
rect 597636 9922 597704 9978
rect 597760 9922 597828 9978
rect 597884 9922 597980 9978
rect -1916 9826 597980 9922
rect 572780 8038 577124 8054
rect 572780 7982 572796 8038
rect 572852 7982 577052 8038
rect 577108 7982 577124 8038
rect 572780 7966 577124 7982
rect 572556 7858 578020 7874
rect 572556 7802 572572 7858
rect 572628 7802 577948 7858
rect 578004 7802 578020 7858
rect 572556 7786 578020 7802
rect 572668 7678 578916 7694
rect 572668 7622 572684 7678
rect 572740 7622 578844 7678
rect 578900 7622 578916 7678
rect 572668 7606 578916 7622
rect 570988 7498 579924 7514
rect 570988 7442 571004 7498
rect 571060 7442 579852 7498
rect 579908 7442 579924 7498
rect 570988 7426 579924 7442
rect -1916 4350 597980 4446
rect -1916 4294 -860 4350
rect -804 4294 -736 4350
rect -680 4294 -612 4350
rect -556 4294 -488 4350
rect -432 4294 3250 4350
rect 3306 4294 3374 4350
rect 3430 4294 3498 4350
rect 3554 4294 3622 4350
rect 3678 4294 21250 4350
rect 21306 4294 21374 4350
rect 21430 4294 21498 4350
rect 21554 4294 21622 4350
rect 21678 4294 39250 4350
rect 39306 4294 39374 4350
rect 39430 4294 39498 4350
rect 39554 4294 39622 4350
rect 39678 4294 57250 4350
rect 57306 4294 57374 4350
rect 57430 4294 57498 4350
rect 57554 4294 57622 4350
rect 57678 4294 75250 4350
rect 75306 4294 75374 4350
rect 75430 4294 75498 4350
rect 75554 4294 75622 4350
rect 75678 4294 93250 4350
rect 93306 4294 93374 4350
rect 93430 4294 93498 4350
rect 93554 4294 93622 4350
rect 93678 4294 111250 4350
rect 111306 4294 111374 4350
rect 111430 4294 111498 4350
rect 111554 4294 111622 4350
rect 111678 4294 129250 4350
rect 129306 4294 129374 4350
rect 129430 4294 129498 4350
rect 129554 4294 129622 4350
rect 129678 4294 147250 4350
rect 147306 4294 147374 4350
rect 147430 4294 147498 4350
rect 147554 4294 147622 4350
rect 147678 4294 165250 4350
rect 165306 4294 165374 4350
rect 165430 4294 165498 4350
rect 165554 4294 165622 4350
rect 165678 4294 183250 4350
rect 183306 4294 183374 4350
rect 183430 4294 183498 4350
rect 183554 4294 183622 4350
rect 183678 4294 201250 4350
rect 201306 4294 201374 4350
rect 201430 4294 201498 4350
rect 201554 4294 201622 4350
rect 201678 4294 219250 4350
rect 219306 4294 219374 4350
rect 219430 4294 219498 4350
rect 219554 4294 219622 4350
rect 219678 4294 237250 4350
rect 237306 4294 237374 4350
rect 237430 4294 237498 4350
rect 237554 4294 237622 4350
rect 237678 4294 255250 4350
rect 255306 4294 255374 4350
rect 255430 4294 255498 4350
rect 255554 4294 255622 4350
rect 255678 4294 273250 4350
rect 273306 4294 273374 4350
rect 273430 4294 273498 4350
rect 273554 4294 273622 4350
rect 273678 4294 291250 4350
rect 291306 4294 291374 4350
rect 291430 4294 291498 4350
rect 291554 4294 291622 4350
rect 291678 4294 309250 4350
rect 309306 4294 309374 4350
rect 309430 4294 309498 4350
rect 309554 4294 309622 4350
rect 309678 4294 327250 4350
rect 327306 4294 327374 4350
rect 327430 4294 327498 4350
rect 327554 4294 327622 4350
rect 327678 4294 345250 4350
rect 345306 4294 345374 4350
rect 345430 4294 345498 4350
rect 345554 4294 345622 4350
rect 345678 4294 363250 4350
rect 363306 4294 363374 4350
rect 363430 4294 363498 4350
rect 363554 4294 363622 4350
rect 363678 4294 381250 4350
rect 381306 4294 381374 4350
rect 381430 4294 381498 4350
rect 381554 4294 381622 4350
rect 381678 4294 399250 4350
rect 399306 4294 399374 4350
rect 399430 4294 399498 4350
rect 399554 4294 399622 4350
rect 399678 4294 417250 4350
rect 417306 4294 417374 4350
rect 417430 4294 417498 4350
rect 417554 4294 417622 4350
rect 417678 4294 435250 4350
rect 435306 4294 435374 4350
rect 435430 4294 435498 4350
rect 435554 4294 435622 4350
rect 435678 4294 453250 4350
rect 453306 4294 453374 4350
rect 453430 4294 453498 4350
rect 453554 4294 453622 4350
rect 453678 4294 471250 4350
rect 471306 4294 471374 4350
rect 471430 4294 471498 4350
rect 471554 4294 471622 4350
rect 471678 4294 489250 4350
rect 489306 4294 489374 4350
rect 489430 4294 489498 4350
rect 489554 4294 489622 4350
rect 489678 4294 507250 4350
rect 507306 4294 507374 4350
rect 507430 4294 507498 4350
rect 507554 4294 507622 4350
rect 507678 4294 525250 4350
rect 525306 4294 525374 4350
rect 525430 4294 525498 4350
rect 525554 4294 525622 4350
rect 525678 4294 543250 4350
rect 543306 4294 543374 4350
rect 543430 4294 543498 4350
rect 543554 4294 543622 4350
rect 543678 4294 561250 4350
rect 561306 4294 561374 4350
rect 561430 4294 561498 4350
rect 561554 4294 561622 4350
rect 561678 4294 579250 4350
rect 579306 4294 579374 4350
rect 579430 4294 579498 4350
rect 579554 4294 579622 4350
rect 579678 4294 596496 4350
rect 596552 4294 596620 4350
rect 596676 4294 596744 4350
rect 596800 4294 596868 4350
rect 596924 4294 597980 4350
rect -1916 4226 597980 4294
rect -1916 4170 -860 4226
rect -804 4170 -736 4226
rect -680 4170 -612 4226
rect -556 4170 -488 4226
rect -432 4170 3250 4226
rect 3306 4170 3374 4226
rect 3430 4170 3498 4226
rect 3554 4170 3622 4226
rect 3678 4170 21250 4226
rect 21306 4170 21374 4226
rect 21430 4170 21498 4226
rect 21554 4170 21622 4226
rect 21678 4170 39250 4226
rect 39306 4170 39374 4226
rect 39430 4170 39498 4226
rect 39554 4170 39622 4226
rect 39678 4170 57250 4226
rect 57306 4170 57374 4226
rect 57430 4170 57498 4226
rect 57554 4170 57622 4226
rect 57678 4170 75250 4226
rect 75306 4170 75374 4226
rect 75430 4170 75498 4226
rect 75554 4170 75622 4226
rect 75678 4170 93250 4226
rect 93306 4170 93374 4226
rect 93430 4170 93498 4226
rect 93554 4170 93622 4226
rect 93678 4170 111250 4226
rect 111306 4170 111374 4226
rect 111430 4170 111498 4226
rect 111554 4170 111622 4226
rect 111678 4170 129250 4226
rect 129306 4170 129374 4226
rect 129430 4170 129498 4226
rect 129554 4170 129622 4226
rect 129678 4170 147250 4226
rect 147306 4170 147374 4226
rect 147430 4170 147498 4226
rect 147554 4170 147622 4226
rect 147678 4170 165250 4226
rect 165306 4170 165374 4226
rect 165430 4170 165498 4226
rect 165554 4170 165622 4226
rect 165678 4170 183250 4226
rect 183306 4170 183374 4226
rect 183430 4170 183498 4226
rect 183554 4170 183622 4226
rect 183678 4170 201250 4226
rect 201306 4170 201374 4226
rect 201430 4170 201498 4226
rect 201554 4170 201622 4226
rect 201678 4170 219250 4226
rect 219306 4170 219374 4226
rect 219430 4170 219498 4226
rect 219554 4170 219622 4226
rect 219678 4170 237250 4226
rect 237306 4170 237374 4226
rect 237430 4170 237498 4226
rect 237554 4170 237622 4226
rect 237678 4170 255250 4226
rect 255306 4170 255374 4226
rect 255430 4170 255498 4226
rect 255554 4170 255622 4226
rect 255678 4170 273250 4226
rect 273306 4170 273374 4226
rect 273430 4170 273498 4226
rect 273554 4170 273622 4226
rect 273678 4170 291250 4226
rect 291306 4170 291374 4226
rect 291430 4170 291498 4226
rect 291554 4170 291622 4226
rect 291678 4170 309250 4226
rect 309306 4170 309374 4226
rect 309430 4170 309498 4226
rect 309554 4170 309622 4226
rect 309678 4170 327250 4226
rect 327306 4170 327374 4226
rect 327430 4170 327498 4226
rect 327554 4170 327622 4226
rect 327678 4170 345250 4226
rect 345306 4170 345374 4226
rect 345430 4170 345498 4226
rect 345554 4170 345622 4226
rect 345678 4170 363250 4226
rect 363306 4170 363374 4226
rect 363430 4170 363498 4226
rect 363554 4170 363622 4226
rect 363678 4170 381250 4226
rect 381306 4170 381374 4226
rect 381430 4170 381498 4226
rect 381554 4170 381622 4226
rect 381678 4170 399250 4226
rect 399306 4170 399374 4226
rect 399430 4170 399498 4226
rect 399554 4170 399622 4226
rect 399678 4170 417250 4226
rect 417306 4170 417374 4226
rect 417430 4170 417498 4226
rect 417554 4170 417622 4226
rect 417678 4170 435250 4226
rect 435306 4170 435374 4226
rect 435430 4170 435498 4226
rect 435554 4170 435622 4226
rect 435678 4170 453250 4226
rect 453306 4170 453374 4226
rect 453430 4170 453498 4226
rect 453554 4170 453622 4226
rect 453678 4170 471250 4226
rect 471306 4170 471374 4226
rect 471430 4170 471498 4226
rect 471554 4170 471622 4226
rect 471678 4170 489250 4226
rect 489306 4170 489374 4226
rect 489430 4170 489498 4226
rect 489554 4170 489622 4226
rect 489678 4170 507250 4226
rect 507306 4170 507374 4226
rect 507430 4170 507498 4226
rect 507554 4170 507622 4226
rect 507678 4170 525250 4226
rect 525306 4170 525374 4226
rect 525430 4170 525498 4226
rect 525554 4170 525622 4226
rect 525678 4170 543250 4226
rect 543306 4170 543374 4226
rect 543430 4170 543498 4226
rect 543554 4170 543622 4226
rect 543678 4170 561250 4226
rect 561306 4170 561374 4226
rect 561430 4170 561498 4226
rect 561554 4170 561622 4226
rect 561678 4170 579250 4226
rect 579306 4170 579374 4226
rect 579430 4170 579498 4226
rect 579554 4170 579622 4226
rect 579678 4170 596496 4226
rect 596552 4170 596620 4226
rect 596676 4170 596744 4226
rect 596800 4170 596868 4226
rect 596924 4170 597980 4226
rect -1916 4102 597980 4170
rect -1916 4046 -860 4102
rect -804 4046 -736 4102
rect -680 4046 -612 4102
rect -556 4046 -488 4102
rect -432 4046 3250 4102
rect 3306 4046 3374 4102
rect 3430 4046 3498 4102
rect 3554 4046 3622 4102
rect 3678 4046 21250 4102
rect 21306 4046 21374 4102
rect 21430 4046 21498 4102
rect 21554 4046 21622 4102
rect 21678 4046 39250 4102
rect 39306 4046 39374 4102
rect 39430 4046 39498 4102
rect 39554 4046 39622 4102
rect 39678 4046 57250 4102
rect 57306 4046 57374 4102
rect 57430 4046 57498 4102
rect 57554 4046 57622 4102
rect 57678 4046 75250 4102
rect 75306 4046 75374 4102
rect 75430 4046 75498 4102
rect 75554 4046 75622 4102
rect 75678 4046 93250 4102
rect 93306 4046 93374 4102
rect 93430 4046 93498 4102
rect 93554 4046 93622 4102
rect 93678 4046 111250 4102
rect 111306 4046 111374 4102
rect 111430 4046 111498 4102
rect 111554 4046 111622 4102
rect 111678 4046 129250 4102
rect 129306 4046 129374 4102
rect 129430 4046 129498 4102
rect 129554 4046 129622 4102
rect 129678 4046 147250 4102
rect 147306 4046 147374 4102
rect 147430 4046 147498 4102
rect 147554 4046 147622 4102
rect 147678 4046 165250 4102
rect 165306 4046 165374 4102
rect 165430 4046 165498 4102
rect 165554 4046 165622 4102
rect 165678 4046 183250 4102
rect 183306 4046 183374 4102
rect 183430 4046 183498 4102
rect 183554 4046 183622 4102
rect 183678 4046 201250 4102
rect 201306 4046 201374 4102
rect 201430 4046 201498 4102
rect 201554 4046 201622 4102
rect 201678 4046 219250 4102
rect 219306 4046 219374 4102
rect 219430 4046 219498 4102
rect 219554 4046 219622 4102
rect 219678 4046 237250 4102
rect 237306 4046 237374 4102
rect 237430 4046 237498 4102
rect 237554 4046 237622 4102
rect 237678 4046 255250 4102
rect 255306 4046 255374 4102
rect 255430 4046 255498 4102
rect 255554 4046 255622 4102
rect 255678 4046 273250 4102
rect 273306 4046 273374 4102
rect 273430 4046 273498 4102
rect 273554 4046 273622 4102
rect 273678 4046 291250 4102
rect 291306 4046 291374 4102
rect 291430 4046 291498 4102
rect 291554 4046 291622 4102
rect 291678 4046 309250 4102
rect 309306 4046 309374 4102
rect 309430 4046 309498 4102
rect 309554 4046 309622 4102
rect 309678 4046 327250 4102
rect 327306 4046 327374 4102
rect 327430 4046 327498 4102
rect 327554 4046 327622 4102
rect 327678 4046 345250 4102
rect 345306 4046 345374 4102
rect 345430 4046 345498 4102
rect 345554 4046 345622 4102
rect 345678 4046 363250 4102
rect 363306 4046 363374 4102
rect 363430 4046 363498 4102
rect 363554 4046 363622 4102
rect 363678 4046 381250 4102
rect 381306 4046 381374 4102
rect 381430 4046 381498 4102
rect 381554 4046 381622 4102
rect 381678 4046 399250 4102
rect 399306 4046 399374 4102
rect 399430 4046 399498 4102
rect 399554 4046 399622 4102
rect 399678 4046 417250 4102
rect 417306 4046 417374 4102
rect 417430 4046 417498 4102
rect 417554 4046 417622 4102
rect 417678 4046 435250 4102
rect 435306 4046 435374 4102
rect 435430 4046 435498 4102
rect 435554 4046 435622 4102
rect 435678 4046 453250 4102
rect 453306 4046 453374 4102
rect 453430 4046 453498 4102
rect 453554 4046 453622 4102
rect 453678 4046 471250 4102
rect 471306 4046 471374 4102
rect 471430 4046 471498 4102
rect 471554 4046 471622 4102
rect 471678 4046 489250 4102
rect 489306 4046 489374 4102
rect 489430 4046 489498 4102
rect 489554 4046 489622 4102
rect 489678 4046 507250 4102
rect 507306 4046 507374 4102
rect 507430 4046 507498 4102
rect 507554 4046 507622 4102
rect 507678 4046 525250 4102
rect 525306 4046 525374 4102
rect 525430 4046 525498 4102
rect 525554 4046 525622 4102
rect 525678 4046 543250 4102
rect 543306 4046 543374 4102
rect 543430 4046 543498 4102
rect 543554 4046 543622 4102
rect 543678 4046 561250 4102
rect 561306 4046 561374 4102
rect 561430 4046 561498 4102
rect 561554 4046 561622 4102
rect 561678 4046 579250 4102
rect 579306 4046 579374 4102
rect 579430 4046 579498 4102
rect 579554 4046 579622 4102
rect 579678 4046 596496 4102
rect 596552 4046 596620 4102
rect 596676 4046 596744 4102
rect 596800 4046 596868 4102
rect 596924 4046 597980 4102
rect -1916 3978 597980 4046
rect -1916 3922 -860 3978
rect -804 3922 -736 3978
rect -680 3922 -612 3978
rect -556 3922 -488 3978
rect -432 3922 3250 3978
rect 3306 3922 3374 3978
rect 3430 3922 3498 3978
rect 3554 3922 3622 3978
rect 3678 3922 21250 3978
rect 21306 3922 21374 3978
rect 21430 3922 21498 3978
rect 21554 3922 21622 3978
rect 21678 3922 39250 3978
rect 39306 3922 39374 3978
rect 39430 3922 39498 3978
rect 39554 3922 39622 3978
rect 39678 3922 57250 3978
rect 57306 3922 57374 3978
rect 57430 3922 57498 3978
rect 57554 3922 57622 3978
rect 57678 3922 75250 3978
rect 75306 3922 75374 3978
rect 75430 3922 75498 3978
rect 75554 3922 75622 3978
rect 75678 3922 93250 3978
rect 93306 3922 93374 3978
rect 93430 3922 93498 3978
rect 93554 3922 93622 3978
rect 93678 3922 111250 3978
rect 111306 3922 111374 3978
rect 111430 3922 111498 3978
rect 111554 3922 111622 3978
rect 111678 3922 129250 3978
rect 129306 3922 129374 3978
rect 129430 3922 129498 3978
rect 129554 3922 129622 3978
rect 129678 3922 147250 3978
rect 147306 3922 147374 3978
rect 147430 3922 147498 3978
rect 147554 3922 147622 3978
rect 147678 3922 165250 3978
rect 165306 3922 165374 3978
rect 165430 3922 165498 3978
rect 165554 3922 165622 3978
rect 165678 3922 183250 3978
rect 183306 3922 183374 3978
rect 183430 3922 183498 3978
rect 183554 3922 183622 3978
rect 183678 3922 201250 3978
rect 201306 3922 201374 3978
rect 201430 3922 201498 3978
rect 201554 3922 201622 3978
rect 201678 3922 219250 3978
rect 219306 3922 219374 3978
rect 219430 3922 219498 3978
rect 219554 3922 219622 3978
rect 219678 3922 237250 3978
rect 237306 3922 237374 3978
rect 237430 3922 237498 3978
rect 237554 3922 237622 3978
rect 237678 3922 255250 3978
rect 255306 3922 255374 3978
rect 255430 3922 255498 3978
rect 255554 3922 255622 3978
rect 255678 3922 273250 3978
rect 273306 3922 273374 3978
rect 273430 3922 273498 3978
rect 273554 3922 273622 3978
rect 273678 3922 291250 3978
rect 291306 3922 291374 3978
rect 291430 3922 291498 3978
rect 291554 3922 291622 3978
rect 291678 3922 309250 3978
rect 309306 3922 309374 3978
rect 309430 3922 309498 3978
rect 309554 3922 309622 3978
rect 309678 3922 327250 3978
rect 327306 3922 327374 3978
rect 327430 3922 327498 3978
rect 327554 3922 327622 3978
rect 327678 3922 345250 3978
rect 345306 3922 345374 3978
rect 345430 3922 345498 3978
rect 345554 3922 345622 3978
rect 345678 3922 363250 3978
rect 363306 3922 363374 3978
rect 363430 3922 363498 3978
rect 363554 3922 363622 3978
rect 363678 3922 381250 3978
rect 381306 3922 381374 3978
rect 381430 3922 381498 3978
rect 381554 3922 381622 3978
rect 381678 3922 399250 3978
rect 399306 3922 399374 3978
rect 399430 3922 399498 3978
rect 399554 3922 399622 3978
rect 399678 3922 417250 3978
rect 417306 3922 417374 3978
rect 417430 3922 417498 3978
rect 417554 3922 417622 3978
rect 417678 3922 435250 3978
rect 435306 3922 435374 3978
rect 435430 3922 435498 3978
rect 435554 3922 435622 3978
rect 435678 3922 453250 3978
rect 453306 3922 453374 3978
rect 453430 3922 453498 3978
rect 453554 3922 453622 3978
rect 453678 3922 471250 3978
rect 471306 3922 471374 3978
rect 471430 3922 471498 3978
rect 471554 3922 471622 3978
rect 471678 3922 489250 3978
rect 489306 3922 489374 3978
rect 489430 3922 489498 3978
rect 489554 3922 489622 3978
rect 489678 3922 507250 3978
rect 507306 3922 507374 3978
rect 507430 3922 507498 3978
rect 507554 3922 507622 3978
rect 507678 3922 525250 3978
rect 525306 3922 525374 3978
rect 525430 3922 525498 3978
rect 525554 3922 525622 3978
rect 525678 3922 543250 3978
rect 543306 3922 543374 3978
rect 543430 3922 543498 3978
rect 543554 3922 543622 3978
rect 543678 3922 561250 3978
rect 561306 3922 561374 3978
rect 561430 3922 561498 3978
rect 561554 3922 561622 3978
rect 561678 3922 579250 3978
rect 579306 3922 579374 3978
rect 579430 3922 579498 3978
rect 579554 3922 579622 3978
rect 579678 3922 596496 3978
rect 596552 3922 596620 3978
rect 596676 3922 596744 3978
rect 596800 3922 596868 3978
rect 596924 3922 597980 3978
rect -1916 3826 597980 3922
rect -956 -160 597020 -64
rect -956 -216 -860 -160
rect -804 -216 -736 -160
rect -680 -216 -612 -160
rect -556 -216 -488 -160
rect -432 -216 3250 -160
rect 3306 -216 3374 -160
rect 3430 -216 3498 -160
rect 3554 -216 3622 -160
rect 3678 -216 21250 -160
rect 21306 -216 21374 -160
rect 21430 -216 21498 -160
rect 21554 -216 21622 -160
rect 21678 -216 39250 -160
rect 39306 -216 39374 -160
rect 39430 -216 39498 -160
rect 39554 -216 39622 -160
rect 39678 -216 57250 -160
rect 57306 -216 57374 -160
rect 57430 -216 57498 -160
rect 57554 -216 57622 -160
rect 57678 -216 75250 -160
rect 75306 -216 75374 -160
rect 75430 -216 75498 -160
rect 75554 -216 75622 -160
rect 75678 -216 93250 -160
rect 93306 -216 93374 -160
rect 93430 -216 93498 -160
rect 93554 -216 93622 -160
rect 93678 -216 111250 -160
rect 111306 -216 111374 -160
rect 111430 -216 111498 -160
rect 111554 -216 111622 -160
rect 111678 -216 129250 -160
rect 129306 -216 129374 -160
rect 129430 -216 129498 -160
rect 129554 -216 129622 -160
rect 129678 -216 147250 -160
rect 147306 -216 147374 -160
rect 147430 -216 147498 -160
rect 147554 -216 147622 -160
rect 147678 -216 165250 -160
rect 165306 -216 165374 -160
rect 165430 -216 165498 -160
rect 165554 -216 165622 -160
rect 165678 -216 183250 -160
rect 183306 -216 183374 -160
rect 183430 -216 183498 -160
rect 183554 -216 183622 -160
rect 183678 -216 201250 -160
rect 201306 -216 201374 -160
rect 201430 -216 201498 -160
rect 201554 -216 201622 -160
rect 201678 -216 219250 -160
rect 219306 -216 219374 -160
rect 219430 -216 219498 -160
rect 219554 -216 219622 -160
rect 219678 -216 237250 -160
rect 237306 -216 237374 -160
rect 237430 -216 237498 -160
rect 237554 -216 237622 -160
rect 237678 -216 255250 -160
rect 255306 -216 255374 -160
rect 255430 -216 255498 -160
rect 255554 -216 255622 -160
rect 255678 -216 273250 -160
rect 273306 -216 273374 -160
rect 273430 -216 273498 -160
rect 273554 -216 273622 -160
rect 273678 -216 291250 -160
rect 291306 -216 291374 -160
rect 291430 -216 291498 -160
rect 291554 -216 291622 -160
rect 291678 -216 309250 -160
rect 309306 -216 309374 -160
rect 309430 -216 309498 -160
rect 309554 -216 309622 -160
rect 309678 -216 327250 -160
rect 327306 -216 327374 -160
rect 327430 -216 327498 -160
rect 327554 -216 327622 -160
rect 327678 -216 345250 -160
rect 345306 -216 345374 -160
rect 345430 -216 345498 -160
rect 345554 -216 345622 -160
rect 345678 -216 363250 -160
rect 363306 -216 363374 -160
rect 363430 -216 363498 -160
rect 363554 -216 363622 -160
rect 363678 -216 381250 -160
rect 381306 -216 381374 -160
rect 381430 -216 381498 -160
rect 381554 -216 381622 -160
rect 381678 -216 399250 -160
rect 399306 -216 399374 -160
rect 399430 -216 399498 -160
rect 399554 -216 399622 -160
rect 399678 -216 417250 -160
rect 417306 -216 417374 -160
rect 417430 -216 417498 -160
rect 417554 -216 417622 -160
rect 417678 -216 435250 -160
rect 435306 -216 435374 -160
rect 435430 -216 435498 -160
rect 435554 -216 435622 -160
rect 435678 -216 453250 -160
rect 453306 -216 453374 -160
rect 453430 -216 453498 -160
rect 453554 -216 453622 -160
rect 453678 -216 471250 -160
rect 471306 -216 471374 -160
rect 471430 -216 471498 -160
rect 471554 -216 471622 -160
rect 471678 -216 489250 -160
rect 489306 -216 489374 -160
rect 489430 -216 489498 -160
rect 489554 -216 489622 -160
rect 489678 -216 507250 -160
rect 507306 -216 507374 -160
rect 507430 -216 507498 -160
rect 507554 -216 507622 -160
rect 507678 -216 525250 -160
rect 525306 -216 525374 -160
rect 525430 -216 525498 -160
rect 525554 -216 525622 -160
rect 525678 -216 543250 -160
rect 543306 -216 543374 -160
rect 543430 -216 543498 -160
rect 543554 -216 543622 -160
rect 543678 -216 561250 -160
rect 561306 -216 561374 -160
rect 561430 -216 561498 -160
rect 561554 -216 561622 -160
rect 561678 -216 579250 -160
rect 579306 -216 579374 -160
rect 579430 -216 579498 -160
rect 579554 -216 579622 -160
rect 579678 -216 596496 -160
rect 596552 -216 596620 -160
rect 596676 -216 596744 -160
rect 596800 -216 596868 -160
rect 596924 -216 597020 -160
rect -956 -284 597020 -216
rect -956 -340 -860 -284
rect -804 -340 -736 -284
rect -680 -340 -612 -284
rect -556 -340 -488 -284
rect -432 -340 3250 -284
rect 3306 -340 3374 -284
rect 3430 -340 3498 -284
rect 3554 -340 3622 -284
rect 3678 -340 21250 -284
rect 21306 -340 21374 -284
rect 21430 -340 21498 -284
rect 21554 -340 21622 -284
rect 21678 -340 39250 -284
rect 39306 -340 39374 -284
rect 39430 -340 39498 -284
rect 39554 -340 39622 -284
rect 39678 -340 57250 -284
rect 57306 -340 57374 -284
rect 57430 -340 57498 -284
rect 57554 -340 57622 -284
rect 57678 -340 75250 -284
rect 75306 -340 75374 -284
rect 75430 -340 75498 -284
rect 75554 -340 75622 -284
rect 75678 -340 93250 -284
rect 93306 -340 93374 -284
rect 93430 -340 93498 -284
rect 93554 -340 93622 -284
rect 93678 -340 111250 -284
rect 111306 -340 111374 -284
rect 111430 -340 111498 -284
rect 111554 -340 111622 -284
rect 111678 -340 129250 -284
rect 129306 -340 129374 -284
rect 129430 -340 129498 -284
rect 129554 -340 129622 -284
rect 129678 -340 147250 -284
rect 147306 -340 147374 -284
rect 147430 -340 147498 -284
rect 147554 -340 147622 -284
rect 147678 -340 165250 -284
rect 165306 -340 165374 -284
rect 165430 -340 165498 -284
rect 165554 -340 165622 -284
rect 165678 -340 183250 -284
rect 183306 -340 183374 -284
rect 183430 -340 183498 -284
rect 183554 -340 183622 -284
rect 183678 -340 201250 -284
rect 201306 -340 201374 -284
rect 201430 -340 201498 -284
rect 201554 -340 201622 -284
rect 201678 -340 219250 -284
rect 219306 -340 219374 -284
rect 219430 -340 219498 -284
rect 219554 -340 219622 -284
rect 219678 -340 237250 -284
rect 237306 -340 237374 -284
rect 237430 -340 237498 -284
rect 237554 -340 237622 -284
rect 237678 -340 255250 -284
rect 255306 -340 255374 -284
rect 255430 -340 255498 -284
rect 255554 -340 255622 -284
rect 255678 -340 273250 -284
rect 273306 -340 273374 -284
rect 273430 -340 273498 -284
rect 273554 -340 273622 -284
rect 273678 -340 291250 -284
rect 291306 -340 291374 -284
rect 291430 -340 291498 -284
rect 291554 -340 291622 -284
rect 291678 -340 309250 -284
rect 309306 -340 309374 -284
rect 309430 -340 309498 -284
rect 309554 -340 309622 -284
rect 309678 -340 327250 -284
rect 327306 -340 327374 -284
rect 327430 -340 327498 -284
rect 327554 -340 327622 -284
rect 327678 -340 345250 -284
rect 345306 -340 345374 -284
rect 345430 -340 345498 -284
rect 345554 -340 345622 -284
rect 345678 -340 363250 -284
rect 363306 -340 363374 -284
rect 363430 -340 363498 -284
rect 363554 -340 363622 -284
rect 363678 -340 381250 -284
rect 381306 -340 381374 -284
rect 381430 -340 381498 -284
rect 381554 -340 381622 -284
rect 381678 -340 399250 -284
rect 399306 -340 399374 -284
rect 399430 -340 399498 -284
rect 399554 -340 399622 -284
rect 399678 -340 417250 -284
rect 417306 -340 417374 -284
rect 417430 -340 417498 -284
rect 417554 -340 417622 -284
rect 417678 -340 435250 -284
rect 435306 -340 435374 -284
rect 435430 -340 435498 -284
rect 435554 -340 435622 -284
rect 435678 -340 453250 -284
rect 453306 -340 453374 -284
rect 453430 -340 453498 -284
rect 453554 -340 453622 -284
rect 453678 -340 471250 -284
rect 471306 -340 471374 -284
rect 471430 -340 471498 -284
rect 471554 -340 471622 -284
rect 471678 -340 489250 -284
rect 489306 -340 489374 -284
rect 489430 -340 489498 -284
rect 489554 -340 489622 -284
rect 489678 -340 507250 -284
rect 507306 -340 507374 -284
rect 507430 -340 507498 -284
rect 507554 -340 507622 -284
rect 507678 -340 525250 -284
rect 525306 -340 525374 -284
rect 525430 -340 525498 -284
rect 525554 -340 525622 -284
rect 525678 -340 543250 -284
rect 543306 -340 543374 -284
rect 543430 -340 543498 -284
rect 543554 -340 543622 -284
rect 543678 -340 561250 -284
rect 561306 -340 561374 -284
rect 561430 -340 561498 -284
rect 561554 -340 561622 -284
rect 561678 -340 579250 -284
rect 579306 -340 579374 -284
rect 579430 -340 579498 -284
rect 579554 -340 579622 -284
rect 579678 -340 596496 -284
rect 596552 -340 596620 -284
rect 596676 -340 596744 -284
rect 596800 -340 596868 -284
rect 596924 -340 597020 -284
rect -956 -408 597020 -340
rect -956 -464 -860 -408
rect -804 -464 -736 -408
rect -680 -464 -612 -408
rect -556 -464 -488 -408
rect -432 -464 3250 -408
rect 3306 -464 3374 -408
rect 3430 -464 3498 -408
rect 3554 -464 3622 -408
rect 3678 -464 21250 -408
rect 21306 -464 21374 -408
rect 21430 -464 21498 -408
rect 21554 -464 21622 -408
rect 21678 -464 39250 -408
rect 39306 -464 39374 -408
rect 39430 -464 39498 -408
rect 39554 -464 39622 -408
rect 39678 -464 57250 -408
rect 57306 -464 57374 -408
rect 57430 -464 57498 -408
rect 57554 -464 57622 -408
rect 57678 -464 75250 -408
rect 75306 -464 75374 -408
rect 75430 -464 75498 -408
rect 75554 -464 75622 -408
rect 75678 -464 93250 -408
rect 93306 -464 93374 -408
rect 93430 -464 93498 -408
rect 93554 -464 93622 -408
rect 93678 -464 111250 -408
rect 111306 -464 111374 -408
rect 111430 -464 111498 -408
rect 111554 -464 111622 -408
rect 111678 -464 129250 -408
rect 129306 -464 129374 -408
rect 129430 -464 129498 -408
rect 129554 -464 129622 -408
rect 129678 -464 147250 -408
rect 147306 -464 147374 -408
rect 147430 -464 147498 -408
rect 147554 -464 147622 -408
rect 147678 -464 165250 -408
rect 165306 -464 165374 -408
rect 165430 -464 165498 -408
rect 165554 -464 165622 -408
rect 165678 -464 183250 -408
rect 183306 -464 183374 -408
rect 183430 -464 183498 -408
rect 183554 -464 183622 -408
rect 183678 -464 201250 -408
rect 201306 -464 201374 -408
rect 201430 -464 201498 -408
rect 201554 -464 201622 -408
rect 201678 -464 219250 -408
rect 219306 -464 219374 -408
rect 219430 -464 219498 -408
rect 219554 -464 219622 -408
rect 219678 -464 237250 -408
rect 237306 -464 237374 -408
rect 237430 -464 237498 -408
rect 237554 -464 237622 -408
rect 237678 -464 255250 -408
rect 255306 -464 255374 -408
rect 255430 -464 255498 -408
rect 255554 -464 255622 -408
rect 255678 -464 273250 -408
rect 273306 -464 273374 -408
rect 273430 -464 273498 -408
rect 273554 -464 273622 -408
rect 273678 -464 291250 -408
rect 291306 -464 291374 -408
rect 291430 -464 291498 -408
rect 291554 -464 291622 -408
rect 291678 -464 309250 -408
rect 309306 -464 309374 -408
rect 309430 -464 309498 -408
rect 309554 -464 309622 -408
rect 309678 -464 327250 -408
rect 327306 -464 327374 -408
rect 327430 -464 327498 -408
rect 327554 -464 327622 -408
rect 327678 -464 345250 -408
rect 345306 -464 345374 -408
rect 345430 -464 345498 -408
rect 345554 -464 345622 -408
rect 345678 -464 363250 -408
rect 363306 -464 363374 -408
rect 363430 -464 363498 -408
rect 363554 -464 363622 -408
rect 363678 -464 381250 -408
rect 381306 -464 381374 -408
rect 381430 -464 381498 -408
rect 381554 -464 381622 -408
rect 381678 -464 399250 -408
rect 399306 -464 399374 -408
rect 399430 -464 399498 -408
rect 399554 -464 399622 -408
rect 399678 -464 417250 -408
rect 417306 -464 417374 -408
rect 417430 -464 417498 -408
rect 417554 -464 417622 -408
rect 417678 -464 435250 -408
rect 435306 -464 435374 -408
rect 435430 -464 435498 -408
rect 435554 -464 435622 -408
rect 435678 -464 453250 -408
rect 453306 -464 453374 -408
rect 453430 -464 453498 -408
rect 453554 -464 453622 -408
rect 453678 -464 471250 -408
rect 471306 -464 471374 -408
rect 471430 -464 471498 -408
rect 471554 -464 471622 -408
rect 471678 -464 489250 -408
rect 489306 -464 489374 -408
rect 489430 -464 489498 -408
rect 489554 -464 489622 -408
rect 489678 -464 507250 -408
rect 507306 -464 507374 -408
rect 507430 -464 507498 -408
rect 507554 -464 507622 -408
rect 507678 -464 525250 -408
rect 525306 -464 525374 -408
rect 525430 -464 525498 -408
rect 525554 -464 525622 -408
rect 525678 -464 543250 -408
rect 543306 -464 543374 -408
rect 543430 -464 543498 -408
rect 543554 -464 543622 -408
rect 543678 -464 561250 -408
rect 561306 -464 561374 -408
rect 561430 -464 561498 -408
rect 561554 -464 561622 -408
rect 561678 -464 579250 -408
rect 579306 -464 579374 -408
rect 579430 -464 579498 -408
rect 579554 -464 579622 -408
rect 579678 -464 596496 -408
rect 596552 -464 596620 -408
rect 596676 -464 596744 -408
rect 596800 -464 596868 -408
rect 596924 -464 597020 -408
rect -956 -532 597020 -464
rect -956 -588 -860 -532
rect -804 -588 -736 -532
rect -680 -588 -612 -532
rect -556 -588 -488 -532
rect -432 -588 3250 -532
rect 3306 -588 3374 -532
rect 3430 -588 3498 -532
rect 3554 -588 3622 -532
rect 3678 -588 21250 -532
rect 21306 -588 21374 -532
rect 21430 -588 21498 -532
rect 21554 -588 21622 -532
rect 21678 -588 39250 -532
rect 39306 -588 39374 -532
rect 39430 -588 39498 -532
rect 39554 -588 39622 -532
rect 39678 -588 57250 -532
rect 57306 -588 57374 -532
rect 57430 -588 57498 -532
rect 57554 -588 57622 -532
rect 57678 -588 75250 -532
rect 75306 -588 75374 -532
rect 75430 -588 75498 -532
rect 75554 -588 75622 -532
rect 75678 -588 93250 -532
rect 93306 -588 93374 -532
rect 93430 -588 93498 -532
rect 93554 -588 93622 -532
rect 93678 -588 111250 -532
rect 111306 -588 111374 -532
rect 111430 -588 111498 -532
rect 111554 -588 111622 -532
rect 111678 -588 129250 -532
rect 129306 -588 129374 -532
rect 129430 -588 129498 -532
rect 129554 -588 129622 -532
rect 129678 -588 147250 -532
rect 147306 -588 147374 -532
rect 147430 -588 147498 -532
rect 147554 -588 147622 -532
rect 147678 -588 165250 -532
rect 165306 -588 165374 -532
rect 165430 -588 165498 -532
rect 165554 -588 165622 -532
rect 165678 -588 183250 -532
rect 183306 -588 183374 -532
rect 183430 -588 183498 -532
rect 183554 -588 183622 -532
rect 183678 -588 201250 -532
rect 201306 -588 201374 -532
rect 201430 -588 201498 -532
rect 201554 -588 201622 -532
rect 201678 -588 219250 -532
rect 219306 -588 219374 -532
rect 219430 -588 219498 -532
rect 219554 -588 219622 -532
rect 219678 -588 237250 -532
rect 237306 -588 237374 -532
rect 237430 -588 237498 -532
rect 237554 -588 237622 -532
rect 237678 -588 255250 -532
rect 255306 -588 255374 -532
rect 255430 -588 255498 -532
rect 255554 -588 255622 -532
rect 255678 -588 273250 -532
rect 273306 -588 273374 -532
rect 273430 -588 273498 -532
rect 273554 -588 273622 -532
rect 273678 -588 291250 -532
rect 291306 -588 291374 -532
rect 291430 -588 291498 -532
rect 291554 -588 291622 -532
rect 291678 -588 309250 -532
rect 309306 -588 309374 -532
rect 309430 -588 309498 -532
rect 309554 -588 309622 -532
rect 309678 -588 327250 -532
rect 327306 -588 327374 -532
rect 327430 -588 327498 -532
rect 327554 -588 327622 -532
rect 327678 -588 345250 -532
rect 345306 -588 345374 -532
rect 345430 -588 345498 -532
rect 345554 -588 345622 -532
rect 345678 -588 363250 -532
rect 363306 -588 363374 -532
rect 363430 -588 363498 -532
rect 363554 -588 363622 -532
rect 363678 -588 381250 -532
rect 381306 -588 381374 -532
rect 381430 -588 381498 -532
rect 381554 -588 381622 -532
rect 381678 -588 399250 -532
rect 399306 -588 399374 -532
rect 399430 -588 399498 -532
rect 399554 -588 399622 -532
rect 399678 -588 417250 -532
rect 417306 -588 417374 -532
rect 417430 -588 417498 -532
rect 417554 -588 417622 -532
rect 417678 -588 435250 -532
rect 435306 -588 435374 -532
rect 435430 -588 435498 -532
rect 435554 -588 435622 -532
rect 435678 -588 453250 -532
rect 453306 -588 453374 -532
rect 453430 -588 453498 -532
rect 453554 -588 453622 -532
rect 453678 -588 471250 -532
rect 471306 -588 471374 -532
rect 471430 -588 471498 -532
rect 471554 -588 471622 -532
rect 471678 -588 489250 -532
rect 489306 -588 489374 -532
rect 489430 -588 489498 -532
rect 489554 -588 489622 -532
rect 489678 -588 507250 -532
rect 507306 -588 507374 -532
rect 507430 -588 507498 -532
rect 507554 -588 507622 -532
rect 507678 -588 525250 -532
rect 525306 -588 525374 -532
rect 525430 -588 525498 -532
rect 525554 -588 525622 -532
rect 525678 -588 543250 -532
rect 543306 -588 543374 -532
rect 543430 -588 543498 -532
rect 543554 -588 543622 -532
rect 543678 -588 561250 -532
rect 561306 -588 561374 -532
rect 561430 -588 561498 -532
rect 561554 -588 561622 -532
rect 561678 -588 579250 -532
rect 579306 -588 579374 -532
rect 579430 -588 579498 -532
rect 579554 -588 579622 -532
rect 579678 -588 596496 -532
rect 596552 -588 596620 -532
rect 596676 -588 596744 -532
rect 596800 -588 596868 -532
rect 596924 -588 597020 -532
rect -956 -684 597020 -588
rect -1916 -1120 597980 -1024
rect -1916 -1176 -1820 -1120
rect -1764 -1176 -1696 -1120
rect -1640 -1176 -1572 -1120
rect -1516 -1176 -1448 -1120
rect -1392 -1176 6970 -1120
rect 7026 -1176 7094 -1120
rect 7150 -1176 7218 -1120
rect 7274 -1176 7342 -1120
rect 7398 -1176 24970 -1120
rect 25026 -1176 25094 -1120
rect 25150 -1176 25218 -1120
rect 25274 -1176 25342 -1120
rect 25398 -1176 42970 -1120
rect 43026 -1176 43094 -1120
rect 43150 -1176 43218 -1120
rect 43274 -1176 43342 -1120
rect 43398 -1176 60970 -1120
rect 61026 -1176 61094 -1120
rect 61150 -1176 61218 -1120
rect 61274 -1176 61342 -1120
rect 61398 -1176 78970 -1120
rect 79026 -1176 79094 -1120
rect 79150 -1176 79218 -1120
rect 79274 -1176 79342 -1120
rect 79398 -1176 96970 -1120
rect 97026 -1176 97094 -1120
rect 97150 -1176 97218 -1120
rect 97274 -1176 97342 -1120
rect 97398 -1176 114970 -1120
rect 115026 -1176 115094 -1120
rect 115150 -1176 115218 -1120
rect 115274 -1176 115342 -1120
rect 115398 -1176 132970 -1120
rect 133026 -1176 133094 -1120
rect 133150 -1176 133218 -1120
rect 133274 -1176 133342 -1120
rect 133398 -1176 150970 -1120
rect 151026 -1176 151094 -1120
rect 151150 -1176 151218 -1120
rect 151274 -1176 151342 -1120
rect 151398 -1176 168970 -1120
rect 169026 -1176 169094 -1120
rect 169150 -1176 169218 -1120
rect 169274 -1176 169342 -1120
rect 169398 -1176 186970 -1120
rect 187026 -1176 187094 -1120
rect 187150 -1176 187218 -1120
rect 187274 -1176 187342 -1120
rect 187398 -1176 204970 -1120
rect 205026 -1176 205094 -1120
rect 205150 -1176 205218 -1120
rect 205274 -1176 205342 -1120
rect 205398 -1176 222970 -1120
rect 223026 -1176 223094 -1120
rect 223150 -1176 223218 -1120
rect 223274 -1176 223342 -1120
rect 223398 -1176 240970 -1120
rect 241026 -1176 241094 -1120
rect 241150 -1176 241218 -1120
rect 241274 -1176 241342 -1120
rect 241398 -1176 258970 -1120
rect 259026 -1176 259094 -1120
rect 259150 -1176 259218 -1120
rect 259274 -1176 259342 -1120
rect 259398 -1176 276970 -1120
rect 277026 -1176 277094 -1120
rect 277150 -1176 277218 -1120
rect 277274 -1176 277342 -1120
rect 277398 -1176 294970 -1120
rect 295026 -1176 295094 -1120
rect 295150 -1176 295218 -1120
rect 295274 -1176 295342 -1120
rect 295398 -1176 312970 -1120
rect 313026 -1176 313094 -1120
rect 313150 -1176 313218 -1120
rect 313274 -1176 313342 -1120
rect 313398 -1176 330970 -1120
rect 331026 -1176 331094 -1120
rect 331150 -1176 331218 -1120
rect 331274 -1176 331342 -1120
rect 331398 -1176 348970 -1120
rect 349026 -1176 349094 -1120
rect 349150 -1176 349218 -1120
rect 349274 -1176 349342 -1120
rect 349398 -1176 366970 -1120
rect 367026 -1176 367094 -1120
rect 367150 -1176 367218 -1120
rect 367274 -1176 367342 -1120
rect 367398 -1176 384970 -1120
rect 385026 -1176 385094 -1120
rect 385150 -1176 385218 -1120
rect 385274 -1176 385342 -1120
rect 385398 -1176 402970 -1120
rect 403026 -1176 403094 -1120
rect 403150 -1176 403218 -1120
rect 403274 -1176 403342 -1120
rect 403398 -1176 420970 -1120
rect 421026 -1176 421094 -1120
rect 421150 -1176 421218 -1120
rect 421274 -1176 421342 -1120
rect 421398 -1176 438970 -1120
rect 439026 -1176 439094 -1120
rect 439150 -1176 439218 -1120
rect 439274 -1176 439342 -1120
rect 439398 -1176 456970 -1120
rect 457026 -1176 457094 -1120
rect 457150 -1176 457218 -1120
rect 457274 -1176 457342 -1120
rect 457398 -1176 474970 -1120
rect 475026 -1176 475094 -1120
rect 475150 -1176 475218 -1120
rect 475274 -1176 475342 -1120
rect 475398 -1176 492970 -1120
rect 493026 -1176 493094 -1120
rect 493150 -1176 493218 -1120
rect 493274 -1176 493342 -1120
rect 493398 -1176 510970 -1120
rect 511026 -1176 511094 -1120
rect 511150 -1176 511218 -1120
rect 511274 -1176 511342 -1120
rect 511398 -1176 528970 -1120
rect 529026 -1176 529094 -1120
rect 529150 -1176 529218 -1120
rect 529274 -1176 529342 -1120
rect 529398 -1176 546970 -1120
rect 547026 -1176 547094 -1120
rect 547150 -1176 547218 -1120
rect 547274 -1176 547342 -1120
rect 547398 -1176 564970 -1120
rect 565026 -1176 565094 -1120
rect 565150 -1176 565218 -1120
rect 565274 -1176 565342 -1120
rect 565398 -1176 582970 -1120
rect 583026 -1176 583094 -1120
rect 583150 -1176 583218 -1120
rect 583274 -1176 583342 -1120
rect 583398 -1176 597456 -1120
rect 597512 -1176 597580 -1120
rect 597636 -1176 597704 -1120
rect 597760 -1176 597828 -1120
rect 597884 -1176 597980 -1120
rect -1916 -1244 597980 -1176
rect -1916 -1300 -1820 -1244
rect -1764 -1300 -1696 -1244
rect -1640 -1300 -1572 -1244
rect -1516 -1300 -1448 -1244
rect -1392 -1300 6970 -1244
rect 7026 -1300 7094 -1244
rect 7150 -1300 7218 -1244
rect 7274 -1300 7342 -1244
rect 7398 -1300 24970 -1244
rect 25026 -1300 25094 -1244
rect 25150 -1300 25218 -1244
rect 25274 -1300 25342 -1244
rect 25398 -1300 42970 -1244
rect 43026 -1300 43094 -1244
rect 43150 -1300 43218 -1244
rect 43274 -1300 43342 -1244
rect 43398 -1300 60970 -1244
rect 61026 -1300 61094 -1244
rect 61150 -1300 61218 -1244
rect 61274 -1300 61342 -1244
rect 61398 -1300 78970 -1244
rect 79026 -1300 79094 -1244
rect 79150 -1300 79218 -1244
rect 79274 -1300 79342 -1244
rect 79398 -1300 96970 -1244
rect 97026 -1300 97094 -1244
rect 97150 -1300 97218 -1244
rect 97274 -1300 97342 -1244
rect 97398 -1300 114970 -1244
rect 115026 -1300 115094 -1244
rect 115150 -1300 115218 -1244
rect 115274 -1300 115342 -1244
rect 115398 -1300 132970 -1244
rect 133026 -1300 133094 -1244
rect 133150 -1300 133218 -1244
rect 133274 -1300 133342 -1244
rect 133398 -1300 150970 -1244
rect 151026 -1300 151094 -1244
rect 151150 -1300 151218 -1244
rect 151274 -1300 151342 -1244
rect 151398 -1300 168970 -1244
rect 169026 -1300 169094 -1244
rect 169150 -1300 169218 -1244
rect 169274 -1300 169342 -1244
rect 169398 -1300 186970 -1244
rect 187026 -1300 187094 -1244
rect 187150 -1300 187218 -1244
rect 187274 -1300 187342 -1244
rect 187398 -1300 204970 -1244
rect 205026 -1300 205094 -1244
rect 205150 -1300 205218 -1244
rect 205274 -1300 205342 -1244
rect 205398 -1300 222970 -1244
rect 223026 -1300 223094 -1244
rect 223150 -1300 223218 -1244
rect 223274 -1300 223342 -1244
rect 223398 -1300 240970 -1244
rect 241026 -1300 241094 -1244
rect 241150 -1300 241218 -1244
rect 241274 -1300 241342 -1244
rect 241398 -1300 258970 -1244
rect 259026 -1300 259094 -1244
rect 259150 -1300 259218 -1244
rect 259274 -1300 259342 -1244
rect 259398 -1300 276970 -1244
rect 277026 -1300 277094 -1244
rect 277150 -1300 277218 -1244
rect 277274 -1300 277342 -1244
rect 277398 -1300 294970 -1244
rect 295026 -1300 295094 -1244
rect 295150 -1300 295218 -1244
rect 295274 -1300 295342 -1244
rect 295398 -1300 312970 -1244
rect 313026 -1300 313094 -1244
rect 313150 -1300 313218 -1244
rect 313274 -1300 313342 -1244
rect 313398 -1300 330970 -1244
rect 331026 -1300 331094 -1244
rect 331150 -1300 331218 -1244
rect 331274 -1300 331342 -1244
rect 331398 -1300 348970 -1244
rect 349026 -1300 349094 -1244
rect 349150 -1300 349218 -1244
rect 349274 -1300 349342 -1244
rect 349398 -1300 366970 -1244
rect 367026 -1300 367094 -1244
rect 367150 -1300 367218 -1244
rect 367274 -1300 367342 -1244
rect 367398 -1300 384970 -1244
rect 385026 -1300 385094 -1244
rect 385150 -1300 385218 -1244
rect 385274 -1300 385342 -1244
rect 385398 -1300 402970 -1244
rect 403026 -1300 403094 -1244
rect 403150 -1300 403218 -1244
rect 403274 -1300 403342 -1244
rect 403398 -1300 420970 -1244
rect 421026 -1300 421094 -1244
rect 421150 -1300 421218 -1244
rect 421274 -1300 421342 -1244
rect 421398 -1300 438970 -1244
rect 439026 -1300 439094 -1244
rect 439150 -1300 439218 -1244
rect 439274 -1300 439342 -1244
rect 439398 -1300 456970 -1244
rect 457026 -1300 457094 -1244
rect 457150 -1300 457218 -1244
rect 457274 -1300 457342 -1244
rect 457398 -1300 474970 -1244
rect 475026 -1300 475094 -1244
rect 475150 -1300 475218 -1244
rect 475274 -1300 475342 -1244
rect 475398 -1300 492970 -1244
rect 493026 -1300 493094 -1244
rect 493150 -1300 493218 -1244
rect 493274 -1300 493342 -1244
rect 493398 -1300 510970 -1244
rect 511026 -1300 511094 -1244
rect 511150 -1300 511218 -1244
rect 511274 -1300 511342 -1244
rect 511398 -1300 528970 -1244
rect 529026 -1300 529094 -1244
rect 529150 -1300 529218 -1244
rect 529274 -1300 529342 -1244
rect 529398 -1300 546970 -1244
rect 547026 -1300 547094 -1244
rect 547150 -1300 547218 -1244
rect 547274 -1300 547342 -1244
rect 547398 -1300 564970 -1244
rect 565026 -1300 565094 -1244
rect 565150 -1300 565218 -1244
rect 565274 -1300 565342 -1244
rect 565398 -1300 582970 -1244
rect 583026 -1300 583094 -1244
rect 583150 -1300 583218 -1244
rect 583274 -1300 583342 -1244
rect 583398 -1300 597456 -1244
rect 597512 -1300 597580 -1244
rect 597636 -1300 597704 -1244
rect 597760 -1300 597828 -1244
rect 597884 -1300 597980 -1244
rect -1916 -1368 597980 -1300
rect -1916 -1424 -1820 -1368
rect -1764 -1424 -1696 -1368
rect -1640 -1424 -1572 -1368
rect -1516 -1424 -1448 -1368
rect -1392 -1424 6970 -1368
rect 7026 -1424 7094 -1368
rect 7150 -1424 7218 -1368
rect 7274 -1424 7342 -1368
rect 7398 -1424 24970 -1368
rect 25026 -1424 25094 -1368
rect 25150 -1424 25218 -1368
rect 25274 -1424 25342 -1368
rect 25398 -1424 42970 -1368
rect 43026 -1424 43094 -1368
rect 43150 -1424 43218 -1368
rect 43274 -1424 43342 -1368
rect 43398 -1424 60970 -1368
rect 61026 -1424 61094 -1368
rect 61150 -1424 61218 -1368
rect 61274 -1424 61342 -1368
rect 61398 -1424 78970 -1368
rect 79026 -1424 79094 -1368
rect 79150 -1424 79218 -1368
rect 79274 -1424 79342 -1368
rect 79398 -1424 96970 -1368
rect 97026 -1424 97094 -1368
rect 97150 -1424 97218 -1368
rect 97274 -1424 97342 -1368
rect 97398 -1424 114970 -1368
rect 115026 -1424 115094 -1368
rect 115150 -1424 115218 -1368
rect 115274 -1424 115342 -1368
rect 115398 -1424 132970 -1368
rect 133026 -1424 133094 -1368
rect 133150 -1424 133218 -1368
rect 133274 -1424 133342 -1368
rect 133398 -1424 150970 -1368
rect 151026 -1424 151094 -1368
rect 151150 -1424 151218 -1368
rect 151274 -1424 151342 -1368
rect 151398 -1424 168970 -1368
rect 169026 -1424 169094 -1368
rect 169150 -1424 169218 -1368
rect 169274 -1424 169342 -1368
rect 169398 -1424 186970 -1368
rect 187026 -1424 187094 -1368
rect 187150 -1424 187218 -1368
rect 187274 -1424 187342 -1368
rect 187398 -1424 204970 -1368
rect 205026 -1424 205094 -1368
rect 205150 -1424 205218 -1368
rect 205274 -1424 205342 -1368
rect 205398 -1424 222970 -1368
rect 223026 -1424 223094 -1368
rect 223150 -1424 223218 -1368
rect 223274 -1424 223342 -1368
rect 223398 -1424 240970 -1368
rect 241026 -1424 241094 -1368
rect 241150 -1424 241218 -1368
rect 241274 -1424 241342 -1368
rect 241398 -1424 258970 -1368
rect 259026 -1424 259094 -1368
rect 259150 -1424 259218 -1368
rect 259274 -1424 259342 -1368
rect 259398 -1424 276970 -1368
rect 277026 -1424 277094 -1368
rect 277150 -1424 277218 -1368
rect 277274 -1424 277342 -1368
rect 277398 -1424 294970 -1368
rect 295026 -1424 295094 -1368
rect 295150 -1424 295218 -1368
rect 295274 -1424 295342 -1368
rect 295398 -1424 312970 -1368
rect 313026 -1424 313094 -1368
rect 313150 -1424 313218 -1368
rect 313274 -1424 313342 -1368
rect 313398 -1424 330970 -1368
rect 331026 -1424 331094 -1368
rect 331150 -1424 331218 -1368
rect 331274 -1424 331342 -1368
rect 331398 -1424 348970 -1368
rect 349026 -1424 349094 -1368
rect 349150 -1424 349218 -1368
rect 349274 -1424 349342 -1368
rect 349398 -1424 366970 -1368
rect 367026 -1424 367094 -1368
rect 367150 -1424 367218 -1368
rect 367274 -1424 367342 -1368
rect 367398 -1424 384970 -1368
rect 385026 -1424 385094 -1368
rect 385150 -1424 385218 -1368
rect 385274 -1424 385342 -1368
rect 385398 -1424 402970 -1368
rect 403026 -1424 403094 -1368
rect 403150 -1424 403218 -1368
rect 403274 -1424 403342 -1368
rect 403398 -1424 420970 -1368
rect 421026 -1424 421094 -1368
rect 421150 -1424 421218 -1368
rect 421274 -1424 421342 -1368
rect 421398 -1424 438970 -1368
rect 439026 -1424 439094 -1368
rect 439150 -1424 439218 -1368
rect 439274 -1424 439342 -1368
rect 439398 -1424 456970 -1368
rect 457026 -1424 457094 -1368
rect 457150 -1424 457218 -1368
rect 457274 -1424 457342 -1368
rect 457398 -1424 474970 -1368
rect 475026 -1424 475094 -1368
rect 475150 -1424 475218 -1368
rect 475274 -1424 475342 -1368
rect 475398 -1424 492970 -1368
rect 493026 -1424 493094 -1368
rect 493150 -1424 493218 -1368
rect 493274 -1424 493342 -1368
rect 493398 -1424 510970 -1368
rect 511026 -1424 511094 -1368
rect 511150 -1424 511218 -1368
rect 511274 -1424 511342 -1368
rect 511398 -1424 528970 -1368
rect 529026 -1424 529094 -1368
rect 529150 -1424 529218 -1368
rect 529274 -1424 529342 -1368
rect 529398 -1424 546970 -1368
rect 547026 -1424 547094 -1368
rect 547150 -1424 547218 -1368
rect 547274 -1424 547342 -1368
rect 547398 -1424 564970 -1368
rect 565026 -1424 565094 -1368
rect 565150 -1424 565218 -1368
rect 565274 -1424 565342 -1368
rect 565398 -1424 582970 -1368
rect 583026 -1424 583094 -1368
rect 583150 -1424 583218 -1368
rect 583274 -1424 583342 -1368
rect 583398 -1424 597456 -1368
rect 597512 -1424 597580 -1368
rect 597636 -1424 597704 -1368
rect 597760 -1424 597828 -1368
rect 597884 -1424 597980 -1368
rect -1916 -1492 597980 -1424
rect -1916 -1548 -1820 -1492
rect -1764 -1548 -1696 -1492
rect -1640 -1548 -1572 -1492
rect -1516 -1548 -1448 -1492
rect -1392 -1548 6970 -1492
rect 7026 -1548 7094 -1492
rect 7150 -1548 7218 -1492
rect 7274 -1548 7342 -1492
rect 7398 -1548 24970 -1492
rect 25026 -1548 25094 -1492
rect 25150 -1548 25218 -1492
rect 25274 -1548 25342 -1492
rect 25398 -1548 42970 -1492
rect 43026 -1548 43094 -1492
rect 43150 -1548 43218 -1492
rect 43274 -1548 43342 -1492
rect 43398 -1548 60970 -1492
rect 61026 -1548 61094 -1492
rect 61150 -1548 61218 -1492
rect 61274 -1548 61342 -1492
rect 61398 -1548 78970 -1492
rect 79026 -1548 79094 -1492
rect 79150 -1548 79218 -1492
rect 79274 -1548 79342 -1492
rect 79398 -1548 96970 -1492
rect 97026 -1548 97094 -1492
rect 97150 -1548 97218 -1492
rect 97274 -1548 97342 -1492
rect 97398 -1548 114970 -1492
rect 115026 -1548 115094 -1492
rect 115150 -1548 115218 -1492
rect 115274 -1548 115342 -1492
rect 115398 -1548 132970 -1492
rect 133026 -1548 133094 -1492
rect 133150 -1548 133218 -1492
rect 133274 -1548 133342 -1492
rect 133398 -1548 150970 -1492
rect 151026 -1548 151094 -1492
rect 151150 -1548 151218 -1492
rect 151274 -1548 151342 -1492
rect 151398 -1548 168970 -1492
rect 169026 -1548 169094 -1492
rect 169150 -1548 169218 -1492
rect 169274 -1548 169342 -1492
rect 169398 -1548 186970 -1492
rect 187026 -1548 187094 -1492
rect 187150 -1548 187218 -1492
rect 187274 -1548 187342 -1492
rect 187398 -1548 204970 -1492
rect 205026 -1548 205094 -1492
rect 205150 -1548 205218 -1492
rect 205274 -1548 205342 -1492
rect 205398 -1548 222970 -1492
rect 223026 -1548 223094 -1492
rect 223150 -1548 223218 -1492
rect 223274 -1548 223342 -1492
rect 223398 -1548 240970 -1492
rect 241026 -1548 241094 -1492
rect 241150 -1548 241218 -1492
rect 241274 -1548 241342 -1492
rect 241398 -1548 258970 -1492
rect 259026 -1548 259094 -1492
rect 259150 -1548 259218 -1492
rect 259274 -1548 259342 -1492
rect 259398 -1548 276970 -1492
rect 277026 -1548 277094 -1492
rect 277150 -1548 277218 -1492
rect 277274 -1548 277342 -1492
rect 277398 -1548 294970 -1492
rect 295026 -1548 295094 -1492
rect 295150 -1548 295218 -1492
rect 295274 -1548 295342 -1492
rect 295398 -1548 312970 -1492
rect 313026 -1548 313094 -1492
rect 313150 -1548 313218 -1492
rect 313274 -1548 313342 -1492
rect 313398 -1548 330970 -1492
rect 331026 -1548 331094 -1492
rect 331150 -1548 331218 -1492
rect 331274 -1548 331342 -1492
rect 331398 -1548 348970 -1492
rect 349026 -1548 349094 -1492
rect 349150 -1548 349218 -1492
rect 349274 -1548 349342 -1492
rect 349398 -1548 366970 -1492
rect 367026 -1548 367094 -1492
rect 367150 -1548 367218 -1492
rect 367274 -1548 367342 -1492
rect 367398 -1548 384970 -1492
rect 385026 -1548 385094 -1492
rect 385150 -1548 385218 -1492
rect 385274 -1548 385342 -1492
rect 385398 -1548 402970 -1492
rect 403026 -1548 403094 -1492
rect 403150 -1548 403218 -1492
rect 403274 -1548 403342 -1492
rect 403398 -1548 420970 -1492
rect 421026 -1548 421094 -1492
rect 421150 -1548 421218 -1492
rect 421274 -1548 421342 -1492
rect 421398 -1548 438970 -1492
rect 439026 -1548 439094 -1492
rect 439150 -1548 439218 -1492
rect 439274 -1548 439342 -1492
rect 439398 -1548 456970 -1492
rect 457026 -1548 457094 -1492
rect 457150 -1548 457218 -1492
rect 457274 -1548 457342 -1492
rect 457398 -1548 474970 -1492
rect 475026 -1548 475094 -1492
rect 475150 -1548 475218 -1492
rect 475274 -1548 475342 -1492
rect 475398 -1548 492970 -1492
rect 493026 -1548 493094 -1492
rect 493150 -1548 493218 -1492
rect 493274 -1548 493342 -1492
rect 493398 -1548 510970 -1492
rect 511026 -1548 511094 -1492
rect 511150 -1548 511218 -1492
rect 511274 -1548 511342 -1492
rect 511398 -1548 528970 -1492
rect 529026 -1548 529094 -1492
rect 529150 -1548 529218 -1492
rect 529274 -1548 529342 -1492
rect 529398 -1548 546970 -1492
rect 547026 -1548 547094 -1492
rect 547150 -1548 547218 -1492
rect 547274 -1548 547342 -1492
rect 547398 -1548 564970 -1492
rect 565026 -1548 565094 -1492
rect 565150 -1548 565218 -1492
rect 565274 -1548 565342 -1492
rect 565398 -1548 582970 -1492
rect 583026 -1548 583094 -1492
rect 583150 -1548 583218 -1492
rect 583274 -1548 583342 -1492
rect 583398 -1548 597456 -1492
rect 597512 -1548 597580 -1492
rect 597636 -1548 597704 -1492
rect 597760 -1548 597828 -1492
rect 597884 -1548 597980 -1492
rect -1916 -1644 597980 -1548
use analog_wrapper  analog_wrapper
timestamp 0
transform 1 0 40000 0 1 240000
box 1258 0 508678 350000
use temp_sensor  temp_sensor
timestamp 0
transform 1 0 560000 0 1 380000
box 0 0 28720 120000
use peri_top  u_peri
timestamp 0
transform 1 0 280000 0 1 70000
box 0 0 38640 100000
use pinmux_top  u_pinmux
timestamp 0
transform 1 0 60000 0 1 30000
box 0 0 180000 200000
use uart_i2c_usb_spi_top  u_uart_i2c_usb_spi
timestamp 0
transform 1 0 350000 0 1 40000
box 0 0 200000 180000
use wb_buttons_leds  wb_buttons_leds
timestamp 0
transform 1 0 554000 0 1 10000
box 0 0 40000 50000
<< labels >>
flabel metal3 s 595560 7112 597000 7336 0 FreeSans 896 0 0 0 io_in[0]
port 0 nsew signal input
flabel metal3 s 595560 403592 597000 403816 0 FreeSans 896 0 0 0 io_in[10]
port 1 nsew signal input
flabel metal3 s 595560 443240 597000 443464 0 FreeSans 896 0 0 0 io_in[11]
port 2 nsew signal input
flabel metal3 s 595560 482888 597000 483112 0 FreeSans 896 0 0 0 io_in[12]
port 3 nsew signal input
flabel metal3 s 595560 522536 597000 522760 0 FreeSans 896 0 0 0 io_in[13]
port 4 nsew signal input
flabel metal3 s 595560 562184 597000 562408 0 FreeSans 896 0 0 0 io_in[14]
port 5 nsew signal input
flabel metal2 s 584696 595560 584920 597000 0 FreeSans 896 90 0 0 io_in[15]
port 6 nsew signal input
flabel metal2 s 518504 595560 518728 597000 0 FreeSans 896 90 0 0 io_in[16]
port 7 nsew signal input
flabel metal2 s 452312 595560 452536 597000 0 FreeSans 896 90 0 0 io_in[17]
port 8 nsew signal input
flabel metal2 s 386120 595560 386344 597000 0 FreeSans 896 90 0 0 io_in[18]
port 9 nsew signal input
flabel metal2 s 319928 595560 320152 597000 0 FreeSans 896 90 0 0 io_in[19]
port 10 nsew signal input
flabel metal3 s 595560 46760 597000 46984 0 FreeSans 896 0 0 0 io_in[1]
port 11 nsew signal input
flabel metal2 s 253736 595560 253960 597000 0 FreeSans 896 90 0 0 io_in[20]
port 12 nsew signal input
flabel metal2 s 187544 595560 187768 597000 0 FreeSans 896 90 0 0 io_in[21]
port 13 nsew signal input
flabel metal2 s 121352 595560 121576 597000 0 FreeSans 896 90 0 0 io_in[22]
port 14 nsew signal input
flabel metal2 s 55160 595560 55384 597000 0 FreeSans 896 90 0 0 io_in[23]
port 15 nsew signal input
flabel metal3 s -960 587160 480 587384 0 FreeSans 896 0 0 0 io_in[24]
port 16 nsew signal input
flabel metal3 s -960 544824 480 545048 0 FreeSans 896 0 0 0 io_in[25]
port 17 nsew signal input
flabel metal3 s -960 502488 480 502712 0 FreeSans 896 0 0 0 io_in[26]
port 18 nsew signal input
flabel metal3 s -960 460152 480 460376 0 FreeSans 896 0 0 0 io_in[27]
port 19 nsew signal input
flabel metal3 s -960 417816 480 418040 0 FreeSans 896 0 0 0 io_in[28]
port 20 nsew signal input
flabel metal3 s -960 375480 480 375704 0 FreeSans 896 0 0 0 io_in[29]
port 21 nsew signal input
flabel metal3 s 595560 86408 597000 86632 0 FreeSans 896 0 0 0 io_in[2]
port 22 nsew signal input
flabel metal3 s -960 333144 480 333368 0 FreeSans 896 0 0 0 io_in[30]
port 23 nsew signal input
flabel metal3 s -960 290808 480 291032 0 FreeSans 896 0 0 0 io_in[31]
port 24 nsew signal input
flabel metal3 s -960 248472 480 248696 0 FreeSans 896 0 0 0 io_in[32]
port 25 nsew signal input
flabel metal3 s -960 206136 480 206360 0 FreeSans 896 0 0 0 io_in[33]
port 26 nsew signal input
flabel metal3 s -960 163800 480 164024 0 FreeSans 896 0 0 0 io_in[34]
port 27 nsew signal input
flabel metal3 s -960 121464 480 121688 0 FreeSans 896 0 0 0 io_in[35]
port 28 nsew signal input
flabel metal3 s -960 79128 480 79352 0 FreeSans 896 0 0 0 io_in[36]
port 29 nsew signal input
flabel metal3 s -960 36792 480 37016 0 FreeSans 896 0 0 0 io_in[37]
port 30 nsew signal input
flabel metal3 s 595560 126056 597000 126280 0 FreeSans 896 0 0 0 io_in[3]
port 31 nsew signal input
flabel metal3 s 595560 165704 597000 165928 0 FreeSans 896 0 0 0 io_in[4]
port 32 nsew signal input
flabel metal3 s 595560 205352 597000 205576 0 FreeSans 896 0 0 0 io_in[5]
port 33 nsew signal input
flabel metal3 s 595560 245000 597000 245224 0 FreeSans 896 0 0 0 io_in[6]
port 34 nsew signal input
flabel metal3 s 595560 284648 597000 284872 0 FreeSans 896 0 0 0 io_in[7]
port 35 nsew signal input
flabel metal3 s 595560 324296 597000 324520 0 FreeSans 896 0 0 0 io_in[8]
port 36 nsew signal input
flabel metal3 s 595560 363944 597000 364168 0 FreeSans 896 0 0 0 io_in[9]
port 37 nsew signal input
flabel metal3 s 595560 33544 597000 33768 0 FreeSans 896 0 0 0 io_oeb[0]
port 38 nsew signal tristate
flabel metal3 s 595560 430024 597000 430248 0 FreeSans 896 0 0 0 io_oeb[10]
port 39 nsew signal tristate
flabel metal3 s 595560 469672 597000 469896 0 FreeSans 896 0 0 0 io_oeb[11]
port 40 nsew signal tristate
flabel metal3 s 595560 509320 597000 509544 0 FreeSans 896 0 0 0 io_oeb[12]
port 41 nsew signal tristate
flabel metal3 s 595560 548968 597000 549192 0 FreeSans 896 0 0 0 io_oeb[13]
port 42 nsew signal tristate
flabel metal3 s 595560 588616 597000 588840 0 FreeSans 896 0 0 0 io_oeb[14]
port 43 nsew signal tristate
flabel metal2 s 540568 595560 540792 597000 0 FreeSans 896 90 0 0 io_oeb[15]
port 44 nsew signal tristate
flabel metal2 s 474376 595560 474600 597000 0 FreeSans 896 90 0 0 io_oeb[16]
port 45 nsew signal tristate
flabel metal2 s 408184 595560 408408 597000 0 FreeSans 896 90 0 0 io_oeb[17]
port 46 nsew signal tristate
flabel metal2 s 341992 595560 342216 597000 0 FreeSans 896 90 0 0 io_oeb[18]
port 47 nsew signal tristate
flabel metal2 s 275800 595560 276024 597000 0 FreeSans 896 90 0 0 io_oeb[19]
port 48 nsew signal tristate
flabel metal3 s 595560 73192 597000 73416 0 FreeSans 896 0 0 0 io_oeb[1]
port 49 nsew signal tristate
flabel metal2 s 209608 595560 209832 597000 0 FreeSans 896 90 0 0 io_oeb[20]
port 50 nsew signal tristate
flabel metal2 s 143416 595560 143640 597000 0 FreeSans 896 90 0 0 io_oeb[21]
port 51 nsew signal tristate
flabel metal2 s 77224 595560 77448 597000 0 FreeSans 896 90 0 0 io_oeb[22]
port 52 nsew signal tristate
flabel metal2 s 11032 595560 11256 597000 0 FreeSans 896 90 0 0 io_oeb[23]
port 53 nsew signal tristate
flabel metal3 s -960 558936 480 559160 0 FreeSans 896 0 0 0 io_oeb[24]
port 54 nsew signal tristate
flabel metal3 s -960 516600 480 516824 0 FreeSans 896 0 0 0 io_oeb[25]
port 55 nsew signal tristate
flabel metal3 s -960 474264 480 474488 0 FreeSans 896 0 0 0 io_oeb[26]
port 56 nsew signal tristate
flabel metal3 s -960 431928 480 432152 0 FreeSans 896 0 0 0 io_oeb[27]
port 57 nsew signal tristate
flabel metal3 s -960 389592 480 389816 0 FreeSans 896 0 0 0 io_oeb[28]
port 58 nsew signal tristate
flabel metal3 s -960 347256 480 347480 0 FreeSans 896 0 0 0 io_oeb[29]
port 59 nsew signal tristate
flabel metal3 s 595560 112840 597000 113064 0 FreeSans 896 0 0 0 io_oeb[2]
port 60 nsew signal tristate
flabel metal3 s -960 304920 480 305144 0 FreeSans 896 0 0 0 io_oeb[30]
port 61 nsew signal tristate
flabel metal3 s -960 262584 480 262808 0 FreeSans 896 0 0 0 io_oeb[31]
port 62 nsew signal tristate
flabel metal3 s -960 220248 480 220472 0 FreeSans 896 0 0 0 io_oeb[32]
port 63 nsew signal tristate
flabel metal3 s -960 177912 480 178136 0 FreeSans 896 0 0 0 io_oeb[33]
port 64 nsew signal tristate
flabel metal3 s -960 135576 480 135800 0 FreeSans 896 0 0 0 io_oeb[34]
port 65 nsew signal tristate
flabel metal3 s -960 93240 480 93464 0 FreeSans 896 0 0 0 io_oeb[35]
port 66 nsew signal tristate
flabel metal3 s -960 50904 480 51128 0 FreeSans 896 0 0 0 io_oeb[36]
port 67 nsew signal tristate
flabel metal3 s -960 8568 480 8792 0 FreeSans 896 0 0 0 io_oeb[37]
port 68 nsew signal tristate
flabel metal3 s 595560 152488 597000 152712 0 FreeSans 896 0 0 0 io_oeb[3]
port 69 nsew signal tristate
flabel metal3 s 595560 192136 597000 192360 0 FreeSans 896 0 0 0 io_oeb[4]
port 70 nsew signal tristate
flabel metal3 s 595560 231784 597000 232008 0 FreeSans 896 0 0 0 io_oeb[5]
port 71 nsew signal tristate
flabel metal3 s 595560 271432 597000 271656 0 FreeSans 896 0 0 0 io_oeb[6]
port 72 nsew signal tristate
flabel metal3 s 595560 311080 597000 311304 0 FreeSans 896 0 0 0 io_oeb[7]
port 73 nsew signal tristate
flabel metal3 s 595560 350728 597000 350952 0 FreeSans 896 0 0 0 io_oeb[8]
port 74 nsew signal tristate
flabel metal3 s 595560 390376 597000 390600 0 FreeSans 896 0 0 0 io_oeb[9]
port 75 nsew signal tristate
flabel metal3 s 595560 20328 597000 20552 0 FreeSans 896 0 0 0 io_out[0]
port 76 nsew signal tristate
flabel metal3 s 595560 416808 597000 417032 0 FreeSans 896 0 0 0 io_out[10]
port 77 nsew signal tristate
flabel metal3 s 595560 456456 597000 456680 0 FreeSans 896 0 0 0 io_out[11]
port 78 nsew signal tristate
flabel metal3 s 595560 496104 597000 496328 0 FreeSans 896 0 0 0 io_out[12]
port 79 nsew signal tristate
flabel metal3 s 595560 535752 597000 535976 0 FreeSans 896 0 0 0 io_out[13]
port 80 nsew signal tristate
flabel metal3 s 595560 575400 597000 575624 0 FreeSans 896 0 0 0 io_out[14]
port 81 nsew signal tristate
flabel metal2 s 562632 595560 562856 597000 0 FreeSans 896 90 0 0 io_out[15]
port 82 nsew signal tristate
flabel metal2 s 496440 595560 496664 597000 0 FreeSans 896 90 0 0 io_out[16]
port 83 nsew signal tristate
flabel metal2 s 430248 595560 430472 597000 0 FreeSans 896 90 0 0 io_out[17]
port 84 nsew signal tristate
flabel metal2 s 364056 595560 364280 597000 0 FreeSans 896 90 0 0 io_out[18]
port 85 nsew signal tristate
flabel metal2 s 297864 595560 298088 597000 0 FreeSans 896 90 0 0 io_out[19]
port 86 nsew signal tristate
flabel metal3 s 595560 59976 597000 60200 0 FreeSans 896 0 0 0 io_out[1]
port 87 nsew signal tristate
flabel metal2 s 231672 595560 231896 597000 0 FreeSans 896 90 0 0 io_out[20]
port 88 nsew signal tristate
flabel metal2 s 165480 595560 165704 597000 0 FreeSans 896 90 0 0 io_out[21]
port 89 nsew signal tristate
flabel metal2 s 99288 595560 99512 597000 0 FreeSans 896 90 0 0 io_out[22]
port 90 nsew signal tristate
flabel metal2 s 33096 595560 33320 597000 0 FreeSans 896 90 0 0 io_out[23]
port 91 nsew signal tristate
flabel metal3 s -960 573048 480 573272 0 FreeSans 896 0 0 0 io_out[24]
port 92 nsew signal tristate
flabel metal3 s -960 530712 480 530936 0 FreeSans 896 0 0 0 io_out[25]
port 93 nsew signal tristate
flabel metal3 s -960 488376 480 488600 0 FreeSans 896 0 0 0 io_out[26]
port 94 nsew signal tristate
flabel metal3 s -960 446040 480 446264 0 FreeSans 896 0 0 0 io_out[27]
port 95 nsew signal tristate
flabel metal3 s -960 403704 480 403928 0 FreeSans 896 0 0 0 io_out[28]
port 96 nsew signal tristate
flabel metal3 s -960 361368 480 361592 0 FreeSans 896 0 0 0 io_out[29]
port 97 nsew signal tristate
flabel metal3 s 595560 99624 597000 99848 0 FreeSans 896 0 0 0 io_out[2]
port 98 nsew signal tristate
flabel metal3 s -960 319032 480 319256 0 FreeSans 896 0 0 0 io_out[30]
port 99 nsew signal tristate
flabel metal3 s -960 276696 480 276920 0 FreeSans 896 0 0 0 io_out[31]
port 100 nsew signal tristate
flabel metal3 s -960 234360 480 234584 0 FreeSans 896 0 0 0 io_out[32]
port 101 nsew signal tristate
flabel metal3 s -960 192024 480 192248 0 FreeSans 896 0 0 0 io_out[33]
port 102 nsew signal tristate
flabel metal3 s -960 149688 480 149912 0 FreeSans 896 0 0 0 io_out[34]
port 103 nsew signal tristate
flabel metal3 s -960 107352 480 107576 0 FreeSans 896 0 0 0 io_out[35]
port 104 nsew signal tristate
flabel metal3 s -960 65016 480 65240 0 FreeSans 896 0 0 0 io_out[36]
port 105 nsew signal tristate
flabel metal3 s -960 22680 480 22904 0 FreeSans 896 0 0 0 io_out[37]
port 106 nsew signal tristate
flabel metal3 s 595560 139272 597000 139496 0 FreeSans 896 0 0 0 io_out[3]
port 107 nsew signal tristate
flabel metal3 s 595560 178920 597000 179144 0 FreeSans 896 0 0 0 io_out[4]
port 108 nsew signal tristate
flabel metal3 s 595560 218568 597000 218792 0 FreeSans 896 0 0 0 io_out[5]
port 109 nsew signal tristate
flabel metal3 s 595560 258216 597000 258440 0 FreeSans 896 0 0 0 io_out[6]
port 110 nsew signal tristate
flabel metal3 s 595560 297864 597000 298088 0 FreeSans 896 0 0 0 io_out[7]
port 111 nsew signal tristate
flabel metal3 s 595560 337512 597000 337736 0 FreeSans 896 0 0 0 io_out[8]
port 112 nsew signal tristate
flabel metal3 s 595560 377160 597000 377384 0 FreeSans 896 0 0 0 io_out[9]
port 113 nsew signal tristate
flabel metal2 s 213192 -960 213416 480 0 FreeSans 896 90 0 0 la_data_in[0]
port 114 nsew signal input
flabel metal2 s 270312 -960 270536 480 0 FreeSans 896 90 0 0 la_data_in[10]
port 115 nsew signal input
flabel metal2 s 276024 -960 276248 480 0 FreeSans 896 90 0 0 la_data_in[11]
port 116 nsew signal input
flabel metal2 s 281736 -960 281960 480 0 FreeSans 896 90 0 0 la_data_in[12]
port 117 nsew signal input
flabel metal2 s 287448 -960 287672 480 0 FreeSans 896 90 0 0 la_data_in[13]
port 118 nsew signal input
flabel metal2 s 293160 -960 293384 480 0 FreeSans 896 90 0 0 la_data_in[14]
port 119 nsew signal input
flabel metal2 s 298872 -960 299096 480 0 FreeSans 896 90 0 0 la_data_in[15]
port 120 nsew signal input
flabel metal2 s 304584 -960 304808 480 0 FreeSans 896 90 0 0 la_data_in[16]
port 121 nsew signal input
flabel metal2 s 310296 -960 310520 480 0 FreeSans 896 90 0 0 la_data_in[17]
port 122 nsew signal input
flabel metal2 s 316008 -960 316232 480 0 FreeSans 896 90 0 0 la_data_in[18]
port 123 nsew signal input
flabel metal2 s 321720 -960 321944 480 0 FreeSans 896 90 0 0 la_data_in[19]
port 124 nsew signal input
flabel metal2 s 218904 -960 219128 480 0 FreeSans 896 90 0 0 la_data_in[1]
port 125 nsew signal input
flabel metal2 s 327432 -960 327656 480 0 FreeSans 896 90 0 0 la_data_in[20]
port 126 nsew signal input
flabel metal2 s 333144 -960 333368 480 0 FreeSans 896 90 0 0 la_data_in[21]
port 127 nsew signal input
flabel metal2 s 338856 -960 339080 480 0 FreeSans 896 90 0 0 la_data_in[22]
port 128 nsew signal input
flabel metal2 s 344568 -960 344792 480 0 FreeSans 896 90 0 0 la_data_in[23]
port 129 nsew signal input
flabel metal2 s 350280 -960 350504 480 0 FreeSans 896 90 0 0 la_data_in[24]
port 130 nsew signal input
flabel metal2 s 355992 -960 356216 480 0 FreeSans 896 90 0 0 la_data_in[25]
port 131 nsew signal input
flabel metal2 s 361704 -960 361928 480 0 FreeSans 896 90 0 0 la_data_in[26]
port 132 nsew signal input
flabel metal2 s 367416 -960 367640 480 0 FreeSans 896 90 0 0 la_data_in[27]
port 133 nsew signal input
flabel metal2 s 373128 -960 373352 480 0 FreeSans 896 90 0 0 la_data_in[28]
port 134 nsew signal input
flabel metal2 s 378840 -960 379064 480 0 FreeSans 896 90 0 0 la_data_in[29]
port 135 nsew signal input
flabel metal2 s 224616 -960 224840 480 0 FreeSans 896 90 0 0 la_data_in[2]
port 136 nsew signal input
flabel metal2 s 384552 -960 384776 480 0 FreeSans 896 90 0 0 la_data_in[30]
port 137 nsew signal input
flabel metal2 s 390264 -960 390488 480 0 FreeSans 896 90 0 0 la_data_in[31]
port 138 nsew signal input
flabel metal2 s 395976 -960 396200 480 0 FreeSans 896 90 0 0 la_data_in[32]
port 139 nsew signal input
flabel metal2 s 401688 -960 401912 480 0 FreeSans 896 90 0 0 la_data_in[33]
port 140 nsew signal input
flabel metal2 s 407400 -960 407624 480 0 FreeSans 896 90 0 0 la_data_in[34]
port 141 nsew signal input
flabel metal2 s 413112 -960 413336 480 0 FreeSans 896 90 0 0 la_data_in[35]
port 142 nsew signal input
flabel metal2 s 418824 -960 419048 480 0 FreeSans 896 90 0 0 la_data_in[36]
port 143 nsew signal input
flabel metal2 s 424536 -960 424760 480 0 FreeSans 896 90 0 0 la_data_in[37]
port 144 nsew signal input
flabel metal2 s 430248 -960 430472 480 0 FreeSans 896 90 0 0 la_data_in[38]
port 145 nsew signal input
flabel metal2 s 435960 -960 436184 480 0 FreeSans 896 90 0 0 la_data_in[39]
port 146 nsew signal input
flabel metal2 s 230328 -960 230552 480 0 FreeSans 896 90 0 0 la_data_in[3]
port 147 nsew signal input
flabel metal2 s 441672 -960 441896 480 0 FreeSans 896 90 0 0 la_data_in[40]
port 148 nsew signal input
flabel metal2 s 447384 -960 447608 480 0 FreeSans 896 90 0 0 la_data_in[41]
port 149 nsew signal input
flabel metal2 s 453096 -960 453320 480 0 FreeSans 896 90 0 0 la_data_in[42]
port 150 nsew signal input
flabel metal2 s 458808 -960 459032 480 0 FreeSans 896 90 0 0 la_data_in[43]
port 151 nsew signal input
flabel metal2 s 464520 -960 464744 480 0 FreeSans 896 90 0 0 la_data_in[44]
port 152 nsew signal input
flabel metal2 s 470232 -960 470456 480 0 FreeSans 896 90 0 0 la_data_in[45]
port 153 nsew signal input
flabel metal2 s 475944 -960 476168 480 0 FreeSans 896 90 0 0 la_data_in[46]
port 154 nsew signal input
flabel metal2 s 481656 -960 481880 480 0 FreeSans 896 90 0 0 la_data_in[47]
port 155 nsew signal input
flabel metal2 s 487368 -960 487592 480 0 FreeSans 896 90 0 0 la_data_in[48]
port 156 nsew signal input
flabel metal2 s 493080 -960 493304 480 0 FreeSans 896 90 0 0 la_data_in[49]
port 157 nsew signal input
flabel metal2 s 236040 -960 236264 480 0 FreeSans 896 90 0 0 la_data_in[4]
port 158 nsew signal input
flabel metal2 s 498792 -960 499016 480 0 FreeSans 896 90 0 0 la_data_in[50]
port 159 nsew signal input
flabel metal2 s 504504 -960 504728 480 0 FreeSans 896 90 0 0 la_data_in[51]
port 160 nsew signal input
flabel metal2 s 510216 -960 510440 480 0 FreeSans 896 90 0 0 la_data_in[52]
port 161 nsew signal input
flabel metal2 s 515928 -960 516152 480 0 FreeSans 896 90 0 0 la_data_in[53]
port 162 nsew signal input
flabel metal2 s 521640 -960 521864 480 0 FreeSans 896 90 0 0 la_data_in[54]
port 163 nsew signal input
flabel metal2 s 527352 -960 527576 480 0 FreeSans 896 90 0 0 la_data_in[55]
port 164 nsew signal input
flabel metal2 s 533064 -960 533288 480 0 FreeSans 896 90 0 0 la_data_in[56]
port 165 nsew signal input
flabel metal2 s 538776 -960 539000 480 0 FreeSans 896 90 0 0 la_data_in[57]
port 166 nsew signal input
flabel metal2 s 544488 -960 544712 480 0 FreeSans 896 90 0 0 la_data_in[58]
port 167 nsew signal input
flabel metal2 s 550200 -960 550424 480 0 FreeSans 896 90 0 0 la_data_in[59]
port 168 nsew signal input
flabel metal2 s 241752 -960 241976 480 0 FreeSans 896 90 0 0 la_data_in[5]
port 169 nsew signal input
flabel metal2 s 555912 -960 556136 480 0 FreeSans 896 90 0 0 la_data_in[60]
port 170 nsew signal input
flabel metal2 s 561624 -960 561848 480 0 FreeSans 896 90 0 0 la_data_in[61]
port 171 nsew signal input
flabel metal2 s 567336 -960 567560 480 0 FreeSans 896 90 0 0 la_data_in[62]
port 172 nsew signal input
flabel metal2 s 573048 -960 573272 480 0 FreeSans 896 90 0 0 la_data_in[63]
port 173 nsew signal input
flabel metal2 s 247464 -960 247688 480 0 FreeSans 896 90 0 0 la_data_in[6]
port 174 nsew signal input
flabel metal2 s 253176 -960 253400 480 0 FreeSans 896 90 0 0 la_data_in[7]
port 175 nsew signal input
flabel metal2 s 258888 -960 259112 480 0 FreeSans 896 90 0 0 la_data_in[8]
port 176 nsew signal input
flabel metal2 s 264600 -960 264824 480 0 FreeSans 896 90 0 0 la_data_in[9]
port 177 nsew signal input
flabel metal2 s 215096 -960 215320 480 0 FreeSans 896 90 0 0 la_data_out[0]
port 178 nsew signal tristate
flabel metal2 s 272216 -960 272440 480 0 FreeSans 896 90 0 0 la_data_out[10]
port 179 nsew signal tristate
flabel metal2 s 277928 -960 278152 480 0 FreeSans 896 90 0 0 la_data_out[11]
port 180 nsew signal tristate
flabel metal2 s 283640 -960 283864 480 0 FreeSans 896 90 0 0 la_data_out[12]
port 181 nsew signal tristate
flabel metal2 s 289352 -960 289576 480 0 FreeSans 896 90 0 0 la_data_out[13]
port 182 nsew signal tristate
flabel metal2 s 295064 -960 295288 480 0 FreeSans 896 90 0 0 la_data_out[14]
port 183 nsew signal tristate
flabel metal2 s 300776 -960 301000 480 0 FreeSans 896 90 0 0 la_data_out[15]
port 184 nsew signal tristate
flabel metal2 s 306488 -960 306712 480 0 FreeSans 896 90 0 0 la_data_out[16]
port 185 nsew signal tristate
flabel metal2 s 312200 -960 312424 480 0 FreeSans 896 90 0 0 la_data_out[17]
port 186 nsew signal tristate
flabel metal2 s 317912 -960 318136 480 0 FreeSans 896 90 0 0 la_data_out[18]
port 187 nsew signal tristate
flabel metal2 s 323624 -960 323848 480 0 FreeSans 896 90 0 0 la_data_out[19]
port 188 nsew signal tristate
flabel metal2 s 220808 -960 221032 480 0 FreeSans 896 90 0 0 la_data_out[1]
port 189 nsew signal tristate
flabel metal2 s 329336 -960 329560 480 0 FreeSans 896 90 0 0 la_data_out[20]
port 190 nsew signal tristate
flabel metal2 s 335048 -960 335272 480 0 FreeSans 896 90 0 0 la_data_out[21]
port 191 nsew signal tristate
flabel metal2 s 340760 -960 340984 480 0 FreeSans 896 90 0 0 la_data_out[22]
port 192 nsew signal tristate
flabel metal2 s 346472 -960 346696 480 0 FreeSans 896 90 0 0 la_data_out[23]
port 193 nsew signal tristate
flabel metal2 s 352184 -960 352408 480 0 FreeSans 896 90 0 0 la_data_out[24]
port 194 nsew signal tristate
flabel metal2 s 357896 -960 358120 480 0 FreeSans 896 90 0 0 la_data_out[25]
port 195 nsew signal tristate
flabel metal2 s 363608 -960 363832 480 0 FreeSans 896 90 0 0 la_data_out[26]
port 196 nsew signal tristate
flabel metal2 s 369320 -960 369544 480 0 FreeSans 896 90 0 0 la_data_out[27]
port 197 nsew signal tristate
flabel metal2 s 375032 -960 375256 480 0 FreeSans 896 90 0 0 la_data_out[28]
port 198 nsew signal tristate
flabel metal2 s 380744 -960 380968 480 0 FreeSans 896 90 0 0 la_data_out[29]
port 199 nsew signal tristate
flabel metal2 s 226520 -960 226744 480 0 FreeSans 896 90 0 0 la_data_out[2]
port 200 nsew signal tristate
flabel metal2 s 386456 -960 386680 480 0 FreeSans 896 90 0 0 la_data_out[30]
port 201 nsew signal tristate
flabel metal2 s 392168 -960 392392 480 0 FreeSans 896 90 0 0 la_data_out[31]
port 202 nsew signal tristate
flabel metal2 s 397880 -960 398104 480 0 FreeSans 896 90 0 0 la_data_out[32]
port 203 nsew signal tristate
flabel metal2 s 403592 -960 403816 480 0 FreeSans 896 90 0 0 la_data_out[33]
port 204 nsew signal tristate
flabel metal2 s 409304 -960 409528 480 0 FreeSans 896 90 0 0 la_data_out[34]
port 205 nsew signal tristate
flabel metal2 s 415016 -960 415240 480 0 FreeSans 896 90 0 0 la_data_out[35]
port 206 nsew signal tristate
flabel metal2 s 420728 -960 420952 480 0 FreeSans 896 90 0 0 la_data_out[36]
port 207 nsew signal tristate
flabel metal2 s 426440 -960 426664 480 0 FreeSans 896 90 0 0 la_data_out[37]
port 208 nsew signal tristate
flabel metal2 s 432152 -960 432376 480 0 FreeSans 896 90 0 0 la_data_out[38]
port 209 nsew signal tristate
flabel metal2 s 437864 -960 438088 480 0 FreeSans 896 90 0 0 la_data_out[39]
port 210 nsew signal tristate
flabel metal2 s 232232 -960 232456 480 0 FreeSans 896 90 0 0 la_data_out[3]
port 211 nsew signal tristate
flabel metal2 s 443576 -960 443800 480 0 FreeSans 896 90 0 0 la_data_out[40]
port 212 nsew signal tristate
flabel metal2 s 449288 -960 449512 480 0 FreeSans 896 90 0 0 la_data_out[41]
port 213 nsew signal tristate
flabel metal2 s 455000 -960 455224 480 0 FreeSans 896 90 0 0 la_data_out[42]
port 214 nsew signal tristate
flabel metal2 s 460712 -960 460936 480 0 FreeSans 896 90 0 0 la_data_out[43]
port 215 nsew signal tristate
flabel metal2 s 466424 -960 466648 480 0 FreeSans 896 90 0 0 la_data_out[44]
port 216 nsew signal tristate
flabel metal2 s 472136 -960 472360 480 0 FreeSans 896 90 0 0 la_data_out[45]
port 217 nsew signal tristate
flabel metal2 s 477848 -960 478072 480 0 FreeSans 896 90 0 0 la_data_out[46]
port 218 nsew signal tristate
flabel metal2 s 483560 -960 483784 480 0 FreeSans 896 90 0 0 la_data_out[47]
port 219 nsew signal tristate
flabel metal2 s 489272 -960 489496 480 0 FreeSans 896 90 0 0 la_data_out[48]
port 220 nsew signal tristate
flabel metal2 s 494984 -960 495208 480 0 FreeSans 896 90 0 0 la_data_out[49]
port 221 nsew signal tristate
flabel metal2 s 237944 -960 238168 480 0 FreeSans 896 90 0 0 la_data_out[4]
port 222 nsew signal tristate
flabel metal2 s 500696 -960 500920 480 0 FreeSans 896 90 0 0 la_data_out[50]
port 223 nsew signal tristate
flabel metal2 s 506408 -960 506632 480 0 FreeSans 896 90 0 0 la_data_out[51]
port 224 nsew signal tristate
flabel metal2 s 512120 -960 512344 480 0 FreeSans 896 90 0 0 la_data_out[52]
port 225 nsew signal tristate
flabel metal2 s 517832 -960 518056 480 0 FreeSans 896 90 0 0 la_data_out[53]
port 226 nsew signal tristate
flabel metal2 s 523544 -960 523768 480 0 FreeSans 896 90 0 0 la_data_out[54]
port 227 nsew signal tristate
flabel metal2 s 529256 -960 529480 480 0 FreeSans 896 90 0 0 la_data_out[55]
port 228 nsew signal tristate
flabel metal2 s 534968 -960 535192 480 0 FreeSans 896 90 0 0 la_data_out[56]
port 229 nsew signal tristate
flabel metal2 s 540680 -960 540904 480 0 FreeSans 896 90 0 0 la_data_out[57]
port 230 nsew signal tristate
flabel metal2 s 546392 -960 546616 480 0 FreeSans 896 90 0 0 la_data_out[58]
port 231 nsew signal tristate
flabel metal2 s 552104 -960 552328 480 0 FreeSans 896 90 0 0 la_data_out[59]
port 232 nsew signal tristate
flabel metal2 s 243656 -960 243880 480 0 FreeSans 896 90 0 0 la_data_out[5]
port 233 nsew signal tristate
flabel metal2 s 557816 -960 558040 480 0 FreeSans 896 90 0 0 la_data_out[60]
port 234 nsew signal tristate
flabel metal2 s 563528 -960 563752 480 0 FreeSans 896 90 0 0 la_data_out[61]
port 235 nsew signal tristate
flabel metal2 s 569240 -960 569464 480 0 FreeSans 896 90 0 0 la_data_out[62]
port 236 nsew signal tristate
flabel metal2 s 574952 -960 575176 480 0 FreeSans 896 90 0 0 la_data_out[63]
port 237 nsew signal tristate
flabel metal2 s 249368 -960 249592 480 0 FreeSans 896 90 0 0 la_data_out[6]
port 238 nsew signal tristate
flabel metal2 s 255080 -960 255304 480 0 FreeSans 896 90 0 0 la_data_out[7]
port 239 nsew signal tristate
flabel metal2 s 260792 -960 261016 480 0 FreeSans 896 90 0 0 la_data_out[8]
port 240 nsew signal tristate
flabel metal2 s 266504 -960 266728 480 0 FreeSans 896 90 0 0 la_data_out[9]
port 241 nsew signal tristate
flabel metal2 s 217000 -960 217224 480 0 FreeSans 896 90 0 0 la_oenb[0]
port 242 nsew signal input
flabel metal2 s 274120 -960 274344 480 0 FreeSans 896 90 0 0 la_oenb[10]
port 243 nsew signal input
flabel metal2 s 279832 -960 280056 480 0 FreeSans 896 90 0 0 la_oenb[11]
port 244 nsew signal input
flabel metal2 s 285544 -960 285768 480 0 FreeSans 896 90 0 0 la_oenb[12]
port 245 nsew signal input
flabel metal2 s 291256 -960 291480 480 0 FreeSans 896 90 0 0 la_oenb[13]
port 246 nsew signal input
flabel metal2 s 296968 -960 297192 480 0 FreeSans 896 90 0 0 la_oenb[14]
port 247 nsew signal input
flabel metal2 s 302680 -960 302904 480 0 FreeSans 896 90 0 0 la_oenb[15]
port 248 nsew signal input
flabel metal2 s 308392 -960 308616 480 0 FreeSans 896 90 0 0 la_oenb[16]
port 249 nsew signal input
flabel metal2 s 314104 -960 314328 480 0 FreeSans 896 90 0 0 la_oenb[17]
port 250 nsew signal input
flabel metal2 s 319816 -960 320040 480 0 FreeSans 896 90 0 0 la_oenb[18]
port 251 nsew signal input
flabel metal2 s 325528 -960 325752 480 0 FreeSans 896 90 0 0 la_oenb[19]
port 252 nsew signal input
flabel metal2 s 222712 -960 222936 480 0 FreeSans 896 90 0 0 la_oenb[1]
port 253 nsew signal input
flabel metal2 s 331240 -960 331464 480 0 FreeSans 896 90 0 0 la_oenb[20]
port 254 nsew signal input
flabel metal2 s 336952 -960 337176 480 0 FreeSans 896 90 0 0 la_oenb[21]
port 255 nsew signal input
flabel metal2 s 342664 -960 342888 480 0 FreeSans 896 90 0 0 la_oenb[22]
port 256 nsew signal input
flabel metal2 s 348376 -960 348600 480 0 FreeSans 896 90 0 0 la_oenb[23]
port 257 nsew signal input
flabel metal2 s 354088 -960 354312 480 0 FreeSans 896 90 0 0 la_oenb[24]
port 258 nsew signal input
flabel metal2 s 359800 -960 360024 480 0 FreeSans 896 90 0 0 la_oenb[25]
port 259 nsew signal input
flabel metal2 s 365512 -960 365736 480 0 FreeSans 896 90 0 0 la_oenb[26]
port 260 nsew signal input
flabel metal2 s 371224 -960 371448 480 0 FreeSans 896 90 0 0 la_oenb[27]
port 261 nsew signal input
flabel metal2 s 376936 -960 377160 480 0 FreeSans 896 90 0 0 la_oenb[28]
port 262 nsew signal input
flabel metal2 s 382648 -960 382872 480 0 FreeSans 896 90 0 0 la_oenb[29]
port 263 nsew signal input
flabel metal2 s 228424 -960 228648 480 0 FreeSans 896 90 0 0 la_oenb[2]
port 264 nsew signal input
flabel metal2 s 388360 -960 388584 480 0 FreeSans 896 90 0 0 la_oenb[30]
port 265 nsew signal input
flabel metal2 s 394072 -960 394296 480 0 FreeSans 896 90 0 0 la_oenb[31]
port 266 nsew signal input
flabel metal2 s 399784 -960 400008 480 0 FreeSans 896 90 0 0 la_oenb[32]
port 267 nsew signal input
flabel metal2 s 405496 -960 405720 480 0 FreeSans 896 90 0 0 la_oenb[33]
port 268 nsew signal input
flabel metal2 s 411208 -960 411432 480 0 FreeSans 896 90 0 0 la_oenb[34]
port 269 nsew signal input
flabel metal2 s 416920 -960 417144 480 0 FreeSans 896 90 0 0 la_oenb[35]
port 270 nsew signal input
flabel metal2 s 422632 -960 422856 480 0 FreeSans 896 90 0 0 la_oenb[36]
port 271 nsew signal input
flabel metal2 s 428344 -960 428568 480 0 FreeSans 896 90 0 0 la_oenb[37]
port 272 nsew signal input
flabel metal2 s 434056 -960 434280 480 0 FreeSans 896 90 0 0 la_oenb[38]
port 273 nsew signal input
flabel metal2 s 439768 -960 439992 480 0 FreeSans 896 90 0 0 la_oenb[39]
port 274 nsew signal input
flabel metal2 s 234136 -960 234360 480 0 FreeSans 896 90 0 0 la_oenb[3]
port 275 nsew signal input
flabel metal2 s 445480 -960 445704 480 0 FreeSans 896 90 0 0 la_oenb[40]
port 276 nsew signal input
flabel metal2 s 451192 -960 451416 480 0 FreeSans 896 90 0 0 la_oenb[41]
port 277 nsew signal input
flabel metal2 s 456904 -960 457128 480 0 FreeSans 896 90 0 0 la_oenb[42]
port 278 nsew signal input
flabel metal2 s 462616 -960 462840 480 0 FreeSans 896 90 0 0 la_oenb[43]
port 279 nsew signal input
flabel metal2 s 468328 -960 468552 480 0 FreeSans 896 90 0 0 la_oenb[44]
port 280 nsew signal input
flabel metal2 s 474040 -960 474264 480 0 FreeSans 896 90 0 0 la_oenb[45]
port 281 nsew signal input
flabel metal2 s 479752 -960 479976 480 0 FreeSans 896 90 0 0 la_oenb[46]
port 282 nsew signal input
flabel metal2 s 485464 -960 485688 480 0 FreeSans 896 90 0 0 la_oenb[47]
port 283 nsew signal input
flabel metal2 s 491176 -960 491400 480 0 FreeSans 896 90 0 0 la_oenb[48]
port 284 nsew signal input
flabel metal2 s 496888 -960 497112 480 0 FreeSans 896 90 0 0 la_oenb[49]
port 285 nsew signal input
flabel metal2 s 239848 -960 240072 480 0 FreeSans 896 90 0 0 la_oenb[4]
port 286 nsew signal input
flabel metal2 s 502600 -960 502824 480 0 FreeSans 896 90 0 0 la_oenb[50]
port 287 nsew signal input
flabel metal2 s 508312 -960 508536 480 0 FreeSans 896 90 0 0 la_oenb[51]
port 288 nsew signal input
flabel metal2 s 514024 -960 514248 480 0 FreeSans 896 90 0 0 la_oenb[52]
port 289 nsew signal input
flabel metal2 s 519736 -960 519960 480 0 FreeSans 896 90 0 0 la_oenb[53]
port 290 nsew signal input
flabel metal2 s 525448 -960 525672 480 0 FreeSans 896 90 0 0 la_oenb[54]
port 291 nsew signal input
flabel metal2 s 531160 -960 531384 480 0 FreeSans 896 90 0 0 la_oenb[55]
port 292 nsew signal input
flabel metal2 s 536872 -960 537096 480 0 FreeSans 896 90 0 0 la_oenb[56]
port 293 nsew signal input
flabel metal2 s 542584 -960 542808 480 0 FreeSans 896 90 0 0 la_oenb[57]
port 294 nsew signal input
flabel metal2 s 548296 -960 548520 480 0 FreeSans 896 90 0 0 la_oenb[58]
port 295 nsew signal input
flabel metal2 s 554008 -960 554232 480 0 FreeSans 896 90 0 0 la_oenb[59]
port 296 nsew signal input
flabel metal2 s 245560 -960 245784 480 0 FreeSans 896 90 0 0 la_oenb[5]
port 297 nsew signal input
flabel metal2 s 559720 -960 559944 480 0 FreeSans 896 90 0 0 la_oenb[60]
port 298 nsew signal input
flabel metal2 s 565432 -960 565656 480 0 FreeSans 896 90 0 0 la_oenb[61]
port 299 nsew signal input
flabel metal2 s 571144 -960 571368 480 0 FreeSans 896 90 0 0 la_oenb[62]
port 300 nsew signal input
flabel metal2 s 576856 -960 577080 480 0 FreeSans 896 90 0 0 la_oenb[63]
port 301 nsew signal input
flabel metal2 s 251272 -960 251496 480 0 FreeSans 896 90 0 0 la_oenb[6]
port 302 nsew signal input
flabel metal2 s 256984 -960 257208 480 0 FreeSans 896 90 0 0 la_oenb[7]
port 303 nsew signal input
flabel metal2 s 262696 -960 262920 480 0 FreeSans 896 90 0 0 la_oenb[8]
port 304 nsew signal input
flabel metal2 s 268408 -960 268632 480 0 FreeSans 896 90 0 0 la_oenb[9]
port 305 nsew signal input
flabel metal2 s 578760 -960 578984 480 0 FreeSans 896 90 0 0 user_clock2
port 306 nsew signal input
flabel metal2 s 580664 -960 580888 480 0 FreeSans 896 90 0 0 user_irq[0]
port 307 nsew signal tristate
flabel metal2 s 582568 -960 582792 480 0 FreeSans 896 90 0 0 user_irq[1]
port 308 nsew signal tristate
flabel metal2 s 584472 -960 584696 480 0 FreeSans 896 90 0 0 user_irq[2]
port 309 nsew signal tristate
flabel metal4 s -956 -684 -336 597308 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -956 -684 597020 -64 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -956 596688 597020 597308 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 596400 -684 597020 597308 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 3154 -1644 3774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 21154 -1644 21774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 39154 -1644 39774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 57154 -1644 57774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 75154 -1644 75774 31350 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 75154 219134 75774 242964 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 93154 -1644 93774 31350 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 93154 219134 93774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 111154 -1644 111774 31350 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 111154 219134 111774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 129154 -1644 129774 31350 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 129154 219134 129774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 147154 -1644 147774 31350 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 147154 219134 147774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 165154 -1644 165774 31350 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 165154 219134 165774 242964 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 183154 -1644 183774 31350 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 183154 219134 183774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 201154 -1644 201774 31350 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 201154 219134 201774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 219154 -1644 219774 31350 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 219154 219134 219774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 237154 -1644 237774 31350 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 237154 219134 237774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 255154 -1644 255774 242964 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 273154 -1644 273774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 291154 -1644 291774 79330 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 291154 158782 291774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 309154 -1644 309774 79330 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 309154 158782 309774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 327154 -1644 327774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 345154 -1644 345774 242964 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 363154 -1644 363774 41266 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 363154 217934 363774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 381154 -1644 381774 41266 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 381154 217934 381774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 399154 -1644 399774 41266 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 399154 217934 399774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 417154 -1644 417774 41266 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 417154 217934 417774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 435154 -1644 435774 40964 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 435154 218572 435774 242964 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 453154 -1644 453774 41266 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 453154 217934 453774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 471154 -1644 471774 41266 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 471154 217934 471774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 489154 -1644 489774 41266 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 489154 217934 489774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 507154 -1644 507774 41266 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 507154 217934 507774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 525154 -1644 525774 40964 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 525154 218572 525774 242964 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 543154 -1644 543774 41266 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 543154 217934 543774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 561154 -1644 561774 11154 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 561154 20830 561774 380034 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 561154 487822 561774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 579154 -1644 579774 10964 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 579154 58428 579774 380034 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 579154 487822 579774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 3826 597980 4446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 21826 597980 22446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 39826 66564 40446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 57826 66564 58446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 75826 66564 76446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 93826 66564 94446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 111826 66564 112446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 129826 66564 130446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 147826 66564 148446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 165826 66564 166446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 183826 66564 184446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 201826 597980 202446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 219826 597980 220446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 237826 597980 238446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 255826 597980 256446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 273826 597980 274446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 291826 597980 292446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 309826 597980 310446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 327826 597980 328446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 345826 597980 346446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 363826 597980 364446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 381826 597980 382446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 399826 597980 400446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 417826 597980 418446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 435826 597980 436446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 453826 597980 454446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 471826 597980 472446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 489826 597980 490446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 507826 597980 508446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 525826 597980 526446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 543826 597980 544446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 561826 597980 562446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 579826 597980 580446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s 239468 39826 597980 40446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s 239468 57826 350740 58446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s 239468 75826 350740 76446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s 239468 93826 350740 94446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s 239468 111826 350740 112446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s 239468 129826 350740 130446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s 239468 147826 350740 148446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s 239468 165826 350740 166446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s 239468 183826 350740 184446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s 545484 57826 597980 58446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s 545484 75826 597980 76446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s 545484 93826 597980 94446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s 545484 111826 597980 112446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s 545484 129826 597980 130446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s 545484 147826 597980 148446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s 545484 165826 597980 166446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s 545484 183826 597980 184446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s -1916 -1644 -1296 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 -1644 597980 -1024 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 597648 597980 598268 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 597360 -1644 597980 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 6874 -1644 7494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 24874 -1644 25494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 42874 -1644 43494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 60874 -1644 61494 31350 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 60874 219134 61494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 78874 -1644 79494 31350 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 78874 219134 79494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 96874 -1644 97494 31350 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 96874 219134 97494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 114874 -1644 115494 31350 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 114874 219134 115494 242964 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 132874 -1644 133494 31350 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 132874 219134 133494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 150874 -1644 151494 31350 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 150874 219134 151494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 168874 -1644 169494 31350 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 168874 219134 169494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 186874 -1644 187494 30964 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 186874 228956 187494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 204874 -1644 205494 31350 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 204874 219134 205494 242964 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 222874 -1644 223494 31350 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 222874 219134 223494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 240874 -1644 241494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 258874 -1644 259494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 276874 -1644 277494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 294874 -1644 295494 70964 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 294874 168604 295494 242964 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 312874 -1644 313494 79330 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 312874 158782 313494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 330874 -1644 331494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 348874 -1644 349494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 366874 -1644 367494 41266 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 366874 217934 367494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 384874 -1644 385494 40964 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 402874 -1644 403494 41266 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 402874 217934 403494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 420874 -1644 421494 41266 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 420874 217934 421494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 438874 -1644 439494 41266 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 438874 217934 439494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 456874 -1644 457494 41266 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 456874 217934 457494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 474874 -1644 475494 40964 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 492874 -1644 493494 41266 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 492874 217934 493494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 510874 -1644 511494 41266 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 510874 217934 511494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 528874 -1644 529494 41266 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 528874 217934 529494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 546874 -1644 547494 41266 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 546874 217934 547494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 564874 -1644 565494 11154 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 564874 20830 565494 379396 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 564874 500556 565494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 582874 -1644 583494 380034 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 582874 487822 583494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 9826 597980 10446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 27826 597980 28446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 45826 66564 46446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 63826 66564 64446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 81826 66564 82446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 99826 66564 100446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 117826 66564 118446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 135826 66564 136446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 153826 66564 154446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 171826 66564 172446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 189826 66564 190446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 207826 597980 208446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 225826 597980 226446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 243826 597980 244446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 261826 597980 262446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 279826 597980 280446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 297826 597980 298446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 315826 597980 316446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 333826 597980 334446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 351826 597980 352446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 369826 597980 370446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 387826 597980 388446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 405826 597980 406446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 423826 597980 424446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 441826 597980 442446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 459826 597980 460446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 477826 597980 478446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 495826 597980 496446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 513826 597980 514446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 531826 597980 532446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 549826 597980 550446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 567826 597980 568446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 585826 597980 586446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s 239468 45826 350740 46446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s 239468 63826 350740 64446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s 239468 81826 350740 82446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s 239468 99826 350740 100446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s 239468 117826 350740 118446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s 239468 135826 350740 136446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s 239468 153826 350740 154446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s 239468 171826 350740 172446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s 239468 189826 350740 190446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s 545484 45826 597980 46446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s 545484 63826 597980 64446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s 545484 81826 597980 82446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s 545484 99826 597980 100446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s 545484 117826 597980 118446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s 545484 135826 597980 136446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s 545484 153826 597980 154446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s 545484 171826 597980 172446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s 545484 189826 597980 190446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal2 s 11368 -960 11592 480 0 FreeSans 896 90 0 0 wb_clk_i
port 312 nsew signal input
flabel metal2 s 13272 -960 13496 480 0 FreeSans 896 90 0 0 wb_rst_i
port 313 nsew signal input
flabel metal2 s 15176 -960 15400 480 0 FreeSans 896 90 0 0 wbs_ack_o
port 314 nsew signal tristate
flabel metal2 s 22792 -960 23016 480 0 FreeSans 896 90 0 0 wbs_adr_i[0]
port 315 nsew signal input
flabel metal2 s 87528 -960 87752 480 0 FreeSans 896 90 0 0 wbs_adr_i[10]
port 316 nsew signal input
flabel metal2 s 93240 -960 93464 480 0 FreeSans 896 90 0 0 wbs_adr_i[11]
port 317 nsew signal input
flabel metal2 s 98952 -960 99176 480 0 FreeSans 896 90 0 0 wbs_adr_i[12]
port 318 nsew signal input
flabel metal2 s 104664 -960 104888 480 0 FreeSans 896 90 0 0 wbs_adr_i[13]
port 319 nsew signal input
flabel metal2 s 110376 -960 110600 480 0 FreeSans 896 90 0 0 wbs_adr_i[14]
port 320 nsew signal input
flabel metal2 s 116088 -960 116312 480 0 FreeSans 896 90 0 0 wbs_adr_i[15]
port 321 nsew signal input
flabel metal2 s 121800 -960 122024 480 0 FreeSans 896 90 0 0 wbs_adr_i[16]
port 322 nsew signal input
flabel metal2 s 127512 -960 127736 480 0 FreeSans 896 90 0 0 wbs_adr_i[17]
port 323 nsew signal input
flabel metal2 s 133224 -960 133448 480 0 FreeSans 896 90 0 0 wbs_adr_i[18]
port 324 nsew signal input
flabel metal2 s 138936 -960 139160 480 0 FreeSans 896 90 0 0 wbs_adr_i[19]
port 325 nsew signal input
flabel metal2 s 30408 -960 30632 480 0 FreeSans 896 90 0 0 wbs_adr_i[1]
port 326 nsew signal input
flabel metal2 s 144648 -960 144872 480 0 FreeSans 896 90 0 0 wbs_adr_i[20]
port 327 nsew signal input
flabel metal2 s 150360 -960 150584 480 0 FreeSans 896 90 0 0 wbs_adr_i[21]
port 328 nsew signal input
flabel metal2 s 156072 -960 156296 480 0 FreeSans 896 90 0 0 wbs_adr_i[22]
port 329 nsew signal input
flabel metal2 s 161784 -960 162008 480 0 FreeSans 896 90 0 0 wbs_adr_i[23]
port 330 nsew signal input
flabel metal2 s 167496 -960 167720 480 0 FreeSans 896 90 0 0 wbs_adr_i[24]
port 331 nsew signal input
flabel metal2 s 173208 -960 173432 480 0 FreeSans 896 90 0 0 wbs_adr_i[25]
port 332 nsew signal input
flabel metal2 s 178920 -960 179144 480 0 FreeSans 896 90 0 0 wbs_adr_i[26]
port 333 nsew signal input
flabel metal2 s 184632 -960 184856 480 0 FreeSans 896 90 0 0 wbs_adr_i[27]
port 334 nsew signal input
flabel metal2 s 190344 -960 190568 480 0 FreeSans 896 90 0 0 wbs_adr_i[28]
port 335 nsew signal input
flabel metal2 s 196056 -960 196280 480 0 FreeSans 896 90 0 0 wbs_adr_i[29]
port 336 nsew signal input
flabel metal2 s 38024 -960 38248 480 0 FreeSans 896 90 0 0 wbs_adr_i[2]
port 337 nsew signal input
flabel metal2 s 201768 -960 201992 480 0 FreeSans 896 90 0 0 wbs_adr_i[30]
port 338 nsew signal input
flabel metal2 s 207480 -960 207704 480 0 FreeSans 896 90 0 0 wbs_adr_i[31]
port 339 nsew signal input
flabel metal2 s 45640 -960 45864 480 0 FreeSans 896 90 0 0 wbs_adr_i[3]
port 340 nsew signal input
flabel metal2 s 53256 -960 53480 480 0 FreeSans 896 90 0 0 wbs_adr_i[4]
port 341 nsew signal input
flabel metal2 s 58968 -960 59192 480 0 FreeSans 896 90 0 0 wbs_adr_i[5]
port 342 nsew signal input
flabel metal2 s 64680 -960 64904 480 0 FreeSans 896 90 0 0 wbs_adr_i[6]
port 343 nsew signal input
flabel metal2 s 70392 -960 70616 480 0 FreeSans 896 90 0 0 wbs_adr_i[7]
port 344 nsew signal input
flabel metal2 s 76104 -960 76328 480 0 FreeSans 896 90 0 0 wbs_adr_i[8]
port 345 nsew signal input
flabel metal2 s 81816 -960 82040 480 0 FreeSans 896 90 0 0 wbs_adr_i[9]
port 346 nsew signal input
flabel metal2 s 17080 -960 17304 480 0 FreeSans 896 90 0 0 wbs_cyc_i
port 347 nsew signal input
flabel metal2 s 24696 -960 24920 480 0 FreeSans 896 90 0 0 wbs_dat_i[0]
port 348 nsew signal input
flabel metal2 s 89432 -960 89656 480 0 FreeSans 896 90 0 0 wbs_dat_i[10]
port 349 nsew signal input
flabel metal2 s 95144 -960 95368 480 0 FreeSans 896 90 0 0 wbs_dat_i[11]
port 350 nsew signal input
flabel metal2 s 100856 -960 101080 480 0 FreeSans 896 90 0 0 wbs_dat_i[12]
port 351 nsew signal input
flabel metal2 s 106568 -960 106792 480 0 FreeSans 896 90 0 0 wbs_dat_i[13]
port 352 nsew signal input
flabel metal2 s 112280 -960 112504 480 0 FreeSans 896 90 0 0 wbs_dat_i[14]
port 353 nsew signal input
flabel metal2 s 117992 -960 118216 480 0 FreeSans 896 90 0 0 wbs_dat_i[15]
port 354 nsew signal input
flabel metal2 s 123704 -960 123928 480 0 FreeSans 896 90 0 0 wbs_dat_i[16]
port 355 nsew signal input
flabel metal2 s 129416 -960 129640 480 0 FreeSans 896 90 0 0 wbs_dat_i[17]
port 356 nsew signal input
flabel metal2 s 135128 -960 135352 480 0 FreeSans 896 90 0 0 wbs_dat_i[18]
port 357 nsew signal input
flabel metal2 s 140840 -960 141064 480 0 FreeSans 896 90 0 0 wbs_dat_i[19]
port 358 nsew signal input
flabel metal2 s 32312 -960 32536 480 0 FreeSans 896 90 0 0 wbs_dat_i[1]
port 359 nsew signal input
flabel metal2 s 146552 -960 146776 480 0 FreeSans 896 90 0 0 wbs_dat_i[20]
port 360 nsew signal input
flabel metal2 s 152264 -960 152488 480 0 FreeSans 896 90 0 0 wbs_dat_i[21]
port 361 nsew signal input
flabel metal2 s 157976 -960 158200 480 0 FreeSans 896 90 0 0 wbs_dat_i[22]
port 362 nsew signal input
flabel metal2 s 163688 -960 163912 480 0 FreeSans 896 90 0 0 wbs_dat_i[23]
port 363 nsew signal input
flabel metal2 s 169400 -960 169624 480 0 FreeSans 896 90 0 0 wbs_dat_i[24]
port 364 nsew signal input
flabel metal2 s 175112 -960 175336 480 0 FreeSans 896 90 0 0 wbs_dat_i[25]
port 365 nsew signal input
flabel metal2 s 180824 -960 181048 480 0 FreeSans 896 90 0 0 wbs_dat_i[26]
port 366 nsew signal input
flabel metal2 s 186536 -960 186760 480 0 FreeSans 896 90 0 0 wbs_dat_i[27]
port 367 nsew signal input
flabel metal2 s 192248 -960 192472 480 0 FreeSans 896 90 0 0 wbs_dat_i[28]
port 368 nsew signal input
flabel metal2 s 197960 -960 198184 480 0 FreeSans 896 90 0 0 wbs_dat_i[29]
port 369 nsew signal input
flabel metal2 s 39928 -960 40152 480 0 FreeSans 896 90 0 0 wbs_dat_i[2]
port 370 nsew signal input
flabel metal2 s 203672 -960 203896 480 0 FreeSans 896 90 0 0 wbs_dat_i[30]
port 371 nsew signal input
flabel metal2 s 209384 -960 209608 480 0 FreeSans 896 90 0 0 wbs_dat_i[31]
port 372 nsew signal input
flabel metal2 s 47544 -960 47768 480 0 FreeSans 896 90 0 0 wbs_dat_i[3]
port 373 nsew signal input
flabel metal2 s 55160 -960 55384 480 0 FreeSans 896 90 0 0 wbs_dat_i[4]
port 374 nsew signal input
flabel metal2 s 60872 -960 61096 480 0 FreeSans 896 90 0 0 wbs_dat_i[5]
port 375 nsew signal input
flabel metal2 s 66584 -960 66808 480 0 FreeSans 896 90 0 0 wbs_dat_i[6]
port 376 nsew signal input
flabel metal2 s 72296 -960 72520 480 0 FreeSans 896 90 0 0 wbs_dat_i[7]
port 377 nsew signal input
flabel metal2 s 78008 -960 78232 480 0 FreeSans 896 90 0 0 wbs_dat_i[8]
port 378 nsew signal input
flabel metal2 s 83720 -960 83944 480 0 FreeSans 896 90 0 0 wbs_dat_i[9]
port 379 nsew signal input
flabel metal2 s 26600 -960 26824 480 0 FreeSans 896 90 0 0 wbs_dat_o[0]
port 380 nsew signal tristate
flabel metal2 s 91336 -960 91560 480 0 FreeSans 896 90 0 0 wbs_dat_o[10]
port 381 nsew signal tristate
flabel metal2 s 97048 -960 97272 480 0 FreeSans 896 90 0 0 wbs_dat_o[11]
port 382 nsew signal tristate
flabel metal2 s 102760 -960 102984 480 0 FreeSans 896 90 0 0 wbs_dat_o[12]
port 383 nsew signal tristate
flabel metal2 s 108472 -960 108696 480 0 FreeSans 896 90 0 0 wbs_dat_o[13]
port 384 nsew signal tristate
flabel metal2 s 114184 -960 114408 480 0 FreeSans 896 90 0 0 wbs_dat_o[14]
port 385 nsew signal tristate
flabel metal2 s 119896 -960 120120 480 0 FreeSans 896 90 0 0 wbs_dat_o[15]
port 386 nsew signal tristate
flabel metal2 s 125608 -960 125832 480 0 FreeSans 896 90 0 0 wbs_dat_o[16]
port 387 nsew signal tristate
flabel metal2 s 131320 -960 131544 480 0 FreeSans 896 90 0 0 wbs_dat_o[17]
port 388 nsew signal tristate
flabel metal2 s 137032 -960 137256 480 0 FreeSans 896 90 0 0 wbs_dat_o[18]
port 389 nsew signal tristate
flabel metal2 s 142744 -960 142968 480 0 FreeSans 896 90 0 0 wbs_dat_o[19]
port 390 nsew signal tristate
flabel metal2 s 34216 -960 34440 480 0 FreeSans 896 90 0 0 wbs_dat_o[1]
port 391 nsew signal tristate
flabel metal2 s 148456 -960 148680 480 0 FreeSans 896 90 0 0 wbs_dat_o[20]
port 392 nsew signal tristate
flabel metal2 s 154168 -960 154392 480 0 FreeSans 896 90 0 0 wbs_dat_o[21]
port 393 nsew signal tristate
flabel metal2 s 159880 -960 160104 480 0 FreeSans 896 90 0 0 wbs_dat_o[22]
port 394 nsew signal tristate
flabel metal2 s 165592 -960 165816 480 0 FreeSans 896 90 0 0 wbs_dat_o[23]
port 395 nsew signal tristate
flabel metal2 s 171304 -960 171528 480 0 FreeSans 896 90 0 0 wbs_dat_o[24]
port 396 nsew signal tristate
flabel metal2 s 177016 -960 177240 480 0 FreeSans 896 90 0 0 wbs_dat_o[25]
port 397 nsew signal tristate
flabel metal2 s 182728 -960 182952 480 0 FreeSans 896 90 0 0 wbs_dat_o[26]
port 398 nsew signal tristate
flabel metal2 s 188440 -960 188664 480 0 FreeSans 896 90 0 0 wbs_dat_o[27]
port 399 nsew signal tristate
flabel metal2 s 194152 -960 194376 480 0 FreeSans 896 90 0 0 wbs_dat_o[28]
port 400 nsew signal tristate
flabel metal2 s 199864 -960 200088 480 0 FreeSans 896 90 0 0 wbs_dat_o[29]
port 401 nsew signal tristate
flabel metal2 s 41832 -960 42056 480 0 FreeSans 896 90 0 0 wbs_dat_o[2]
port 402 nsew signal tristate
flabel metal2 s 205576 -960 205800 480 0 FreeSans 896 90 0 0 wbs_dat_o[30]
port 403 nsew signal tristate
flabel metal2 s 211288 -960 211512 480 0 FreeSans 896 90 0 0 wbs_dat_o[31]
port 404 nsew signal tristate
flabel metal2 s 49448 -960 49672 480 0 FreeSans 896 90 0 0 wbs_dat_o[3]
port 405 nsew signal tristate
flabel metal2 s 57064 -960 57288 480 0 FreeSans 896 90 0 0 wbs_dat_o[4]
port 406 nsew signal tristate
flabel metal2 s 62776 -960 63000 480 0 FreeSans 896 90 0 0 wbs_dat_o[5]
port 407 nsew signal tristate
flabel metal2 s 68488 -960 68712 480 0 FreeSans 896 90 0 0 wbs_dat_o[6]
port 408 nsew signal tristate
flabel metal2 s 74200 -960 74424 480 0 FreeSans 896 90 0 0 wbs_dat_o[7]
port 409 nsew signal tristate
flabel metal2 s 79912 -960 80136 480 0 FreeSans 896 90 0 0 wbs_dat_o[8]
port 410 nsew signal tristate
flabel metal2 s 85624 -960 85848 480 0 FreeSans 896 90 0 0 wbs_dat_o[9]
port 411 nsew signal tristate
flabel metal2 s 28504 -960 28728 480 0 FreeSans 896 90 0 0 wbs_sel_i[0]
port 412 nsew signal input
flabel metal2 s 36120 -960 36344 480 0 FreeSans 896 90 0 0 wbs_sel_i[1]
port 413 nsew signal input
flabel metal2 s 43736 -960 43960 480 0 FreeSans 896 90 0 0 wbs_sel_i[2]
port 414 nsew signal input
flabel metal2 s 51352 -960 51576 480 0 FreeSans 896 90 0 0 wbs_sel_i[3]
port 415 nsew signal input
flabel metal2 s 18984 -960 19208 480 0 FreeSans 896 90 0 0 wbs_stb_i
port 416 nsew signal input
flabel metal2 s 20888 -960 21112 480 0 FreeSans 896 90 0 0 wbs_we_i
port 417 nsew signal input
rlabel via4 579166 40384 579166 40384 0 vdd
rlabel via4 589166 46384 589166 46384 0 vss
rlabel metal2 85400 230174 85400 230174 0 i2c_rst_n
rlabel metal2 456792 226632 456792 226632 0 i2cm_clk_i
rlabel metal2 474824 225078 474824 225078 0 i2cm_clk_o
rlabel metal2 491400 224742 491400 224742 0 i2cm_clk_oen
rlabel metal2 185752 230118 185752 230118 0 i2cm_data_i
rlabel metal2 524104 226632 524104 226632 0 i2cm_data_o
rlabel metal2 171416 230230 171416 230230 0 i2cm_data_oen
rlabel metal3 551334 134792 551334 134792 0 i2cm_intr_o
rlabel metal2 187544 592522 187544 592522 0 io_in[21]
rlabel metal2 121352 592578 121352 592578 0 io_in[22]
rlabel metal2 55160 593194 55160 593194 0 io_in[23]
rlabel metal3 19110 587160 19110 587160 0 io_in[24]
rlabel metal3 3150 544824 3150 544824 0 io_in[25]
rlabel metal3 36330 168056 36330 168056 0 io_in[26]
rlabel metal3 7350 460152 7350 460152 0 io_in[27]
rlabel metal3 38010 145208 38010 145208 0 io_in[28]
rlabel metal3 9030 375480 9030 375480 0 io_in[29]
rlabel metal3 9926 333144 9926 333144 0 io_in[30]
rlabel metal4 22792 202104 22792 202104 0 io_in[31]
rlabel metal4 27832 175056 27832 175056 0 io_in[32]
rlabel metal4 29512 147112 29512 147112 0 io_in[33]
rlabel metal3 6510 163800 6510 163800 0 io_in[34]
rlabel metal3 7350 121464 7350 121464 0 io_in[35]
rlabel metal3 2422 79128 2422 79128 0 io_in[36]
rlabel metal3 2310 36904 2310 36904 0 io_in[37]
rlabel metal3 592256 60424 592256 60424 0 io_in[5]
rlabel metal3 592368 60312 592368 60312 0 io_in[6]
rlabel metal3 593082 430136 593082 430136 0 io_oeb[10]
rlabel metal3 584794 548968 584794 548968 0 io_oeb[13]
rlabel metal2 572152 544278 572152 544278 0 io_oeb[14]
rlabel metal4 540792 589512 540792 589512 0 io_oeb[15]
rlabel metal4 474600 589512 474600 589512 0 io_oeb[16]
rlabel metal2 566776 544390 566776 544390 0 io_oeb[17]
rlabel metal3 564312 503944 564312 503944 0 io_oeb[18]
rlabel metal2 563192 501326 563192 501326 0 io_oeb[19]
rlabel metal2 209832 592522 209832 592522 0 io_oeb[20]
rlabel metal2 143416 593138 143416 593138 0 io_oeb[21]
rlabel metal4 77336 589288 77336 589288 0 io_oeb[22]
rlabel metal2 53816 203224 53816 203224 0 io_oeb[23]
rlabel metal3 18270 558936 18270 558936 0 io_oeb[24]
rlabel metal3 17430 516600 17430 516600 0 io_oeb[25]
rlabel metal3 3206 474264 3206 474264 0 io_oeb[26]
rlabel metal4 31080 291144 31080 291144 0 io_oeb[27]
rlabel metal3 4830 389592 4830 389592 0 io_oeb[28]
rlabel metal4 29400 236712 29400 236712 0 io_oeb[29]
rlabel metal3 16590 304920 16590 304920 0 io_oeb[30]
rlabel metal3 3262 262584 3262 262584 0 io_oeb[31]
rlabel metal3 2422 220248 2422 220248 0 io_oeb[32]
rlabel metal3 4886 177912 4886 177912 0 io_oeb[33]
rlabel metal3 2310 135576 2310 135576 0 io_oeb[34]
rlabel metal3 3150 93240 3150 93240 0 io_oeb[35]
rlabel metal4 5096 49392 5096 49392 0 io_oeb[36]
rlabel metal3 2310 8792 2310 8792 0 io_oeb[37]
rlabel metal3 594314 231896 594314 231896 0 io_oeb[5]
rlabel metal5 592312 30150 592312 30150 0 io_oeb[6]
rlabel metal3 586026 311080 586026 311080 0 io_oeb[7]
rlabel metal3 591402 350728 591402 350728 0 io_oeb[8]
rlabel metal3 593194 390376 593194 390376 0 io_oeb[9]
rlabel metal3 589736 379736 589736 379736 0 io_out[10]
rlabel metal3 591962 535752 591962 535752 0 io_out[13]
rlabel metal3 591066 575400 591066 575400 0 io_out[14]
rlabel metal2 562744 593082 562744 593082 0 io_out[15]
rlabel metal2 496664 593306 496664 593306 0 io_out[16]
rlabel metal2 430472 593250 430472 593250 0 io_out[17]
rlabel metal2 364280 593194 364280 593194 0 io_out[18]
rlabel metal2 298088 593138 298088 593138 0 io_out[19]
rlabel metal2 231784 593082 231784 593082 0 io_out[20]
rlabel metal2 165480 593082 165480 593082 0 io_out[21]
rlabel metal2 99288 592634 99288 592634 0 io_out[22]
rlabel metal2 33096 397082 33096 397082 0 io_out[23]
rlabel metal4 27720 380072 27720 380072 0 io_out[24]
rlabel metal4 22680 353192 22680 353192 0 io_out[25]
rlabel metal3 2310 488376 2310 488376 0 io_out[26]
rlabel metal3 9870 446040 9870 446040 0 io_out[27]
rlabel metal3 2366 403704 2366 403704 0 io_out[28]
rlabel metal3 19166 361368 19166 361368 0 io_out[29]
rlabel metal4 57064 119336 57064 119336 0 io_out[30]
rlabel metal3 17486 276696 17486 276696 0 io_out[31]
rlabel metal4 44520 165480 44520 165480 0 io_out[32]
rlabel metal3 20790 192024 20790 192024 0 io_out[33]
rlabel metal3 35490 72856 35490 72856 0 io_out[34]
rlabel metal3 2366 107352 2366 107352 0 io_out[35]
rlabel metal3 2310 65016 2310 65016 0 io_out[36]
rlabel metal3 2366 22904 2366 22904 0 io_out[37]
rlabel metal3 592298 297864 592298 297864 0 io_out[7]
rlabel metal3 593418 337512 593418 337512 0 io_out[8]
rlabel metal2 590184 376320 590184 376320 0 io_out[9]
rlabel metal3 241542 220696 241542 220696 0 reg_peri_ack
rlabel metal3 241094 81592 241094 81592 0 reg_peri_addr\[0\]
rlabel metal4 275576 74928 275576 74928 0 reg_peri_addr\[10\]
rlabel metal3 241150 79576 241150 79576 0 reg_peri_addr\[1\]
rlabel metal3 241374 77560 241374 77560 0 reg_peri_addr\[2\]
rlabel metal3 242270 75544 242270 75544 0 reg_peri_addr\[3\]
rlabel metal3 257390 73528 257390 73528 0 reg_peri_addr\[4\]
rlabel metal3 241598 71512 241598 71512 0 reg_peri_addr\[5\]
rlabel metal3 241654 69496 241654 69496 0 reg_peri_addr\[6\]
rlabel metal3 241542 67480 241542 67480 0 reg_peri_addr\[7\]
rlabel metal3 241430 65464 241430 65464 0 reg_peri_addr\[8\]
rlabel metal3 241486 63448 241486 63448 0 reg_peri_addr\[9\]
rlabel metal3 241598 89656 241598 89656 0 reg_peri_be\[0\]
rlabel metal3 241542 87640 241542 87640 0 reg_peri_be\[1\]
rlabel metal3 241038 85624 241038 85624 0 reg_peri_be\[2\]
rlabel metal3 240982 83608 240982 83608 0 reg_peri_be\[3\]
rlabel metal3 241374 57400 241374 57400 0 reg_peri_cs
rlabel metal3 243054 218680 243054 218680 0 reg_peri_rdata\[0\]
rlabel metal3 275674 152936 275674 152936 0 reg_peri_rdata\[10\]
rlabel metal4 261240 174160 261240 174160 0 reg_peri_rdata\[11\]
rlabel metal3 254814 194488 254814 194488 0 reg_peri_rdata\[12\]
rlabel metal4 262920 171024 262920 171024 0 reg_peri_rdata\[13\]
rlabel metal4 257880 169456 257880 169456 0 reg_peri_rdata\[14\]
rlabel metal3 243894 188440 243894 188440 0 reg_peri_rdata\[15\]
rlabel metal3 273994 146216 273994 146216 0 reg_peri_rdata\[16\]
rlabel metal3 264754 145096 264754 145096 0 reg_peri_rdata\[17\]
rlabel metal4 264712 163184 264712 163184 0 reg_peri_rdata\[18\]
rlabel metal3 265650 142856 265650 142856 0 reg_peri_rdata\[19\]
rlabel metal4 266280 189840 266280 189840 0 reg_peri_rdata\[1\]
rlabel metal3 266490 141736 266490 141736 0 reg_peri_rdata\[20\]
rlabel metal3 277410 140616 277410 140616 0 reg_peri_rdata\[21\]
rlabel metal3 263130 139496 263130 139496 0 reg_peri_rdata\[22\]
rlabel metal3 240982 172312 240982 172312 0 reg_peri_rdata\[23\]
rlabel metal3 255710 170296 255710 170296 0 reg_peri_rdata\[24\]
rlabel metal4 261352 153440 261352 153440 0 reg_peri_rdata\[25\]
rlabel metal3 243950 166264 243950 166264 0 reg_peri_rdata\[26\]
rlabel metal4 263032 149072 263032 149072 0 reg_peri_rdata\[27\]
rlabel metal3 242270 162232 242270 162232 0 reg_peri_rdata\[28\]
rlabel metal3 274890 131656 274890 131656 0 reg_peri_rdata\[29\]
rlabel metal3 246414 214648 246414 214648 0 reg_peri_rdata\[2\]
rlabel metal4 257992 145040 257992 145040 0 reg_peri_rdata\[30\]
rlabel metal3 277354 129416 277354 129416 0 reg_peri_rdata\[31\]
rlabel metal3 241486 212632 241486 212632 0 reg_peri_rdata\[3\]
rlabel metal3 245574 210616 245574 210616 0 reg_peri_rdata\[4\]
rlabel metal3 241374 208600 241374 208600 0 reg_peri_rdata\[5\]
rlabel metal3 241542 206584 241542 206584 0 reg_peri_rdata\[6\]
rlabel metal3 241430 204568 241430 204568 0 reg_peri_rdata\[7\]
rlabel metal3 241598 202552 241598 202552 0 reg_peri_rdata\[8\]
rlabel metal4 264600 177968 264600 177968 0 reg_peri_rdata\[9\]
rlabel metal3 240982 154168 240982 154168 0 reg_peri_wdata\[0\]
rlabel metal3 266434 117096 266434 117096 0 reg_peri_wdata\[10\]
rlabel metal4 258216 123984 258216 123984 0 reg_peri_wdata\[11\]
rlabel metal3 262290 114856 262290 114856 0 reg_peri_wdata\[12\]
rlabel metal3 274162 113736 274162 113736 0 reg_peri_wdata\[13\]
rlabel metal3 241654 125944 241654 125944 0 reg_peri_wdata\[14\]
rlabel metal3 243054 123928 243054 123928 0 reg_peri_wdata\[15\]
rlabel metal3 241374 121912 241374 121912 0 reg_peri_wdata\[16\]
rlabel metal3 241486 119896 241486 119896 0 reg_peri_wdata\[17\]
rlabel metal3 241542 117880 241542 117880 0 reg_peri_wdata\[18\]
rlabel metal3 241766 115864 241766 115864 0 reg_peri_wdata\[19\]
rlabel metal4 264600 139664 264600 139664 0 reg_peri_wdata\[1\]
rlabel metal3 241094 113848 241094 113848 0 reg_peri_wdata\[20\]
rlabel metal3 241038 111832 241038 111832 0 reg_peri_wdata\[21\]
rlabel metal3 241150 109816 241150 109816 0 reg_peri_wdata\[22\]
rlabel metal3 240982 107800 240982 107800 0 reg_peri_wdata\[23\]
rlabel metal3 241542 105784 241542 105784 0 reg_peri_wdata\[24\]
rlabel metal4 275576 100968 275576 100968 0 reg_peri_wdata\[25\]
rlabel metal4 273896 100464 273896 100464 0 reg_peri_wdata\[26\]
rlabel metal3 240982 99736 240982 99736 0 reg_peri_wdata\[27\]
rlabel metal3 239960 97594 239960 97594 0 reg_peri_wdata\[28\]
rlabel metal3 241794 95704 241794 95704 0 reg_peri_wdata\[29\]
rlabel metal3 241542 150136 241542 150136 0 reg_peri_wdata\[2\]
rlabel metal3 239960 93870 239960 93870 0 reg_peri_wdata\[30\]
rlabel metal3 240982 91672 240982 91672 0 reg_peri_wdata\[31\]
rlabel metal3 241374 148120 241374 148120 0 reg_peri_wdata\[3\]
rlabel metal3 241430 146104 241430 146104 0 reg_peri_wdata\[4\]
rlabel metal3 241542 144088 241542 144088 0 reg_peri_wdata\[5\]
rlabel metal3 241486 142072 241486 142072 0 reg_peri_wdata\[6\]
rlabel metal3 241598 140056 241598 140056 0 reg_peri_wdata\[7\]
rlabel metal3 241710 138040 241710 138040 0 reg_peri_wdata\[8\]
rlabel metal4 275576 120008 275576 120008 0 reg_peri_wdata\[9\]
rlabel metal3 277354 75656 277354 75656 0 reg_peri_wr
rlabel metal2 289912 200326 289912 200326 0 rtc_clk
rlabel metal2 309848 171094 309848 171094 0 rtc_intr
rlabel metal2 424984 225512 424984 225512 0 sspim_rst_n
rlabel metal4 193256 228536 193256 228536 0 sspim_sck
rlabel metal3 239344 231896 239344 231896 0 sspim_si
rlabel metal2 240184 228144 240184 228144 0 sspim_so
rlabel metal2 242984 225176 242984 225176 0 sspim_ssn\[0\]
rlabel metal2 214424 231126 214424 231126 0 sspim_ssn\[1\]
rlabel metal3 551334 193928 551334 193928 0 sspim_ssn\[2\]
rlabel metal3 374752 232456 374752 232456 0 sspim_ssn\[3\]
rlabel metal2 78470 229432 78470 229432 0 uart_rst_n\[0\]
rlabel metal2 71064 231070 71064 231070 0 uart_rst_n\[1\]
rlabel metal3 291998 55384 291998 55384 0 uart_rxd\[0\]
rlabel metal4 350168 43288 350168 43288 0 uart_rxd\[1\]
rlabel metal4 350616 44184 350616 44184 0 uart_txd\[0\]
rlabel metal3 241486 49336 241486 49336 0 uart_txd\[1\]
rlabel metal2 106904 230342 106904 230342 0 usb_clk
rlabel metal3 291774 47320 291774 47320 0 usb_dn_i
rlabel metal3 239960 40866 239960 40866 0 usb_dn_o
rlabel metal4 349608 40824 349608 40824 0 usb_dp_i
rlabel metal4 437640 37016 437640 37016 0 usb_dp_o
rlabel metal3 225736 232120 225736 232120 0 usb_intr_o
rlabel metal3 240982 43288 240982 43288 0 usb_oen
rlabel metal2 241976 226184 241976 226184 0 usb_rst_n
rlabel metal3 73360 26936 73360 26936 0 user_clock2
rlabel metal2 562968 6720 562968 6720 0 user_irq[0]
rlabel metal2 582568 2422 582568 2422 0 user_irq[1]
rlabel metal2 584472 2366 584472 2366 0 user_irq[2]
rlabel metal2 69510 30072 69510 30072 0 wb_clk_i
rlabel metal2 78232 25858 78232 25858 0 wb_rst_i
rlabel metal3 350616 216230 350616 216230 0 wbs_ack_o
rlabel metal2 101528 27426 101528 27426 0 wbs_adr_i[0]
rlabel metal2 570318 10136 570318 10136 0 wbs_adr_i[10]
rlabel metal2 93464 1470 93464 1470 0 wbs_adr_i[11]
rlabel metal2 99064 1526 99064 1526 0 wbs_adr_i[12]
rlabel metal2 572600 9842 572600 9842 0 wbs_adr_i[13]
rlabel metal2 110600 1638 110600 1638 0 wbs_adr_i[14]
rlabel metal2 116312 1694 116312 1694 0 wbs_adr_i[15]
rlabel metal2 122024 3150 122024 3150 0 wbs_adr_i[16]
rlabel metal2 127624 3206 127624 3206 0 wbs_adr_i[17]
rlabel metal2 572824 378266 572824 378266 0 wbs_adr_i[18]
rlabel metal2 139272 280 139272 280 0 wbs_adr_i[19]
rlabel metal2 99736 26754 99736 26754 0 wbs_adr_i[1]
rlabel metal2 144984 336 144984 336 0 wbs_adr_i[20]
rlabel metal2 571032 378280 571032 378280 0 wbs_adr_i[21]
rlabel metal3 570640 376600 570640 376600 0 wbs_adr_i[22]
rlabel metal2 162008 462 162008 462 0 wbs_adr_i[23]
rlabel metal2 167720 3374 167720 3374 0 wbs_adr_i[24]
rlabel metal2 569240 7336 569240 7336 0 wbs_adr_i[25]
rlabel metal2 567000 5208 567000 5208 0 wbs_adr_i[26]
rlabel metal2 184856 6384 184856 6384 0 wbs_adr_i[27]
rlabel metal2 190568 4158 190568 4158 0 wbs_adr_i[28]
rlabel metal2 196280 4214 196280 4214 0 wbs_adr_i[29]
rlabel metal2 97944 24850 97944 24850 0 wbs_adr_i[2]
rlabel metal3 568064 376824 568064 376824 0 wbs_adr_i[30]
rlabel metal2 564424 6384 564424 6384 0 wbs_adr_i[31]
rlabel metal2 96152 28266 96152 28266 0 wbs_adr_i[3]
rlabel metal2 94360 27370 94360 27370 0 wbs_adr_i[4]
rlabel metal2 92568 29106 92568 29106 0 wbs_adr_i[5]
rlabel metal2 90776 29218 90776 29218 0 wbs_adr_i[6]
rlabel metal2 70504 3206 70504 3206 0 wbs_adr_i[7]
rlabel metal2 76328 3262 76328 3262 0 wbs_adr_i[8]
rlabel metal2 569016 9898 569016 9898 0 wbs_adr_i[9]
rlabel metal3 586656 376488 586656 376488 0 wbs_cyc_i
rlabel metal2 24920 2366 24920 2366 0 wbs_dat_i[0]
rlabel metal2 147994 30072 147994 30072 0 wbs_dat_i[10]
rlabel metal3 144536 26656 144536 26656 0 wbs_dat_i[11]
rlabel metal2 144536 27482 144536 27482 0 wbs_dat_i[12]
rlabel metal2 106568 8358 106568 8358 0 wbs_dat_i[13]
rlabel metal2 112504 3318 112504 3318 0 wbs_dat_i[14]
rlabel metal2 117992 10094 117992 10094 0 wbs_dat_i[15]
rlabel metal2 123704 6734 123704 6734 0 wbs_dat_i[16]
rlabel metal3 557354 430472 557354 430472 0 wbs_dat_i[17]
rlabel metal2 134848 20160 134848 20160 0 wbs_dat_i[18]
rlabel metal2 131992 29274 131992 29274 0 wbs_dat_i[19]
rlabel metal2 164066 30072 164066 30072 0 wbs_dat_i[1]
rlabel metal2 146216 26264 146216 26264 0 wbs_dat_i[20]
rlabel metal2 128408 25522 128408 25522 0 wbs_dat_i[21]
rlabel via4 451976 39495 451976 39495 0 wbs_dat_i[22]
rlabel metal2 124824 29106 124824 29106 0 wbs_dat_i[23]
rlabel metal2 123032 29050 123032 29050 0 wbs_dat_i[24]
rlabel metal2 121240 28770 121240 28770 0 wbs_dat_i[25]
rlabel metal2 119448 26362 119448 26362 0 wbs_dat_i[26]
rlabel metal2 117656 28826 117656 28826 0 wbs_dat_i[27]
rlabel metal2 115864 28938 115864 28938 0 wbs_dat_i[28]
rlabel metal2 423570 40040 423570 40040 0 wbs_dat_i[29]
rlabel metal2 162456 28714 162456 28714 0 wbs_dat_i[2]
rlabel metal4 238504 31039 238504 31039 0 wbs_dat_i[30]
rlabel metal4 209384 24235 209384 24235 0 wbs_dat_i[31]
rlabel metal2 47544 9030 47544 9030 0 wbs_dat_i[3]
rlabel metal2 55160 10878 55160 10878 0 wbs_dat_i[4]
rlabel metal2 520646 40040 520646 40040 0 wbs_dat_i[5]
rlabel metal2 516488 39858 516488 39858 0 wbs_dat_i[6]
rlabel metal2 72296 13342 72296 13342 0 wbs_dat_i[7]
rlabel metal2 78008 13174 78008 13174 0 wbs_dat_i[8]
rlabel metal3 519904 38696 519904 38696 0 wbs_dat_i[9]
rlabel metal2 26824 2310 26824 2310 0 wbs_dat_o[0]
rlabel metal2 91336 13286 91336 13286 0 wbs_dat_o[10]
rlabel metal2 97048 6510 97048 6510 0 wbs_dat_o[11]
rlabel metal4 209944 30016 209944 30016 0 wbs_dat_o[12]
rlabel metal3 347018 140616 347018 140616 0 wbs_dat_o[13]
rlabel metal2 114408 4942 114408 4942 0 wbs_dat_o[14]
rlabel metal2 119896 9142 119896 9142 0 wbs_dat_o[15]
rlabel metal2 193256 23912 193256 23912 0 wbs_dat_o[16]
rlabel metal3 192640 24472 192640 24472 0 wbs_dat_o[17]
rlabel metal2 240296 36008 240296 36008 0 wbs_dat_o[18]
rlabel metal2 142856 7518 142856 7518 0 wbs_dat_o[19]
rlabel metal3 350056 205478 350056 205478 0 wbs_dat_o[1]
rlabel metal2 148456 13398 148456 13398 0 wbs_dat_o[20]
rlabel metal2 242984 36792 242984 36792 0 wbs_dat_o[21]
rlabel metal4 349944 35000 349944 35000 0 wbs_dat_o[22]
rlabel metal2 165816 4046 165816 4046 0 wbs_dat_o[23]
rlabel metal2 171416 12894 171416 12894 0 wbs_dat_o[24]
rlabel metal4 350504 34776 350504 34776 0 wbs_dat_o[25]
rlabel metal2 349832 34776 349832 34776 0 wbs_dat_o[26]
rlabel metal2 239400 41328 239400 41328 0 wbs_dat_o[27]
rlabel metal2 242872 42672 242872 42672 0 wbs_dat_o[28]
rlabel metal2 171416 29162 171416 29162 0 wbs_dat_o[29]
rlabel metal3 130144 21224 130144 21224 0 wbs_dat_o[2]
rlabel metal2 169624 29050 169624 29050 0 wbs_dat_o[30]
rlabel metal2 167832 29106 167832 29106 0 wbs_dat_o[31]
rlabel metal2 49448 7406 49448 7406 0 wbs_dat_o[3]
rlabel metal2 57288 2310 57288 2310 0 wbs_dat_o[4]
rlabel metal2 214298 30072 214298 30072 0 wbs_dat_o[5]
rlabel metal2 212562 30072 212562 30072 0 wbs_dat_o[6]
rlabel metal2 74424 2702 74424 2702 0 wbs_dat_o[7]
rlabel metal2 209048 28938 209048 28938 0 wbs_dat_o[8]
rlabel metal2 207382 30072 207382 30072 0 wbs_dat_o[9]
rlabel metal2 28728 4046 28728 4046 0 wbs_sel_i[0]
rlabel metal2 117544 28840 117544 28840 0 wbs_sel_i[1]
rlabel metal2 43960 3150 43960 3150 0 wbs_sel_i[2]
rlabel metal2 51576 4102 51576 4102 0 wbs_sel_i[3]
rlabel metal3 585592 376600 585592 376600 0 wbs_stb_i
rlabel metal2 21112 462 21112 462 0 wbs_we_i
<< properties >>
string FIXED_BBOX 0 0 596040 596040
<< end >>
