VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO uart_i2c_usb_spi_top
  CLASS BLOCK ;
  FOREIGN uart_i2c_usb_spi_top ;
  ORIGIN 0.000 0.000 ;
  SIZE 850.000 BY 1000.000 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 19.940 15.380 26.140 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 119.940 15.380 126.140 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 219.940 15.380 226.140 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 319.940 15.380 326.140 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 419.940 15.380 426.140 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 519.940 15.380 526.140 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 619.940 15.380 626.140 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 719.940 15.380 726.140 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 819.940 15.380 826.140 984.220 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 69.940 15.380 76.140 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 169.940 15.380 176.140 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 269.940 15.380 276.140 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 369.940 15.380 376.140 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 469.940 15.380 476.140 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 569.940 15.380 576.140 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 669.940 15.380 676.140 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 769.940 15.380 776.140 984.220 ;
    END
  END VSS
  PIN app_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 85.120 4.000 85.680 ;
    END
  END app_clk
  PIN cfg_cska_uart[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 17.632000 ;
    ANTENNADIFFAREA 3.283200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 51.520 4.000 52.080 ;
    END
  END cfg_cska_uart[0]
  PIN cfg_cska_uart[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 8.816000 ;
    ANTENNADIFFAREA 1.641600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 40.320 4.000 40.880 ;
    END
  END cfg_cska_uart[1]
  PIN cfg_cska_uart[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.408000 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 29.120 4.000 29.680 ;
    END
  END cfg_cska_uart[2]
  PIN cfg_cska_uart[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 17.920 4.000 18.480 ;
    END
  END cfg_cska_uart[3]
  PIN i2c_rstn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 593.600 0.000 594.160 4.000 ;
    END
  END i2c_rstn
  PIN i2cm_intr_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 525.280 996.000 525.840 1000.000 ;
    END
  END i2cm_intr_o
  PIN reg_ack
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 981.120 4.000 981.680 ;
    END
  END reg_ack
  PIN reg_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 208.320 4.000 208.880 ;
    END
  END reg_addr[0]
  PIN reg_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 197.120 4.000 197.680 ;
    END
  END reg_addr[1]
  PIN reg_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 185.920 4.000 186.480 ;
    END
  END reg_addr[2]
  PIN reg_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 174.720 4.000 175.280 ;
    END
  END reg_addr[3]
  PIN reg_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 163.520 4.000 164.080 ;
    END
  END reg_addr[4]
  PIN reg_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 152.320 4.000 152.880 ;
    END
  END reg_addr[5]
  PIN reg_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 141.120 4.000 141.680 ;
    END
  END reg_addr[6]
  PIN reg_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 129.920 4.000 130.480 ;
    END
  END reg_addr[7]
  PIN reg_addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 118.720 4.000 119.280 ;
    END
  END reg_addr[8]
  PIN reg_be[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 253.120 4.000 253.680 ;
    END
  END reg_be[0]
  PIN reg_be[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 241.920 4.000 242.480 ;
    END
  END reg_be[1]
  PIN reg_be[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 230.720 4.000 231.280 ;
    END
  END reg_be[2]
  PIN reg_be[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 219.520 4.000 220.080 ;
    END
  END reg_be[3]
  PIN reg_cs
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 96.320 4.000 96.880 ;
    END
  END reg_cs
  PIN reg_rdata[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 969.920 4.000 970.480 ;
    END
  END reg_rdata[0]
  PIN reg_rdata[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 857.920 4.000 858.480 ;
    END
  END reg_rdata[10]
  PIN reg_rdata[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 846.720 4.000 847.280 ;
    END
  END reg_rdata[11]
  PIN reg_rdata[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 835.520 4.000 836.080 ;
    END
  END reg_rdata[12]
  PIN reg_rdata[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 824.320 4.000 824.880 ;
    END
  END reg_rdata[13]
  PIN reg_rdata[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 813.120 4.000 813.680 ;
    END
  END reg_rdata[14]
  PIN reg_rdata[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 801.920 4.000 802.480 ;
    END
  END reg_rdata[15]
  PIN reg_rdata[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 790.720 4.000 791.280 ;
    END
  END reg_rdata[16]
  PIN reg_rdata[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 779.520 4.000 780.080 ;
    END
  END reg_rdata[17]
  PIN reg_rdata[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 768.320 4.000 768.880 ;
    END
  END reg_rdata[18]
  PIN reg_rdata[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 757.120 4.000 757.680 ;
    END
  END reg_rdata[19]
  PIN reg_rdata[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 958.720 4.000 959.280 ;
    END
  END reg_rdata[1]
  PIN reg_rdata[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 745.920 4.000 746.480 ;
    END
  END reg_rdata[20]
  PIN reg_rdata[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 734.720 4.000 735.280 ;
    END
  END reg_rdata[21]
  PIN reg_rdata[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 723.520 4.000 724.080 ;
    END
  END reg_rdata[22]
  PIN reg_rdata[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 712.320 4.000 712.880 ;
    END
  END reg_rdata[23]
  PIN reg_rdata[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 701.120 4.000 701.680 ;
    END
  END reg_rdata[24]
  PIN reg_rdata[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 689.920 4.000 690.480 ;
    END
  END reg_rdata[25]
  PIN reg_rdata[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 678.720 4.000 679.280 ;
    END
  END reg_rdata[26]
  PIN reg_rdata[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 667.520 4.000 668.080 ;
    END
  END reg_rdata[27]
  PIN reg_rdata[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 656.320 4.000 656.880 ;
    END
  END reg_rdata[28]
  PIN reg_rdata[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 645.120 4.000 645.680 ;
    END
  END reg_rdata[29]
  PIN reg_rdata[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 947.520 4.000 948.080 ;
    END
  END reg_rdata[2]
  PIN reg_rdata[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 633.920 4.000 634.480 ;
    END
  END reg_rdata[30]
  PIN reg_rdata[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 622.720 4.000 623.280 ;
    END
  END reg_rdata[31]
  PIN reg_rdata[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 936.320 4.000 936.880 ;
    END
  END reg_rdata[3]
  PIN reg_rdata[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 925.120 4.000 925.680 ;
    END
  END reg_rdata[4]
  PIN reg_rdata[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 913.920 4.000 914.480 ;
    END
  END reg_rdata[5]
  PIN reg_rdata[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 902.720 4.000 903.280 ;
    END
  END reg_rdata[6]
  PIN reg_rdata[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 891.520 4.000 892.080 ;
    END
  END reg_rdata[7]
  PIN reg_rdata[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 880.320 4.000 880.880 ;
    END
  END reg_rdata[8]
  PIN reg_rdata[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 869.120 4.000 869.680 ;
    END
  END reg_rdata[9]
  PIN reg_wdata[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 611.520 4.000 612.080 ;
    END
  END reg_wdata[0]
  PIN reg_wdata[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 499.520 4.000 500.080 ;
    END
  END reg_wdata[10]
  PIN reg_wdata[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 488.320 4.000 488.880 ;
    END
  END reg_wdata[11]
  PIN reg_wdata[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 477.120 4.000 477.680 ;
    END
  END reg_wdata[12]
  PIN reg_wdata[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 465.920 4.000 466.480 ;
    END
  END reg_wdata[13]
  PIN reg_wdata[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 454.720 4.000 455.280 ;
    END
  END reg_wdata[14]
  PIN reg_wdata[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 443.520 4.000 444.080 ;
    END
  END reg_wdata[15]
  PIN reg_wdata[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 432.320 4.000 432.880 ;
    END
  END reg_wdata[16]
  PIN reg_wdata[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 421.120 4.000 421.680 ;
    END
  END reg_wdata[17]
  PIN reg_wdata[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 409.920 4.000 410.480 ;
    END
  END reg_wdata[18]
  PIN reg_wdata[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 398.720 4.000 399.280 ;
    END
  END reg_wdata[19]
  PIN reg_wdata[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 600.320 4.000 600.880 ;
    END
  END reg_wdata[1]
  PIN reg_wdata[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 387.520 4.000 388.080 ;
    END
  END reg_wdata[20]
  PIN reg_wdata[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 376.320 4.000 376.880 ;
    END
  END reg_wdata[21]
  PIN reg_wdata[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 365.120 4.000 365.680 ;
    END
  END reg_wdata[22]
  PIN reg_wdata[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 353.920 4.000 354.480 ;
    END
  END reg_wdata[23]
  PIN reg_wdata[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 342.720 4.000 343.280 ;
    END
  END reg_wdata[24]
  PIN reg_wdata[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 331.520 4.000 332.080 ;
    END
  END reg_wdata[25]
  PIN reg_wdata[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 320.320 4.000 320.880 ;
    END
  END reg_wdata[26]
  PIN reg_wdata[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 309.120 4.000 309.680 ;
    END
  END reg_wdata[27]
  PIN reg_wdata[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 297.920 4.000 298.480 ;
    END
  END reg_wdata[28]
  PIN reg_wdata[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 286.720 4.000 287.280 ;
    END
  END reg_wdata[29]
  PIN reg_wdata[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 589.120 4.000 589.680 ;
    END
  END reg_wdata[2]
  PIN reg_wdata[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 275.520 4.000 276.080 ;
    END
  END reg_wdata[30]
  PIN reg_wdata[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 264.320 4.000 264.880 ;
    END
  END reg_wdata[31]
  PIN reg_wdata[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 577.920 4.000 578.480 ;
    END
  END reg_wdata[3]
  PIN reg_wdata[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 566.720 4.000 567.280 ;
    END
  END reg_wdata[4]
  PIN reg_wdata[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 555.520 4.000 556.080 ;
    END
  END reg_wdata[5]
  PIN reg_wdata[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 544.320 4.000 544.880 ;
    END
  END reg_wdata[6]
  PIN reg_wdata[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 533.120 4.000 533.680 ;
    END
  END reg_wdata[7]
  PIN reg_wdata[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 521.920 4.000 522.480 ;
    END
  END reg_wdata[8]
  PIN reg_wdata[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 510.720 4.000 511.280 ;
    END
  END reg_wdata[9]
  PIN reg_wr
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 107.520 4.000 108.080 ;
    END
  END reg_wr
  PIN scl_pad_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 21.280 996.000 21.840 1000.000 ;
    END
  END scl_pad_i
  PIN scl_pad_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 54.880 996.000 55.440 1000.000 ;
    END
  END scl_pad_o
  PIN scl_pad_oen_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 88.480 996.000 89.040 1000.000 ;
    END
  END scl_pad_oen_o
  PIN sda_pad_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 122.080 996.000 122.640 1000.000 ;
    END
  END sda_pad_i
  PIN sda_pad_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 155.680 996.000 156.240 1000.000 ;
    END
  END sda_pad_o
  PIN sda_padoen_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 189.280 996.000 189.840 1000.000 ;
    END
  END sda_padoen_o
  PIN spi_rstn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 592.480 996.000 593.040 1000.000 ;
    END
  END spi_rstn
  PIN sspim_sck
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 626.080 996.000 626.640 1000.000 ;
    END
  END sspim_sck
  PIN sspim_si
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 659.680 996.000 660.240 1000.000 ;
    END
  END sspim_si
  PIN sspim_so
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 693.280 996.000 693.840 1000.000 ;
    END
  END sspim_so
  PIN sspim_ssn[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 827.680 996.000 828.240 1000.000 ;
    END
  END sspim_ssn[0]
  PIN sspim_ssn[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 794.080 996.000 794.640 1000.000 ;
    END
  END sspim_ssn[1]
  PIN sspim_ssn[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 760.480 996.000 761.040 1000.000 ;
    END
  END sspim_ssn[2]
  PIN sspim_ssn[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 726.880 996.000 727.440 1000.000 ;
    END
  END sspim_ssn[3]
  PIN uart_rstn[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 424.480 0.000 425.040 4.000 ;
    END
  END uart_rstn[0]
  PIN uart_rstn[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 255.360 0.000 255.920 4.000 ;
    END
  END uart_rstn[1]
  PIN uart_rxd[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 222.880 996.000 223.440 1000.000 ;
    END
  END uart_rxd[0]
  PIN uart_rxd[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 290.080 996.000 290.640 1000.000 ;
    END
  END uart_rxd[1]
  PIN uart_txd[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 256.480 996.000 257.040 1000.000 ;
    END
  END uart_txd[0]
  PIN uart_txd[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal2 ;
        RECT 323.680 996.000 324.240 1000.000 ;
    END
  END uart_txd[1]
  PIN usb_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 86.240 0.000 86.800 4.000 ;
    END
  END usb_clk
  PIN usb_in_dn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 390.880 996.000 391.440 1000.000 ;
    END
  END usb_in_dn
  PIN usb_in_dp
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 357.280 996.000 357.840 1000.000 ;
    END
  END usb_in_dp
  PIN usb_intr_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 558.880 996.000 559.440 1000.000 ;
    END
  END usb_intr_o
  PIN usb_out_dn
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal2 ;
        RECT 458.080 996.000 458.640 1000.000 ;
    END
  END usb_out_dn
  PIN usb_out_dp
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 424.480 996.000 425.040 1000.000 ;
    END
  END usb_out_dp
  PIN usb_out_tx_oen
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 491.680 996.000 492.240 1000.000 ;
    END
  END usb_out_tx_oen
  PIN usb_rstn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 762.720 0.000 763.280 4.000 ;
    END
  END usb_rstn
  PIN wbd_clk_int
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 62.720 4.000 63.280 ;
    END
  END wbd_clk_int
  PIN wbd_clk_uart
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 73.920 4.000 74.480 ;
    END
  END wbd_clk_uart
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 842.800 984.890 ;
      LAYER Metal2 ;
        RECT 7.420 995.700 20.980 996.660 ;
        RECT 22.140 995.700 54.580 996.660 ;
        RECT 55.740 995.700 88.180 996.660 ;
        RECT 89.340 995.700 121.780 996.660 ;
        RECT 122.940 995.700 155.380 996.660 ;
        RECT 156.540 995.700 188.980 996.660 ;
        RECT 190.140 995.700 222.580 996.660 ;
        RECT 223.740 995.700 256.180 996.660 ;
        RECT 257.340 995.700 289.780 996.660 ;
        RECT 290.940 995.700 323.380 996.660 ;
        RECT 324.540 995.700 356.980 996.660 ;
        RECT 358.140 995.700 390.580 996.660 ;
        RECT 391.740 995.700 424.180 996.660 ;
        RECT 425.340 995.700 457.780 996.660 ;
        RECT 458.940 995.700 491.380 996.660 ;
        RECT 492.540 995.700 524.980 996.660 ;
        RECT 526.140 995.700 558.580 996.660 ;
        RECT 559.740 995.700 592.180 996.660 ;
        RECT 593.340 995.700 625.780 996.660 ;
        RECT 626.940 995.700 659.380 996.660 ;
        RECT 660.540 995.700 692.980 996.660 ;
        RECT 694.140 995.700 726.580 996.660 ;
        RECT 727.740 995.700 760.180 996.660 ;
        RECT 761.340 995.700 793.780 996.660 ;
        RECT 794.940 995.700 827.380 996.660 ;
        RECT 828.540 995.700 841.540 996.660 ;
        RECT 7.420 4.300 841.540 995.700 ;
        RECT 7.420 4.000 85.940 4.300 ;
        RECT 87.100 4.000 255.060 4.300 ;
        RECT 256.220 4.000 424.180 4.300 ;
        RECT 425.340 4.000 593.300 4.300 ;
        RECT 594.460 4.000 762.420 4.300 ;
        RECT 763.580 4.000 841.540 4.300 ;
      LAYER Metal3 ;
        RECT 3.500 981.980 841.590 984.900 ;
        RECT 4.300 980.820 841.590 981.980 ;
        RECT 3.500 970.780 841.590 980.820 ;
        RECT 4.300 969.620 841.590 970.780 ;
        RECT 3.500 959.580 841.590 969.620 ;
        RECT 4.300 958.420 841.590 959.580 ;
        RECT 3.500 948.380 841.590 958.420 ;
        RECT 4.300 947.220 841.590 948.380 ;
        RECT 3.500 937.180 841.590 947.220 ;
        RECT 4.300 936.020 841.590 937.180 ;
        RECT 3.500 925.980 841.590 936.020 ;
        RECT 4.300 924.820 841.590 925.980 ;
        RECT 3.500 914.780 841.590 924.820 ;
        RECT 4.300 913.620 841.590 914.780 ;
        RECT 3.500 903.580 841.590 913.620 ;
        RECT 4.300 902.420 841.590 903.580 ;
        RECT 3.500 892.380 841.590 902.420 ;
        RECT 4.300 891.220 841.590 892.380 ;
        RECT 3.500 881.180 841.590 891.220 ;
        RECT 4.300 880.020 841.590 881.180 ;
        RECT 3.500 869.980 841.590 880.020 ;
        RECT 4.300 868.820 841.590 869.980 ;
        RECT 3.500 858.780 841.590 868.820 ;
        RECT 4.300 857.620 841.590 858.780 ;
        RECT 3.500 847.580 841.590 857.620 ;
        RECT 4.300 846.420 841.590 847.580 ;
        RECT 3.500 836.380 841.590 846.420 ;
        RECT 4.300 835.220 841.590 836.380 ;
        RECT 3.500 825.180 841.590 835.220 ;
        RECT 4.300 824.020 841.590 825.180 ;
        RECT 3.500 813.980 841.590 824.020 ;
        RECT 4.300 812.820 841.590 813.980 ;
        RECT 3.500 802.780 841.590 812.820 ;
        RECT 4.300 801.620 841.590 802.780 ;
        RECT 3.500 791.580 841.590 801.620 ;
        RECT 4.300 790.420 841.590 791.580 ;
        RECT 3.500 780.380 841.590 790.420 ;
        RECT 4.300 779.220 841.590 780.380 ;
        RECT 3.500 769.180 841.590 779.220 ;
        RECT 4.300 768.020 841.590 769.180 ;
        RECT 3.500 757.980 841.590 768.020 ;
        RECT 4.300 756.820 841.590 757.980 ;
        RECT 3.500 746.780 841.590 756.820 ;
        RECT 4.300 745.620 841.590 746.780 ;
        RECT 3.500 735.580 841.590 745.620 ;
        RECT 4.300 734.420 841.590 735.580 ;
        RECT 3.500 724.380 841.590 734.420 ;
        RECT 4.300 723.220 841.590 724.380 ;
        RECT 3.500 713.180 841.590 723.220 ;
        RECT 4.300 712.020 841.590 713.180 ;
        RECT 3.500 701.980 841.590 712.020 ;
        RECT 4.300 700.820 841.590 701.980 ;
        RECT 3.500 690.780 841.590 700.820 ;
        RECT 4.300 689.620 841.590 690.780 ;
        RECT 3.500 679.580 841.590 689.620 ;
        RECT 4.300 678.420 841.590 679.580 ;
        RECT 3.500 668.380 841.590 678.420 ;
        RECT 4.300 667.220 841.590 668.380 ;
        RECT 3.500 657.180 841.590 667.220 ;
        RECT 4.300 656.020 841.590 657.180 ;
        RECT 3.500 645.980 841.590 656.020 ;
        RECT 4.300 644.820 841.590 645.980 ;
        RECT 3.500 634.780 841.590 644.820 ;
        RECT 4.300 633.620 841.590 634.780 ;
        RECT 3.500 623.580 841.590 633.620 ;
        RECT 4.300 622.420 841.590 623.580 ;
        RECT 3.500 612.380 841.590 622.420 ;
        RECT 4.300 611.220 841.590 612.380 ;
        RECT 3.500 601.180 841.590 611.220 ;
        RECT 4.300 600.020 841.590 601.180 ;
        RECT 3.500 589.980 841.590 600.020 ;
        RECT 4.300 588.820 841.590 589.980 ;
        RECT 3.500 578.780 841.590 588.820 ;
        RECT 4.300 577.620 841.590 578.780 ;
        RECT 3.500 567.580 841.590 577.620 ;
        RECT 4.300 566.420 841.590 567.580 ;
        RECT 3.500 556.380 841.590 566.420 ;
        RECT 4.300 555.220 841.590 556.380 ;
        RECT 3.500 545.180 841.590 555.220 ;
        RECT 4.300 544.020 841.590 545.180 ;
        RECT 3.500 533.980 841.590 544.020 ;
        RECT 4.300 532.820 841.590 533.980 ;
        RECT 3.500 522.780 841.590 532.820 ;
        RECT 4.300 521.620 841.590 522.780 ;
        RECT 3.500 511.580 841.590 521.620 ;
        RECT 4.300 510.420 841.590 511.580 ;
        RECT 3.500 500.380 841.590 510.420 ;
        RECT 4.300 499.220 841.590 500.380 ;
        RECT 3.500 489.180 841.590 499.220 ;
        RECT 4.300 488.020 841.590 489.180 ;
        RECT 3.500 477.980 841.590 488.020 ;
        RECT 4.300 476.820 841.590 477.980 ;
        RECT 3.500 466.780 841.590 476.820 ;
        RECT 4.300 465.620 841.590 466.780 ;
        RECT 3.500 455.580 841.590 465.620 ;
        RECT 4.300 454.420 841.590 455.580 ;
        RECT 3.500 444.380 841.590 454.420 ;
        RECT 4.300 443.220 841.590 444.380 ;
        RECT 3.500 433.180 841.590 443.220 ;
        RECT 4.300 432.020 841.590 433.180 ;
        RECT 3.500 421.980 841.590 432.020 ;
        RECT 4.300 420.820 841.590 421.980 ;
        RECT 3.500 410.780 841.590 420.820 ;
        RECT 4.300 409.620 841.590 410.780 ;
        RECT 3.500 399.580 841.590 409.620 ;
        RECT 4.300 398.420 841.590 399.580 ;
        RECT 3.500 388.380 841.590 398.420 ;
        RECT 4.300 387.220 841.590 388.380 ;
        RECT 3.500 377.180 841.590 387.220 ;
        RECT 4.300 376.020 841.590 377.180 ;
        RECT 3.500 365.980 841.590 376.020 ;
        RECT 4.300 364.820 841.590 365.980 ;
        RECT 3.500 354.780 841.590 364.820 ;
        RECT 4.300 353.620 841.590 354.780 ;
        RECT 3.500 343.580 841.590 353.620 ;
        RECT 4.300 342.420 841.590 343.580 ;
        RECT 3.500 332.380 841.590 342.420 ;
        RECT 4.300 331.220 841.590 332.380 ;
        RECT 3.500 321.180 841.590 331.220 ;
        RECT 4.300 320.020 841.590 321.180 ;
        RECT 3.500 309.980 841.590 320.020 ;
        RECT 4.300 308.820 841.590 309.980 ;
        RECT 3.500 298.780 841.590 308.820 ;
        RECT 4.300 297.620 841.590 298.780 ;
        RECT 3.500 287.580 841.590 297.620 ;
        RECT 4.300 286.420 841.590 287.580 ;
        RECT 3.500 276.380 841.590 286.420 ;
        RECT 4.300 275.220 841.590 276.380 ;
        RECT 3.500 265.180 841.590 275.220 ;
        RECT 4.300 264.020 841.590 265.180 ;
        RECT 3.500 253.980 841.590 264.020 ;
        RECT 4.300 252.820 841.590 253.980 ;
        RECT 3.500 242.780 841.590 252.820 ;
        RECT 4.300 241.620 841.590 242.780 ;
        RECT 3.500 231.580 841.590 241.620 ;
        RECT 4.300 230.420 841.590 231.580 ;
        RECT 3.500 220.380 841.590 230.420 ;
        RECT 4.300 219.220 841.590 220.380 ;
        RECT 3.500 209.180 841.590 219.220 ;
        RECT 4.300 208.020 841.590 209.180 ;
        RECT 3.500 197.980 841.590 208.020 ;
        RECT 4.300 196.820 841.590 197.980 ;
        RECT 3.500 186.780 841.590 196.820 ;
        RECT 4.300 185.620 841.590 186.780 ;
        RECT 3.500 175.580 841.590 185.620 ;
        RECT 4.300 174.420 841.590 175.580 ;
        RECT 3.500 164.380 841.590 174.420 ;
        RECT 4.300 163.220 841.590 164.380 ;
        RECT 3.500 153.180 841.590 163.220 ;
        RECT 4.300 152.020 841.590 153.180 ;
        RECT 3.500 141.980 841.590 152.020 ;
        RECT 4.300 140.820 841.590 141.980 ;
        RECT 3.500 130.780 841.590 140.820 ;
        RECT 4.300 129.620 841.590 130.780 ;
        RECT 3.500 119.580 841.590 129.620 ;
        RECT 4.300 118.420 841.590 119.580 ;
        RECT 3.500 108.380 841.590 118.420 ;
        RECT 4.300 107.220 841.590 108.380 ;
        RECT 3.500 97.180 841.590 107.220 ;
        RECT 4.300 96.020 841.590 97.180 ;
        RECT 3.500 85.980 841.590 96.020 ;
        RECT 4.300 84.820 841.590 85.980 ;
        RECT 3.500 74.780 841.590 84.820 ;
        RECT 4.300 73.620 841.590 74.780 ;
        RECT 3.500 63.580 841.590 73.620 ;
        RECT 4.300 62.420 841.590 63.580 ;
        RECT 3.500 52.380 841.590 62.420 ;
        RECT 4.300 51.220 841.590 52.380 ;
        RECT 3.500 41.180 841.590 51.220 ;
        RECT 4.300 40.020 841.590 41.180 ;
        RECT 3.500 29.980 841.590 40.020 ;
        RECT 4.300 28.820 841.590 29.980 ;
        RECT 3.500 18.780 841.590 28.820 ;
        RECT 4.300 17.620 841.590 18.780 ;
        RECT 3.500 15.540 841.590 17.620 ;
      LAYER Metal4 ;
        RECT 9.660 20.810 19.640 981.030 ;
        RECT 26.440 20.810 69.640 981.030 ;
        RECT 76.440 20.810 119.640 981.030 ;
        RECT 126.440 20.810 169.640 981.030 ;
        RECT 176.440 20.810 219.640 981.030 ;
        RECT 226.440 20.810 269.640 981.030 ;
        RECT 276.440 20.810 319.640 981.030 ;
        RECT 326.440 20.810 369.640 981.030 ;
        RECT 376.440 20.810 419.640 981.030 ;
        RECT 426.440 20.810 469.640 981.030 ;
        RECT 476.440 20.810 519.640 981.030 ;
        RECT 526.440 20.810 569.640 981.030 ;
        RECT 576.440 20.810 619.640 981.030 ;
        RECT 626.440 20.810 669.640 981.030 ;
        RECT 676.440 20.810 719.640 981.030 ;
        RECT 726.440 20.810 769.640 981.030 ;
        RECT 776.440 20.810 819.640 981.030 ;
        RECT 826.440 20.810 838.180 981.030 ;
      LAYER Metal5 ;
        RECT 13.500 47.930 832.100 887.170 ;
  END
END uart_i2c_usb_spi_top
END LIBRARY

