* NGSPICE file created from temp_sensor.ext - technology: gf180mcuD

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_2 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_4 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_4 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_4 A1 A2 A3 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_4 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_3 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_2 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_2 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__invz_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__invz_2 EN I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_1 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_4 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__invz_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__invz_4 EN I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__invz_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__invz_1 EN I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_4 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_2 A1 A2 A3 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__invz_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__invz_3 EN I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_2 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_2 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_4 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_2 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_4 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_4 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_2 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_1 A1 A2 A3 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_4 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_2 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_4 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_4 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tiel abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tiel ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_12 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_12 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_8 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_12 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_12 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_2 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_2 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_2 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_8 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_12 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_12 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_4 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_4 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_2 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_4 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_1 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_8 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_3 I Z VDD VNW VPW VSS
.ends

.subckt temp_sensor VDD VSS io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6]
+ io_out[7]
XFILLER_0_27_60 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_4 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_188 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1206__A1 _0346_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_288 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_269 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_68_581 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1724__CLK net11 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xdec1._061_ dec1.i_tens dec1._001_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_55_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_199 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_15 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_temp1.dac.parallel_cells\[0\].vdac_batch.einvp_batch\[0\].vref_I temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1270_ net25 _0684_ _0778_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_64_14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_155 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_136 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_158 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_214 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_350 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0985_ _0509_ _0407_ _0408_ _0510_ _0511_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_0_14_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_383 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_66 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1606_ ctr\[3\] clknet_1_0__leaf__0318_ _0320_ _0193_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__0962__A3 _0440_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_4 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1537_ _0782_ _0294_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_1468_ _0522_ _0791_ _0111_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1399_ _0236_ _0070_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_57_518 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1747__CLK net12 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_65_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_252 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_191 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_88_687 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_239 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xdec1._113_ dec1._047_ dec1._040_ dec1._051_ dec1._039_ dec1._002_ dec1._052_ VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_36_350 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1322_ cal_lut\[28\] _0780_ _0801_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_75_35 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_75_24 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1253_ _0704_ _0762_ _0763_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1184_ _0689_ _0690_ _0695_ _0698_ _0699_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__1621__B ctr\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_62_543 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_255 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0968_ _0455_ _0460_ _0494_ _0433_ cal_lut\[2\] _0495_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai32_4
X_0899_ _0358_ _0365_ _0356_ _0413_ _0427_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_64_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_283 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0871__A2 _0395_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_401 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_18_361 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_297 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_397 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_76_624 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0836__I _0363_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_136 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0822_ ctr\[9\] ctr\[8\] _0351_ _0352_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_9_27 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_203 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_331 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_364 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0917__A3 _0355_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_45 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_78 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_61 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1305_ _0794_ _0017_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1236_ _0697_ _0746_ _0747_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1167_ net5 _0682_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_3
X_1098_ cal_lut\[65\] _0622_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_74_220 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_312 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1030__A2 _0407_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[3\].vref_I temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_dec1._090__A1 dec1.i_bin\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_73_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_201 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_117 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_25_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_286 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_191 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_109 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_278 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1021__A2 _0377_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_356 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_0_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_56_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1021_ cal_lut\[58\] _0377_ _0379_ cal_lut\[64\] _0546_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__1808__CLK net15 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_401 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_88_378 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_264 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1854_ _0206_ clknet_1_1__leaf_io_in[0] ctr\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_21_95 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1785_ _0137_ net12 cal_lut\[138\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_97_33 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1012__A2 _0512_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_dec1._072__A1 dec1.i_bin\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1219_ _0728_ _0729_ _0731_ clknet_1_1__leaf_io_in[0] io_out[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_47_220 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_35_395 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_286 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1490__A2 _0255_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_28 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_348 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1242__A2 _0709_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_278 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1570_ _0531_ _0289_ _0171_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_21_153 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_39 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtemp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[6\].pupd temp1.dac.parallel_cells\[3\].vdac_batch.en_pupd
+ temp1.dac.parallel_cells\[3\].vdac_batch.npu_pd temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__invz_2
XTAP_TAPCELL_ROW_1_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_92_711 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_49_476 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtemp1.dac.parallel_cells\[2\].vdac_batch._4_ temp1.dac.i_data\[2\] temp1.dac.i_data\[5\]
+ temp1.dac.parallel_cells\[2\].vdac_batch._1_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__1780__CLK net8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1004_ _0528_ _0436_ _0529_ _0530_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_32_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_381 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_94 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1837_ _0189_ net10 cal_lut\[190\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__0992__A1 _0360_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_153 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1768_ _0120_ net12 cal_lut\[121\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1699_ _0051_ net17 cal_lut\[52\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_79_131 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_304 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1472__A2 _0240_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_186 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_23_332 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_381 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_90_373 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_267 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1653__CLK net11 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1160__A1 ctr\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_46_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtemp1.dac.vdac_single._4_ net20 net21 temp1.dac.vdac_single._1_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_5_128 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_340 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0974__A1 _0360_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1622_ _0348_ _0327_ _0783_ _0202_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1553_ _0560_ _0289_ _0160_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1484_ cal_lut\[120\] _0240_ _0272_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__1624__B _0783_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_50 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1151__A1 _0346_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[6\].vref_I temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1454__A2 _0240_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_82 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_201 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_20_313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_245 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xtemp1.dac.vdac_single.einvp_batch\[0\].pupd temp1.dac.vdac_single.en_pupd temp1.dac.vdac_single.npu_pd
+ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__invz_2
XFILLER_0_94_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_373 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1676__CLK net11 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xdec1._060_ dec1.i_bin\[0\] dec1._000_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_55_307 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_381 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_204 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_384 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_80_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1699__CLK net17 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_373 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0984_ cal_lut\[21\] _0510_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__0947__A1 _0360_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1605_ _0365_ clknet_1_0__leaf__0318_ _0782_ _0320_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_1_153 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1536_ _0293_ _0150_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1467_ _0478_ _0790_ _0110_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1398_ cal_lut\[70\] _0802_ _0236_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_57_519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0883__B1 _0403_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_229 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_65_563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_292 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1427__A2 _0791_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_242 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_220 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_310 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_321 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_170 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_88_688 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xdec1._112_ dec1._047_ dec1._050_ dec1._051_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__1841__CLK clknet_1_0__leaf_io_in[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1418__A2 _0791_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__0929__A1 _0360_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_384 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1354__A1 cal_lut\[47\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1321_ _0800_ _0027_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1106__A1 _0368_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1252_ _0585_ _0687_ _0760_ _0761_ _0762_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1183_ _0696_ _0697_ _0690_ _0698_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1409__A2 _0240_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0880__A3 _0406_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xtemp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[11\].pupd temp1.dac.parallel_cells\[4\].vdac_batch.en_pupd
+ temp1.dac.parallel_cells\[4\].vdac_batch.npu_pd temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__invz_2
XFILLER_0_24_73 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_62_544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_284 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_181 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0967_ _0464_ _0468_ _0481_ _0493_ _0494_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XPHY_EDGE_ROW_12_Right_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_42_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0898_ cal_lut\[109\] _0426_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_10_240 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1714__CLK net9 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_273 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1519_ _0608_ _0289_ _0137_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_65_80 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_207 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_21_Right_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_77_273 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_373 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_30_Right_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_60_195 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_76_625 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_14_Left_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_28_148 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_416 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_276 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_321 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0821_ _0344_ _0350_ _0351_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_43_129 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_298 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_23_Left_121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_24_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1737__CLK net16 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_86 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1304_ cal_lut\[17\] _0780_ _0794_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1235_ seg1.o_segments\[4\] _0691_ _0746_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_32_Left_130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1166_ net7 _0681_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_35_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1097_ _0611_ _0614_ _0617_ _0620_ _0621_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_0_19_137 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_126 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1263__B1 _0770_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_310 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_129 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1566__A1 cal_lut\[168\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0908__A4 _0391_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_184 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_2_281 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_73_606 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0844__A3 _0367_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_81_650 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_416 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_298 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_213 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_302 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_173 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_346 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_27 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1020_ _0368_ cal_lut\[130\] _0373_ _0545_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_88_346 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_56_221 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1853_ _0205_ clknet_1_1__leaf_io_in[0] ctr\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_12_271 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_235 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1784_ _0136_ net10 cal_lut\[137\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xfanout8 net13 net8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_12_313 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_195 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1012__A3 _0525_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_379 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_4_228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_82 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1218_ _0680_ _0730_ _0731_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_94_305 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1149_ _0670_ _0671_ dec1.i_bin\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XTAP_TAPCELL_ROW_35_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_92 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1003__A3 _0391_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_18 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_257 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_165 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_1_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_92_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_30 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1003_ _0376_ cal_lut\[99\] _0391_ _0413_ _0529_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
Xtemp1.dac.parallel_cells\[2\].vdac_batch._3_ temp1.dac.i_data\[2\] temp1.dac.parallel_cells\[2\].vdac_batch.npu_pd
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_88_187 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_254 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_276 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_298 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_224 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1836_ _0188_ net10 cal_lut\[189\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_6_Right_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_4_310 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_365 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1767_ _0119_ net12 cal_lut\[120\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_4_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_12_165 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1698_ _0050_ net17 cal_lut\[51\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_73_80 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_338 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xtemp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[6\].vref temp1.dac.parallel_cells\[3\].vdac_batch.en_vref
+ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__invz_4
XTAP_TAPCELL_ROW_23_333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_202 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_192 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_50_238 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_46_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_371 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtemp1.dac.vdac_single._3_ net19 temp1.dac.vdac_single.npu_pd VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_93_190 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_59_Right_59 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_14_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1621_ ctr\[2\] _0347_ ctr\[3\] _0327_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_78_14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1552_ _0516_ _0289_ _0159_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1483_ _0271_ _0119_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input3_I io_in[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_68_Right_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_6_Left_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_76_124 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_43_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_319 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_179 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_77_Right_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_91_138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout8_I net13 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_268 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_257 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_205 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0965__A2 _0445_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_25_290 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1819_ _0171_ net14 cal_lut\[172\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_7_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_293 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1390__A2 _0802_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_86_Right_86 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_95_Right_95 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_43_439 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_483 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_171 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_193 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1770__CLK net10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xtemp1.dac.vdac_single.einvp_batch\[0\].vref temp1.dac.vdac_single.en_vref temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__invz_1
XANTENNA__1381__A2 _0805_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_79_Left_177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__0892__A1 _0360_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_39_360 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_168 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_88_Left_186 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_0983_ cal_lut\[45\] _0509_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_14_238 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_35 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1604_ ctr\[2\] clknet_1_1__leaf__0318_ _0319_ _0192_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1535_ cal_lut\[150\] _0255_ _0293_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XPHY_EDGE_ROW_97_Left_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1372__A2 _0805_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1466_ _0426_ _0791_ _0109_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1397_ _0235_ _0069_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_38_83 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_94 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1124__A2 _0440_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_65_564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_271 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_146 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtemp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[4\].pupd temp1.dac.parallel_cells\[4\].vdac_batch.en_pupd
+ temp1.dac.parallel_cells\[4\].vdac_batch.npu_pd temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__invz_2
XFILLER_0_45_330 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_45_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1793__CLK net13 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1060__A1 _0357_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_366 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1115__A2 _0357_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_88_689 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0874__A1 _0359_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xdec1._111_ dec1._048_ dec1._026_ dec1._049_ dec1._050_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_95_274 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_374 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_344 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_388 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1320_ cal_lut\[27\] _0783_ _0800_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__1354__A2 _0802_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1251_ _0345_ _0701_ _0687_ _0761_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1182_ _0681_ _0693_ _0697_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__1666__CLK net17 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_308 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_dec1._061__I dec1.i_tens VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_62_545 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_235 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_341 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_385 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_300 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_171 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0966_ _0483_ _0486_ _0489_ _0492_ _0493_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_42_355 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1042__A1 _0390_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1593__A2 _0782_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_0897_ _0376_ _0421_ _0422_ _0423_ _0424_ _0425_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai32_2
XANTENNA__1345__A2 _0791_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1518_ _0779_ _0289_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_1449_ _0258_ _0098_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__0856__A1 _0358_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_80 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_127 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_311 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtemp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[11\].vref temp1.dac.parallel_cells\[4\].vdac_batch.en_vref
+ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__invz_3
XANTENNA__1033__A1 _0359_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1336__A2 _0802_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_temp1.dac.vdac_single.einvp_batch\[0\].vref_I temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1689__CLK net16 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0847__A1 _0368_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_263 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_0820_ _0345_ ctr\[6\] _0349_ _0350_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_3_249 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1327__A2 _0802_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_30 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1303_ _0576_ _0791_ _0016_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1234_ _0357_ _0583_ _0691_ _0584_ _0745_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1165_ clknet_1_1__leaf_io_in[0] _0680_ _0678_ _0673_ temp1.i_precharge_n VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1096_ _0618_ _0436_ _0619_ _0620_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1263__A1 temp1.dac.i_enable VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_255 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1015__A1 _0357_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_314 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1566__A2 _0294_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_0949_ cal_lut\[86\] _0476_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_42_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1831__CLK net17 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_293 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1318__A2 _0783_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0829__A1 _0356_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_73_607 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_81_651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1254__A1 temp1.dac.i_data\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1557__A2 _0294_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_314 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_185 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1309__A2 _0790_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[6\].vref_I temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1704__CLK net8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_233 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_31 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1852_ _0204_ clknet_1_1__leaf_io_in[0] ctr\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_42 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_12_272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1783_ _0135_ net10 cal_lut\[136\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1548__A2 _0294_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1854__CLK clknet_1_1__leaf_io_in[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout9 net13 net9 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_12_347 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_4_229 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1217_ _0678_ _0684_ _0730_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_94_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1148_ cal_lut\[6\] _0433_ _0357_ _0671_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_1079_ cal_lut\[83\] _0602_ _0386_ cal_lut\[77\] _0603_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_35_397 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_233 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0995__B1 _0423_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_409 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_111 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1003__A4 _0413_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_144 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1727__CLK net16 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_380 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_51_Left_149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_53_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0986__B1 _0403_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_409 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_144 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_19 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_188 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_60_Left_158 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_92_713 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1002_ cal_lut\[147\] _0528_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_76_306 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_52 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_214 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0977__B1 _0386_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_300 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_378 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1835_ _0187_ net13 cal_lut\[188\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_4_333 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1766_ _0118_ net12 cal_lut\[119\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__0992__A3 _0378_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1697_ _0049_ net18 cal_lut\[50\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_32_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_103 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_328 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0968__B1 _0433_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_160 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_46_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_158 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_225 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_383 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1620__A1 _0783_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0974__A3 _0373_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_228 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1620_ _0783_ _0326_ _0201_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1_314 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_26 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1551_ _0472_ _0289_ _0158_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1482_ cal_lut\[119\] _0255_ _0271_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__1136__B1 _0402_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_74 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_62 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_236 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_191 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_20_315 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1611__A1 _0368_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1818_ _0170_ net14 cal_lut\[171\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_4_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1749_ _0101_ net10 cal_lut\[102\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_68_70 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_67_158 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_350 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_169 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_51_484 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_342 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_103 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_temp1.dac.parallel_cells\[2\].vdac_batch._4__A2 temp1.dac.i_data\[5\] VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_136 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0982_ cal_lut\[165\] _0389_ _0392_ cal_lut\[123\] _0507_ _0508_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_13_43 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_342 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0947__A3 _0378_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1603_ _0355_ clknet_1_1__leaf__0318_ _0782_ _0319_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1534_ _0618_ _0289_ _0149_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_59_7 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_51 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1465_ _0264_ _0108_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1396_ cal_lut\[69\] _0805_ _0235_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__0883__A2 _0402_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_200 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_266 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_80 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_56_510 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_220 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xdec1._110_ dec1._028_ dec1._034_ dec1._049_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__0929__A3 _0373_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xtemp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[4\].vref temp1.dac.parallel_cells\[4\].vdac_batch.en_vref
+ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__invz_3
XFILLER_0_11_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1250_ _0757_ _0758_ _0759_ _0760_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1106__A3 _0373_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1181_ ctr\[2\] _0696_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
Xtemp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[3\].pupd temp1.dac.parallel_cells\[2\].vdac_batch.en_pupd
+ temp1.dac.parallel_cells\[2\].vdac_batch.npu_pd temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__invz_2
XFILLER_0_24_53 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_64 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_62_546 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_225 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_70_590 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_312 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_161 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0965_ _0490_ _0445_ _0491_ _0492_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__1042__A2 _0363_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_0896_ cal_lut\[85\] _0424_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_10_242 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1517_ _0288_ _0136_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1448_ cal_lut\[98\] _0255_ _0258_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1379_ cal_lut\[60\] _0802_ _0227_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__0856__A2 _0365_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1760__CLK net15 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_278 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_289 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_109 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_dec1._093__A1 dec1.i_bin\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_415 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_117 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_275 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_201 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_183 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_33 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_164 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_66 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_26 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1302_ _0532_ _0790_ _0015_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_dec1._084__A1 dec1.i_bin\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1233_ ctr\[6\] _0744_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__1783__CLK net10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1164_ _0346_ _0672_ _0680_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1095_ _0376_ cal_lut\[101\] _0391_ _0413_ _0619_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_19_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_128 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1263__A2 _0684_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_161 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout17_I net18 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_278 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0948_ cal_lut\[38\] _0475_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_30_304 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_164 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0879_ _0359_ _0390_ _0363_ _0406_ _0407_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_62_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__0829__A2 _0357_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_73_608 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_81_652 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1254__A2 _0709_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_131 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1656__CLK net16 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_dec1._066__A1 dec1.i_bin\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1190__A1 _0356_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_362 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_381 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_201 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1851_ _0203_ clknet_1_1__leaf_io_in[0] ctr\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_12_273 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1782_ _0134_ net10 cal_lut\[135\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1196__B _0684_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_36 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_12_337 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1216_ temp1.dac.i_data\[2\] _0709_ _0684_ _0729_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1147_ _0656_ _0662_ _0663_ _0669_ _0670_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
XFILLER_0_79_348 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1484__A2 _0240_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1078_ _0368_ _0365_ _0356_ _0401_ _0602_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
XTAP_TAPCELL_ROW_35_398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_278 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1679__CLK net8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0995__A1 _0376_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_101 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_189 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_temp1.dac.parallel_cells\[1\].vdac_batch._7__I temp1.dac.i_enable VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_278 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1163__A1 ctr\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xtemp1.dac._5_ temp1.dac._1_ temp1.dac.i_data\[5\] temp1.dac._0_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1001_ _0526_ _0432_ _0433_ _0527_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__1466__A2 _0791_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1821__CLK net14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_86 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_379 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_312 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1834_ _0186_ net12 cal_lut\[187\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xtemp1.dac.parallel_cells\[0\].vdac_batch._8_ temp1.dac.parallel_cells\[0\].vdac_batch._0_
+ temp1.dac.parallel_cells\[0\].vdac_batch._1_ temp1.dac.parallel_cells\[0\].vdac_batch.en_vref
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_12_112 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1765_ _0117_ net12 cal_lut\[118\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_145 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1696_ _0048_ net17 cal_lut\[49\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_189 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_321 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__0968__A1 _0455_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_226 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1090__B1 _0445_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1448__A2 _0255_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1844__CLK clknet_1_1__leaf_io_in[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_137 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_259 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_270 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_281 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1550_ _0417_ _0289_ _0157_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1481_ _0270_ _0118_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_94_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch._5__A1 temp1.dac.i_enable VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1439__A2 _0805_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_118 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_204 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_85 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_310 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_321 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_181 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_20_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1817_ _0169_ net14 cal_lut\[170\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_72_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1748_ _0100_ net12 cal_lut\[101\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1717__CLK net11 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1679_ _0031_ net8 cal_lut\[32\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_295 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_148 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_373 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_51_485 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_376 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_19 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_59_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0892__A3 _0378_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_148 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_362 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_159 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0981_ _0505_ _0395_ _0397_ _0506_ _0507_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_0_54_321 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_118 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_354 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1602_ _0317_ _0318_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_22_240 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_295 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1533_ _0572_ _0289_ _0148_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1464_ cal_lut\[108\] _0240_ _0264_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__1109__A1 _0433_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1395_ _0234_ _0068_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_9_234 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_45_354 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_72_162 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_398 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_60_357 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1348__A1 cal_lut\[42\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0859__B1 _0386_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0874__A3 _0401_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_416 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_321 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_36_354 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_181 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_302 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1180_ seg1.o_segments\[0\] _0691_ _0692_ _0694_ _0695_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_24_32 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_547 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1027__B1 _0392_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_0964_ _0376_ cal_lut\[116\] _0413_ _0406_ _0491_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XTAP_TAPCELL_ROW_70_591 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0895_ _0359_ _0365_ _0356_ _0385_ _0423_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_42_379 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1516_ cal_lut\[136\] _0255_ _0288_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_64_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_84 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_31 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1447_ _0257_ _0097_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1378_ _0612_ _0791_ _0059_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_65_61 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__0856__A3 _0355_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_298 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_82 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtemp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[3\].vref temp1.dac.parallel_cells\[2\].vdac_batch.en_vref
+ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__invz_3
XFILLER_0_18_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_18_365 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_335 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1033__A3 _0394_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_198 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0847__A3 _0373_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_243 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_224 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_162 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_45 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_49 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1301_ _0488_ _0790_ _0014_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1232_ net22 _0731_ _0742_ _0743_ io_out[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_35_42 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1163_ ctr\[7\] _0672_ _0679_ temp1.dac.i_data\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_1094_ cal_lut\[149\] _0618_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_35_53 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_90_697 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_324 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_173 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0947_ _0360_ _0472_ _0378_ _0418_ _0473_ _0474_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_0_82_290 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0878_ _0405_ _0406_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_2_251 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_416 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_140 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_279 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_205 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_195 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_29_363 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1850_ _0202_ clknet_1_1__leaf_io_in[0] ctr\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_21_33 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1781_ _0133_ net8 cal_lut\[134\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_24_121 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_77 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_305 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_360 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1750__CLK net10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1215_ _0363_ _0687_ _0726_ _0727_ _0704_ _0728_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_1_10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1146_ cal_lut\[12\] _0587_ _0664_ _0668_ _0669_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_1_87 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_47_202 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1077_ cal_lut\[89\] _0599_ _0600_ cal_lut\[23\] _0601_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[9\].vref_I temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xtemp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd temp1.dac.parallel_cells\[3\].vdac_batch.en_pupd
+ temp1.dac.parallel_cells\[3\].vdac_batch.npu_pd temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__invz_2
XTAP_TAPCELL_ROW_35_399 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_238 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1406__I _0779_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_3_220 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_308 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_38_213 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_26_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_216 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__0986__A2 _0402_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1773__CLK net10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_271 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_135 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_168 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_157 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xtemp1.dac._4_ temp1.dac.i_enable temp1.dac._1_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_16_33 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1000_ cal_lut\[141\] _0526_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_17_300 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_279 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_65 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_205 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0977__A2 _0383_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_76 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1833_ _0185_ net2 cal_lut\[186\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xtemp1.dac.parallel_cells\[0\].vdac_batch._7_ temp1.dac.i_enable temp1.dac.parallel_cells\[0\].vdac_batch._0_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_52_260 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1764_ _0116_ net14 cal_lut\[117\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_157 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1695_ _0047_ net18 cal_lut\[48\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_0_201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_73_50 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_73_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_79_135 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1129_ cal_lut\[96\] _0595_ _0377_ cal_lut\[60\] _0652_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_79_179 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_341 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_311 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1090__A1 _0376_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1796__CLK net12 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1090__B2 _0613_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_260 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1145__A2 _0666_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_19_Right_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_19_290 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1081__B2 cal_lut\[47\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1081__A1 cal_lut\[155\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_344 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_411 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_349 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_28_Right_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1480_ cal_lut\[118\] _0240_ _0270_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__1669__CLK net17 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0895__A1 _0359_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_37_406 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_37_Right_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_43_20 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_43_53 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_45_450 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_20_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_238 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1072__A1 _0368_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_46_Right_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1816_ _0168_ net14 cal_lut\[169\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_25_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_271 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_198 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1747_ _0099_ net12 cal_lut\[100\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1678_ _0030_ net11 cal_lut\[31\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1127__A2 _0386_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0886__A1 _0359_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_55_Right_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_67_138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_311 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_160 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_171 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_51_486 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1063__A1 _0360_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_64_Right_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_23_208 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_2_Left_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_31_241 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_39_Left_137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1366__A2 _0802_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1811__CLK net13 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1118__A2 _0395_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0877__A1 _0365_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_59_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_73_Right_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_48_Left_146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_39_330 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0980_ cal_lut\[105\] _0506_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_13_45 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_171 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_82_Right_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_6_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1054__A1 _0358_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_27 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1601_ temp_delay_last clknet_1_0__leaf__0316_ _0317_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_57_Left_155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_1_157 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_135 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1532_ _0528_ _0289_ _0147_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1463_ _0263_ _0107_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_91_Right_91 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1394_ cal_lut\[68\] _0805_ _0234_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA_input1_I io_in[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0868__A1 _0362_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_66_Left_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_89_296 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_224 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_268 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_279 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_322 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_75_Left_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1596__A2 _0780_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_314 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_325 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_185 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1348__A2 _0802_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1834__CLK net12 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_84_Left_182 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1520__A2 _0779_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_512 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_266 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_93_Left_191 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1587__A2 _0294_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_18 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_79_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1324__I _0779_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_87_681 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1707__CLK net11 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_200 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_548 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_119 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1857__CLK clknet_1_0__leaf_io_in[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xdec1._099_ dec1._031_ dec1._034_ dec1._028_ dec1._039_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XANTENNA__1578__A2 _0780_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_0963_ cal_lut\[176\] _0490_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_70_592 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_347 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1042__A4 _0384_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_185 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0894_ _0390_ _0363_ _0365_ _0356_ _0422_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_1515_ _0287_ _0135_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_57_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_288 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1446_ cal_lut\[97\] _0240_ _0257_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1377_ _0226_ _0058_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1502__A2 _0779_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_84 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1266__A1 ctr\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_50 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_417 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_277 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_303 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1569__A2 _0289_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_111 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1009__A1 _0376_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_325 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_185 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_13 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_199 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_28 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1300_ _0442_ _0790_ _0013_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__0940__B1 _0408_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_88 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1231_ temp1.dac.i_data\[3\] _0709_ _0684_ _0743_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1496__A1 cal_lut\[126\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1162_ ctr\[6\] _0672_ _0679_ temp1.dac.i_data\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XANTENNA__0893__I cal_lut\[37\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1093_ _0615_ _0395_ _0616_ _0617_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_59_200 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1248__A1 ctr\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_203 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_90_698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_314 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_111 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_100 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0946_ cal_lut\[80\] _0473_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_30_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_42_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0877_ _0365_ _0355_ _0405_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__0931__B1 _0379_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1429_ cal_lut\[89\] _0240_ _0248_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA_temp1.dcdc_EN temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_ VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1239__A1 ctr\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0922__B1 _0433_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_364 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_417 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_225 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1780_ _0132_ net8 cal_lut\[133\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_71_239 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_27 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_155 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_199 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_1_1__f_temp1.i_precharge_n clknet_0_temp1.i_precharge_n clknet_1_1__leaf_temp1.i_precharge_n
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_1214_ _0696_ _0701_ _0687_ _0727_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1145_ _0665_ _0666_ _0667_ _0668_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_94_309 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1076_ _0360_ _0413_ _0406_ _0600_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_62_41 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1641__A1 _0783_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0995__A3 _0422_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_291 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0929_ _0360_ cal_lut\[32\] _0373_ _0456_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_70_261 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_3_221 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_11_Left_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_26_345 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_372 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_20_Left_118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
Xtemp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref temp1.dac.parallel_cells\[3\].vdac_batch.en_vref
+ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__invz_3
Xtemp1.dac.parallel_cells\[1\].vdac_batch.einvp_batch\[0\].pupd temp1.dac.parallel_cells\[1\].vdac_batch.en_pupd
+ temp1.dac.parallel_cells\[1\].vdac_batch.npu_pd temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__invz_2
XFILLER_0_29_258 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1623__A1 ctr\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_239 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1832_ _0184_ net17 cal_lut\[185\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xtemp1.dac.parallel_cells\[0\].vdac_batch._6_ temp1.dac.parallel_cells\[0\].vdac_batch._2_
+ temp1.dac.parallel_cells\[0\].vdac_batch.en_pupd VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1763_ _0115_ net14 cal_lut\[116\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1694_ _0046_ net18 cal_lut\[47\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_57_85 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_202 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_48_470 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1128_ _0360_ cal_lut\[36\] _0373_ _0651_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1059_ _0368_ _0357_ _0584_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__1614__A1 ctr\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0968__A3 _0494_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_272 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1605__A1 _0365_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1740__CLK net15 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_375 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1081__A2 _0452_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_283 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_94_39 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0895__A2 _0365_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_37_407 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_451 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_228 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1072__A2 _0413_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_194 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_122 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_133 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1815_ _0167_ net13 cal_lut\[168\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1746_ _0098_ net12 cal_lut\[99\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_220 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1677_ _0029_ net11 cal_lut\[30\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_84_50 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_68_576 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1763__CLK net14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_342 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_51_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_261 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_197 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0877__A2 _0355_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_161 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_39 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1600_ net24 _0347_ _0677_ _0316_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1531_ _0484_ _0289_ _0146_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1462_ cal_lut\[107\] _0255_ _0263_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_38_32 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1393_ _0233_ _0067_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_38_87 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1786__CLK net12 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0868__A2 _0363_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_20 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_275 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1293__A2 _0790_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_258 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_286 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1729_ _0081_ net16 cal_lut\[82\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__0859__A2 _0383_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_513 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1284__A2 _0780_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_278 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_301 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_345 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_183 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1659__CLK net14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_79_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_87_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1027__A2 _0389_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_345 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0962_ _0487_ _0401_ _0440_ _0441_ _0488_ _0489_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai32_2
Xdec1._098_ dec1._028_ dec1._034_ dec1._036_ dec1._037_ dec1._038_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_6_239 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0893_ cal_lut\[37\] _0421_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1514_ cal_lut\[135\] _0779_ _0287_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_10_256 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1445_ _0256_ _0096_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1376_ cal_lut\[58\] _0802_ _0226_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_77_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1801__CLK net10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_315 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_123 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_dec1._078__A1 dec1.i_bin\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_407 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_164 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_292 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_10_47 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_18 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1193__A1 _0684_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1230_ _0362_ _0687_ _0704_ _0741_ _0742_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_1161_ _0345_ _0672_ _0679_ temp1.dac.i_data\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__1496__A2 _0240_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1092_ _0376_ cal_lut\[119\] _0413_ _0406_ _0616_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_35_44 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1824__CLK net2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_418 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_237 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_90_699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_259 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0945_ cal_lut\[158\] _0472_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_0876_ cal_lut\[43\] _0404_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1420__A2 _0790_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_297 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1245__I _0357_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_51 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1428_ _0564_ _0790_ _0088_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1359_ _0217_ _0049_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_65_204 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_410 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1411__A2 _0805_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1478__A2 _0255_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1847__CLK clknet_1_1__leaf_io_in[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_72_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_237 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_68 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_123 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1402__A2 _0802_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_384 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1065__I _0397_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_395 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__0913__A1 _0359_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1213_ _0688_ _0725_ _0726_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_95_725 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1469__A2 _0791_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1144_ cal_lut\[72\] _0383_ _0589_ cal_lut\[108\] _0667_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1075_ _0376_ _0369_ _0401_ _0599_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_1_67 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_345 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout15_I net2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_0928_ _0453_ _0454_ _0455_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_70_240 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_251 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0859_ cal_lut\[67\] _0383_ _0386_ cal_lut\[73\] _0387_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_11_340 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0904__A1 _0358_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_3_222 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_26_346 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_340 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_38_215 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_384 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1632__A2 _0351_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_259 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_390 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_24 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_181 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_29_248 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1831_ _0183_ net17 cal_lut\[184\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_84_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xtemp1.dac.parallel_cells\[0\].vdac_batch._5_ temp1.dac.i_enable temp1.dac.parallel_cells\[0\].vdac_batch._1_
+ temp1.dac.parallel_cells\[0\].vdac_batch._2_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_52_251 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1762_ _0114_ net14 cal_lut\[115\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1693_ _0045_ net17 cal_lut\[46\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_32_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_48_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1127_ cal_lut\[78\] _0386_ _0650_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_137 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1058_ _0543_ _0548_ _0582_ _0433_ cal_lut\[4\] _0583_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai32_4
XFILLER_0_90_357 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_7_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1090__A3 _0367_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xtemp1.dac.parallel_cells\[1\].vdac_batch.einvp_batch\[0\].vref temp1.dac.parallel_cells\[1\].vdac_batch.en_vref
+ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__invz_3
XFILLER_0_43_251 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1692__CLK net17 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_1_Right_1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_11_170 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_129 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_343 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_229 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_34_273 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xseg1._58_ seg1._22_ seg1._24_ seg1._25_ seg1.o_segments\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__0895__A3 _0356_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_37_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_452 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_66 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1814_ _0166_ net12 cal_lut\[167\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_72_357 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_4_167 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1518__I _0779_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1745_ _0097_ net12 cal_lut\[98\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1676_ _0028_ net11 cal_lut\[29\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__0886__A3 _0355_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_68_577 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_416 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref_I temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_321 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_354 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1063__A3 _0355_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_346 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_240 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_232 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_310 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1112__B _0357_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_332 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_42_433 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1054__A3 _0413_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_346 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_121 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_232 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1530_ _0435_ _0289_ _0145_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1461_ _0550_ _0791_ _0106_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1392_ cal_lut\[67\] _0805_ _0233_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_77_416 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_346 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_154 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_327 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1728_ _0080_ net16 cal_lut\[81\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1659_ _0011_ net14 cal_lut\[12\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_95_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1730__CLK net16 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xtemp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].pupd temp1.dac.parallel_cells\[3\].vdac_batch.en_pupd
+ temp1.dac.parallel_cells\[3\].vdac_batch.npu_pd temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__invz_2
XTAP_TAPCELL_ROW_56_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_224 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_313 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_173 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_121 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1107__B _0630_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_79_639 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_87_683 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_24 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_202 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_57 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_121 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0961_ cal_lut\[14\] _0488_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xdec1._097_ dec1._018_ dec1._019_ dec1._037_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_54_187 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0892_ _0360_ _0417_ _0378_ _0418_ _0419_ _0420_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai32_2
XANTENNA__1753__CLK net10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1513_ _0286_ _0134_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_50_393 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1444_ cal_lut\[96\] _0255_ _0256_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1375_ _0225_ _0057_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_65_31 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_52 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_63 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_279 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_154 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_327 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_102 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_84_664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_216 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1009__A3 _0413_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_154 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_290 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1776__CLK net8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_305 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_382 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0940__A2 _0407_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1160_ ctr\[4\] _0672_ _0679_ temp1.dac.i_data\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_1091_ cal_lut\[191\] _0615_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_15_285 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_66 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_290 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_165 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_113 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0944_ _0469_ _0414_ _0470_ _0471_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_0875_ _0362_ _0364_ _0384_ _0403_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_0_2_221 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__0931__A2 _0377_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1427_ _0520_ _0791_ _0087_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_97_308 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1649__CLK net8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1358_ cal_lut\[49\] _0805_ _0217_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1289_ _0789_ _0006_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1799__CLK net9 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_187 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_135 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_29_366 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_72_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1238__I0 _0675_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_293 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0913__A2 _0365_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1212_ _0343_ _0724_ _0690_ _0725_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_95_726 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1143_ _0368_ cal_lut\[132\] _0373_ _0666_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1074_ _0590_ _0591_ _0594_ _0597_ _0598_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_62_54 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_7_302 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0927_ _0368_ cal_lut\[134\] _0370_ _0454_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_0858_ _0384_ _0385_ _0386_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__1157__A2 _0678_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0904__A2 _0390_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_3_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xtemp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].pupd temp1.dac.parallel_cells\[4\].vdac_batch.en_pupd
+ temp1.dac.parallel_cells\[4\].vdac_batch.npu_pd temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__invz_2
XTAP_TAPCELL_ROW_26_347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_344 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_34_391 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1396__A2 _0805_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_127 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1814__CLK net12 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1148__A2 _0433_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1320__A2 _0783_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_171 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_205 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_216 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_84_300 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1830_ _0182_ net17 cal_lut\[183\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xtemp1.dac.parallel_cells\[0\].vdac_batch._4_ temp1.dac.i_data\[0\] temp1.dac.i_data\[5\]
+ temp1.dac.parallel_cells\[0\].vdac_batch._1_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__1387__A2 _0802_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1761_ _0113_ net15 cal_lut\[114\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1692_ _0044_ net17 cal_lut\[45\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_149 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_31 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_0_204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1126_ _0648_ _0649_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1311__A2 _0791_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1057_ _0552_ _0556_ _0569_ _0581_ _0582_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_75_311 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1075__A1 _0376_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_303 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_325 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1837__CLK net10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1378__A2 _0791_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_241 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_dec1._123__B2 dec1.i_tens VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1550__A2 _0289_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1302__A2 _0790_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1066__A1 cal_lut\[107\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_dec1._114__A1 dec1.i_tens VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xseg1._57_ seg1._11_ seg1._04_ seg1._06_ seg1._25_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_34_296 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_37_409 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_45 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_45_453 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1057__A1 _0552_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_208 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_303 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_314 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1813_ _0165_ net13 cal_lut\[166\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_4_124 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_241 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1744_ _0096_ net12 cal_lut\[97\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_7_67 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_78 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_255 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1675_ _0027_ net15 cal_lut\[28\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_68_31 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_15_Right_15 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1532__A2 _0289_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0886__A4 _0413_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_68_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_24_Right_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1109_ _0433_ _0632_ _0633_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_48_311 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1048__A1 _0358_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1599__A2 _0780_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1063__A4 _0413_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_31_222 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_33_Right_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[2\].vref_I temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1523__A2 _0791_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_42_Right_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_17_Left_115 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_42_434 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1054__A4 _0406_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_314 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_185 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_100 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_144 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_51_Right_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_22_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1460_ _0506_ _0791_ _0105_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_26_Left_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1391_ _0232_ _0066_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_38_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_45 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1514__A2 _0779_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_60_Right_60 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_54_33 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_255 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1682__CLK net11 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_35_Left_133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_89_277 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_288 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_238 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_21 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_314 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_166 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_44_Left_142 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1727_ _0079_ net16 cal_lut\[80\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1658_ _0010_ net15 cal_lut\[11\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1589_ cal_lut\[184\] _0294_ _0313_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__1269__A1 temp1.dac.i_enable VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_53_Left_151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_56_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_258 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_347 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_62_Left_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_5_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_87_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_417 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtemp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].vref temp1.dac.parallel_cells\[3\].vdac_batch.en_vref
+ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__invz_3
XFILLER_0_27_325 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_111 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0960_ cal_lut\[170\] _0487_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xdec1._096_ dec1._028_ dec1._035_ dec1._027_ dec1._036_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_27_347 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_57 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0891_ cal_lut\[79\] _0419_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xtemp1.inv2_3 clknet_1_0__leaf_net23 net24 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
X_1512_ cal_lut\[134\] _0255_ _0286_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_10_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_258 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1443_ _0782_ _0255_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_49_88 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1374_ cal_lut\[57\] _0805_ _0225_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_65_65 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_203 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_236 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_42 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_269 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1423__A1 cal_lut\[84\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_339 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_158 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_84_665 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_100 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_228 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1009__A4 _0406_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_57 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1090_ _0376_ _0612_ _0367_ _0445_ _0613_ _0614_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_0_27_111 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_15_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_144 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1720__CLK net11 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xdec1._079_ dec1._011_ dec1._010_ dec1._014_ dec1._019_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_27_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0943_ _0360_ cal_lut\[92\] _0394_ _0470_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_15_328 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0874_ _0359_ _0369_ _0401_ _0402_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_82_294 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_53 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1426_ _0476_ _0790_ _0086_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1357_ _0216_ _0048_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1288_ cal_lut\[6\] _0780_ _0789_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__1644__A1 _0783_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_temp1.dac.parallel_cells\[3\].vdac_batch._4__A1 temp1.dac.i_data\[3\] VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0922__A3 _0449_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1743__CLK net13 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_217 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtemp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[5\].pupd temp1.dac.parallel_cells\[4\].vdac_batch.en_pupd
+ temp1.dac.parallel_cells\[4\].vdac_batch.npu_pd temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__invz_2
XFILLER_0_64_261 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_19 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__0913__A3 _0356_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1211_ _0720_ _0722_ _0723_ _0724_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_46_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_95_727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1142_ cal_lut\[114\] _0596_ _0665_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_9_Left_107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_1_14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1073_ cal_lut\[95\] _0595_ _0596_ cal_lut\[113\] _0597_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_1_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_33 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_44 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1626__A1 _0783_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_88 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0926_ cal_lut\[152\] _0452_ _0453_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_55_272 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_220 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_1_0__f_io_in[0]_I clknet_0_io_in[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1537__I _0782_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_0857_ _0362_ _0363_ _0385_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_0_11_331 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0904__A3 _0363_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1409_ cal_lut\[75\] _0240_ _0242_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XPHY_EDGE_ROW_89_Right_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1766__CLK net12 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1617__A1 _0346_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_26_348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1093__A2 _0395_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_34_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_275 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_92_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1608__A1 ctr\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_331 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_312 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1760_ _0112_ net15 cal_lut\[113\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xtemp1.dac.parallel_cells\[0\].vdac_batch._3_ temp1.dac.i_data\[0\] temp1.dac.parallel_cells\[0\].vdac_batch.npu_pd
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xtemp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref temp1.dac.parallel_cells\[4\].vdac_batch.en_vref
+ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__invz_3
XFILLER_0_4_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_242 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_253 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1691_ _0043_ net17 cal_lut\[44\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_52_264 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1789__CLK net14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_21 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_0_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1125_ cal_lut\[150\] _0647_ _0379_ cal_lut\[66\] _0648_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_temp1.dac.parallel_cells\[0\].vdac_batch._7__I temp1.dac.i_enable VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1056_ _0571_ _0574_ _0577_ _0580_ _0581_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XTAP_TAPCELL_ROW_23_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_133 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_31_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0909_ _0376_ cal_lut\[97\] _0391_ _0413_ _0437_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__1216__B _0684_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_161 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_345 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_19_272 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_348 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_294 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_242 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xseg1._56_ dec1.o_dec\[1\] seg1._03_ seg1._00_ seg1._24_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_27_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_45_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_301 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_57 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1057__A2 _0556_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_131 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1812_ _0164_ net13 cal_lut\[165\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_25_275 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1743_ _0095_ net13 cal_lut\[96\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_4_169 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_223 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1674_ _0026_ net15 cal_lut\[27\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_342 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_40_289 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_68_579 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1296__A2 _0780_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1108_ cal_lut\[125\] _0392_ _0632_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_48_323 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_120 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1804__CLK net16 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1039_ cal_lut\[88\] _0564_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_75_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_16_242 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_297 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_42_435 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_381 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xseg1._39_ dec1.o_dec\[1\] dec1.o_dec\[0\] seg1._12_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__0970__A1 _0357_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1390_ cal_lut\[66\] _0802_ _0232_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_89_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_223 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1278__A2 _0783_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1827__CLK net2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_153 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_326 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1450__A2 _0255_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_99 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_189 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_0_io_in[0] io_in[0] clknet_0_io_in[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_85_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1726_ _0078_ net15 cal_lut\[79\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1657_ _0009_ net15 cal_lut\[10\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1588_ _0312_ _0183_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1269__A2 _0709_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_226 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_337 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1441__A2 _0240_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0952__A1 _0390_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_87_685 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_39_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_175 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xdec1._095_ dec1._015_ dec1._030_ dec1._034_ dec1._035_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_0890_ _0359_ _0366_ _0355_ _0385_ _0418_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_50_351 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtemp1.inv2_4 clknet_1_1__leaf_net23 net25 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
X_1511_ _0285_ _0133_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1442_ _0254_ _0095_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_49_67 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0943__A1 _0360_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1373_ _0224_ _0056_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_81_10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1120__A1 _0368_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_61_541 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1423__A2 _0805_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_307 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_253 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1187__A1 _0346_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1709_ _0061_ net8 cal_lut\[62\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_84_666 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_167 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_17 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_384 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1672__CLK net15 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_9_252 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0925__A1 _0360_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1102__A1 _0360_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_248 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_207 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_1_0__f_net23 clknet_0_net23 clknet_1_0__leaf_net23 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_15_287 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xdec1._078_ dec1.i_bin\[3\] dec1._017_ dec1._018_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_42_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0942_ cal_lut\[8\] _0469_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_0873_ _0362_ _0363_ _0401_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XPHY_EDGE_ROW_81_Left_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_76_43 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1425_ _0424_ _0791_ _0085_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1356_ cal_lut\[48\] _0802_ _0216_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1287_ _0788_ _0005_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_90_Left_188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__0852__B1 _0379_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_251 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_137 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1695__CLK net18 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_temp1.dac.parallel_cells\[3\].vdac_batch._4__A2 temp1.dac.i_data\[5\] VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_384 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1580__A1 _0613_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_603 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_12_268 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_170 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_376 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0913__A4 _0413_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1210_ ctr\[4\] _0694_ _0723_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_95_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1141_ _0368_ cal_lut\[120\] _0413_ _0406_ _0664_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_1072_ _0368_ _0413_ _0592_ _0596_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_1_48 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_59 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_56 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_337 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_402 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0925_ _0360_ _0367_ _0452_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_55_295 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_60 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xtemp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[5\].vref temp1.dac.parallel_cells\[4\].vdac_batch.en_vref
+ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__invz_3
XFILLER_0_30_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0856_ _0358_ _0365_ _0355_ _0384_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XANTENNA_temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[2\].vref_I temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_298 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_20 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0904__A4 _0406_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1408_ _0241_ _0074_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1339_ _0810_ _0035_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1617__A2 _0791_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_26_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_34_393 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_251 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_381 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1710__CLK net8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_92_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1860__CLK clknet_1_0__leaf_io_in[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_343 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_365 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_48 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_262 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1690_ _0042_ net17 cal_lut\[43\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_57_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_89 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_0_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1124_ _0381_ _0440_ _0647_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1055_ _0578_ _0445_ _0579_ _0580_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_73_66 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_99 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1075__A3 _0401_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_335 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0822__A3 _0351_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_240 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_70 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_fanout13_I net2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_31_374 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_416 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0908_ _0358_ _0362_ _0364_ _0391_ _0436_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_43_254 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_276 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_340 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0839_ _0362_ _0364_ _0366_ _0355_ _0367_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XANTENNA__1733__CLK net18 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_162 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_335 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_78_173 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_54_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_198 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_284 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_221 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xseg1._55_ seg1._00_ seg1._23_ seg1._10_ seg1.o_segments\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_89_416 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_36 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1057__A3 _0569_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_346 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1811_ _0163_ net13 cal_lut\[164\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_84_165 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_198 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_4_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_416 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_137 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_202 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1756__CLK net15 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1742_ _0094_ net15 cal_lut\[95\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_80_371 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1673_ _0025_ net15 cal_lut\[26\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_68_11 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_257 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_376 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_30_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_32 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_54 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_87 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_36_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_5_Right_5 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1107_ _0360_ _0629_ _0378_ _0630_ _0631_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_1038_ cal_lut\[40\] _0563_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1048__A3 _0391_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_346 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_265 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_279 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_302 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_42_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1779__CLK net8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_338 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_50_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_213 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xseg1._38_ seg1._00_ seg1._11_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_22_279 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_10_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_207 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_121 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_124 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1725_ _0077_ net15 cal_lut\[78\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_78_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_190 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1656_ _0008_ net16 cal_lut\[9\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1587_ cal_lut\[183\] _0294_ _0312_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_68_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_305 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0952__A2 _0363_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_205 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_238 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xdec1._094_ dec1._011_ dec1._021_ dec1._019_ dec1.i_bin\[2\] dec1._034_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_54_146 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_308 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_360 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1196__A2 _0709_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1510_ cal_lut\[133\] _0779_ _0285_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_49_24 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1441_ cal_lut\[95\] _0240_ _0254_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1372_ cal_lut\[56\] _0805_ _0224_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_4_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_631 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1120__A2 cal_lut\[102\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_55 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_146 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_382 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_298 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1708_ _0060_ net9 cal_lut\[61\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1639_ _0353_ _0337_ _0783_ _0209_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_69_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_227 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_84_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1817__CLK net14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__0925__A2 _0367_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_9_253 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1350__A2 _0790_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_59 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1102__A2 _0362_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0861__A1 _0359_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_124 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0941_ cal_lut\[182\] _0402_ _0403_ cal_lut\[50\] _0467_ _0468_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XTAP_TAPCELL_ROW_15_288 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xdec1._077_ dec1._010_ dec1._012_ dec1._014_ dec1._017_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_0872_ cal_lut\[163\] _0389_ _0392_ cal_lut\[121\] _0399_ _0400_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_23_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_33 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1424_ _0247_ _0084_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_76_88 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1355_ _0215_ _0047_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1286_ cal_lut\[5\] _0780_ _0788_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_81_648 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_157 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_263 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_296 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_41_160 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1580__A2 _0780_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1332__A2 _0805_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0843__A1 _0368_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_271 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_12_269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_274 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1020__A1 _0368_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_193 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1571__A2 _0289_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_95_729 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1140_ _0364_ cal_lut\[30\] _0384_ _0390_ _0663_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_1_16 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1071_ _0360_ _0394_ _0595_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__1087__A1 _0360_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_349 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0924_ _0357_ _0450_ _0451_ dec1.i_bin\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_0855_ _0358_ _0381_ _0382_ _0383_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_70_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1407_ cal_lut\[74\] _0240_ _0241_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__1314__A2 _0780_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1338_ cal_lut\[35\] _0802_ _0810_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_36_91 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1269_ temp1.dac.i_enable _0709_ _0776_ _0777_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1078__A1 _0368_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1662__CLK net17 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[15\].vref_I temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_34_394 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_263 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1553__A2 _0289_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_28 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1069__A1 _0360_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_314 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1241__A1 _0368_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_222 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_417 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1544__A2 _0294_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1685__CLK net16 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1123_ _0642_ _0643_ _0644_ _0645_ _0646_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__1603__B _0782_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1054_ _0358_ cal_lut\[118\] _0413_ _0406_ _0579_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_87_185 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_146 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_263 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_93 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_31_375 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0907_ cal_lut\[145\] _0435_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_3_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0838_ _0365_ _0366_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_4
XFILLER_0_11_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1535__A2 _0255_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_39_420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_314 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_325 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_241 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_263 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_380 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_277 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xseg1._54_ seg1._12_ seg1._22_ seg1._23_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__0982__B1 _0392_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1526__A2 _0255_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_59 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1462__A1 cal_lut\[107\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_133 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1810_ _0162_ net10 cal_lut\[163\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_72_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1741_ _0093_ net15 cal_lut\[94\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1672_ _0024_ net15 cal_lut\[25\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_80_383 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_23 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_45 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1106_ _0368_ cal_lut\[131\] _0373_ _0630_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
XTAP_TAPCELL_ROW_36_401 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1048__A4 _0413_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1037_ _0359_ _0560_ _0378_ _0418_ _0561_ _0562_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_0_90_103 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1205__A1 _0365_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_391 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1700__CLK net17 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_171 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1294__I _0782_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1508__A2 _0255_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1850__CLK clknet_1_1__leaf_io_in[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_11_Right_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_39_369 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_437 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xtemp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[2\].pupd temp1.dac.parallel_cells\[3\].vdac_batch.en_pupd
+ temp1.dac.parallel_cells\[3\].vdac_batch.npu_pd temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__invz_2
XTAP_TAPCELL_ROW_50_481 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_350 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_225 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_203 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xseg1._37_ seg1._00_ seg1._09_ seg1._10_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1_119 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_20_Right_20 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_38_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_89_214 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1723__CLK net11 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_103 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_380 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1724_ _0076_ net11 cal_lut\[77\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_85_8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1655_ _0007_ net16 cal_lut\[8\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_79_99 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1586_ _0311_ _0182_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_13_Left_111 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_95_76 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_22_Left_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_44_91 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1289__I _0789_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_263 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_158 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0937__B1 _0392_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1746__CLK net12 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_409 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_28 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_122 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xdec1._093_ dec1.i_bin\[1\] dec1._026_ dec1._032_ dec1._033_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XTAP_TAPCELL_ROW_70_587 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_169 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0831__I _0358_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1148__B _0357_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xtemp1.dac.parallel_cells\[3\].vdac_batch._8_ temp1.dac.parallel_cells\[3\].vdac_batch._0_
+ temp1.dac.parallel_cells\[3\].vdac_batch._1_ temp1.dac.parallel_cells\[3\].vdac_batch.en_vref
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA_temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[2\].vref_I temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1440_ _0253_ _0094_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__0943__A3 _0394_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1371_ _0223_ _0055_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_65_57 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1120__A3 _0391_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1611__B _0782_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_228 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_23 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_67 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_83 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_350 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_5_233 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_277 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1707_ _0059_ net11 cal_lut\[60\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1638_ _0343_ _0352_ _0337_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1569_ _0487_ _0289_ _0170_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1769__CLK net10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1647__A1 _0783_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_84_668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtemp1.dac.vdac_single._3__19 net19 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__tiel
Xfanout10 net13 net10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_83_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_286 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_128 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_9_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_59_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0940_ _0465_ _0407_ _0408_ _0466_ _0467_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai22_2
XTAP_TAPCELL_ROW_15_289 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xdec1._076_ dec1._007_ dec1._013_ dec1._015_ dec1._016_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_27_136 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0871_ _0393_ _0395_ _0397_ _0398_ _0399_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_0_2_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1423_ cal_lut\[84\] _0805_ _0247_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_48_8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1354_ cal_lut\[47\] _0802_ _0215_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1285_ _0787_ _0004_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1629__A1 _0783_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch._3__I temp1.dac.i_data\[4\] VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_77 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0852__A2 _0377_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_81_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_103 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_136 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_275 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_6_235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_264 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_286 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_191 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_297 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_356 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1070_ cal_lut\[71\] _0383_ _0593_ cal_lut\[17\] _0594_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__1087__A2 _0608_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_345 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0923_ _0365_ _0357_ _0451_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_0854_ _0365_ _0355_ _0382_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_23_150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_49_Right_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_11_356 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1406_ _0779_ _0240_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_1337_ _0809_ _0034_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_36_81 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1268_ _0687_ _0774_ _0775_ _0709_ _0776_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XPHY_EDGE_ROW_58_Right_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1199_ _0697_ _0712_ _0713_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1078__A2 _0365_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1807__CLK net16 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_348 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_242 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_201 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_245 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_67_Right_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_5_Left_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[5\].vref_I temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_76_Right_76 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_69_301 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1069__A2 _0413_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_25_340 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_39 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_220 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_404 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_37_264 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_85_Right_85 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_52_256 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_94_Right_94 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_57_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_13 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1122_ cal_lut\[90\] _0599_ _0600_ cal_lut\[24\] _0645_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XPHY_EDGE_ROW_69_Left_167 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1053_ cal_lut\[178\] _0578_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_87_120 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_87_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1480__A2 _0240_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_61 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_50 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_158 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_286 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_31_376 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_234 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0906_ _0431_ _0432_ _0433_ _0434_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_2
XPHY_EDGE_ROW_78_Left_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_0837_ dbg3\[1\] _0365_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_12
XFILLER_0_11_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_80 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_87_Left_185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_39_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_201 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_96_Left_194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
Xseg1._53_ dec1.o_dec\[2\] seg1._13_ seg1._22_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_43_16 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1462__A2 _0255_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_123 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_167 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_189 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_267 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1740_ _0092_ net15 cal_lut\[93\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1671_ _0023_ net15 cal_lut\[24\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1652__CLK net11 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1105_ cal_lut\[161\] _0629_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_36_402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1036_ cal_lut\[82\] _0561_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_33_82 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_16_267 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0964__A1 _0376_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_59_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1141__A1 _0368_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_67_571 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_326 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1444__A2 _0255_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_348 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_137 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_50_482 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1675__CLK net15 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xseg1._36_ seg1._08_ seg1._09_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_54_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1435__A2 _0240_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_318 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1723_ _0075_ net11 cal_lut\[76\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1609__B _0782_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtemp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[2\].vref temp1.dac.parallel_cells\[3\].vdac_batch.en_vref
+ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__invz_3
X_1654_ _0006_ net15 cal_lut\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1585_ cal_lut\[182\] _0294_ _0311_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xtemp1.dac.parallel_cells\[1\].vdac_batch.einvp_batch\[1\].pupd temp1.dac.parallel_cells\[1\].vdac_batch.en_pupd
+ temp1.dac.parallel_cells\[1\].vdac_batch.npu_pd temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__invz_2
XANTENNA__0882__B1 _0408_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1019_ _0360_ cal_lut\[34\] _0373_ _0544_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__1426__A2 _0790_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_137 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1698__CLK net17 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_297 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__0952__A4 _0384_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1254__B _0684_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1114__A1 _0635_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_292 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_262 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_251 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xdec1._092_ dec1._027_ dec1._028_ dec1._031_ dec1._032_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__1417__A2 _0790_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_70_588 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_39 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_321 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtemp1.dac.parallel_cells\[3\].vdac_batch._7_ temp1.dac.i_enable temp1.dac.parallel_cells\[3\].vdac_batch._0_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_49_26 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1370_ cal_lut\[55\] _0805_ _0223_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_4_39 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_78_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1120__A4 _0413_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_207 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1840__CLK clknet_1_1__leaf_io_in[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_51 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_273 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_201 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_384 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1706_ _0058_ net9 cal_lut\[59\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1637_ _0783_ _0336_ _0208_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1568_ _0439_ _0289_ _0169_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1499_ _0279_ _0127_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_84_669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout11 net13 net11 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_76_251 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_276 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_181 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_9_255 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1713__CLK net11 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_251 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_262 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xdec1._075_ dec1._011_ dec1._014_ dec1._015_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_0870_ cal_lut\[103\] _0398_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_42_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_287 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_181 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_41_Left_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_23_343 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_237 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtemp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[0\].pupd temp1.dac.parallel_cells\[4\].vdac_batch.en_pupd
+ temp1.dac.parallel_cells\[4\].vdac_batch.npu_pd temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__invz_2
X_1422_ _0246_ _0083_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1353_ _0553_ _0791_ _0046_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1284_ cal_lut\[4\] _0780_ _0787_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XPHY_EDGE_ROW_50_Left_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_92_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1622__B _0783_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_240 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_159 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_181 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0999_ _0515_ _0518_ _0521_ _0524_ _0525_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_74_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1736__CLK net18 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_6_236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_90 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0843__A3 _0370_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1020__A3 _0373_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1087__A3 _0422_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_28_360 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0922_ _0372_ _0388_ _0449_ _0433_ cal_lut\[1\] _0450_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai32_4
XANTENNA__1759__CLK net15 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_276 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0853_ _0362_ _0364_ _0381_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_70_224 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1405_ _0239_ _0073_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1336_ cal_lut\[34\] _0802_ _0809_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_94_720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput1 io_in[1] net1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1267_ ctr\[1\] _0687_ _0775_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1198_ seg1.o_segments\[1\] _0691_ _0712_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1078__A3 _0356_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_279 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1262__B _0684_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_335 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_25_341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_243 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_213 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_268 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1121_ cal_lut\[54\] _0403_ _0604_ cal_lut\[48\] _0644_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XTAP_TAPCELL_ROW_48_466 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1052_ _0575_ _0401_ _0440_ _0441_ _0576_ _0577_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_0_75_327 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_137 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_31_377 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0905_ _0384_ _0413_ _0433_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_43_268 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0836_ _0363_ _0364_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_8
XFILLER_0_37_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1319_ _0799_ _0026_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_78_165 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_93_135 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_276 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xseg1._52_ seg1._20_ seg1._21_ seg1.o_segments\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_34_268 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0982__A2 _0389_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_181 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_338 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_360 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_202 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1670_ _0022_ net16 cal_lut\[23\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_25_279 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_227 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_290 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_24 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1104_ _0623_ _0624_ _0627_ _0628_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
XTAP_TAPCELL_ROW_36_403 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1035_ cal_lut\[160\] _0560_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_48_338 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout11_I net13 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_371 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0819_ ctr\[4\] _0348_ _0349_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1799_ _0151_ net9 cal_lut\[152\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_3_195 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_59_528 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_572 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_90 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_360 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_227 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xseg1._35_ dec1.o_dec\[1\] dec1.o_dec\[2\] dec1.o_dec\[0\] seg1._08_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_15_290 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_271 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_28 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_16 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_135 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_382 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_416 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_190 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1722_ _0074_ net9 cal_lut\[75\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_53_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1653_ _0005_ net11 cal_lut\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_9_Right_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_21_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1584_ _0310_ _0181_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_95_67 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1018_ _0541_ _0542_ _0543_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_8_221 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_243 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_360 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_265 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_330 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__0937__A2 _0389_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1362__A2 _0805_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0873__A1 _0362_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_260 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_271 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xdec1._091_ dec1._015_ dec1._030_ dec1._031_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_35_330 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_70_589 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtemp1.dac.parallel_cells\[1\].vdac_batch.einvp_batch\[1\].vref temp1.dac.parallel_cells\[1\].vdac_batch.en_vref
+ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__invz_3
Xtemp1.dac.parallel_cells\[3\].vdac_batch._6_ temp1.dac.parallel_cells\[3\].vdac_batch._2_
+ temp1.dac.parallel_cells\[3\].vdac_batch.en_pupd VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_2_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_396 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1792__CLK net12 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_208 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1353__A2 _0791_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_78_634 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0864__A1 _0376_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_85 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1705_ _0057_ net8 cal_lut\[58\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_5_257 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_279 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_73 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_333 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0919__A2 _0445_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1636_ _0352_ _0335_ _0336_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_41_377 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[5\].vref_I temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_60 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1567_ _0306_ _0168_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1344__A2 _0790_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1498_ cal_lut\[127\] _0779_ _0279_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__0855__A1 _0358_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1665__CLK net14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout12 net13 net12 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_76_241 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_80 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_274 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_341 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1583__A2 _0294_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_9_256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1099__A1 _0368_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_75_615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0846__A1 _0360_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xdec1._074_ dec1.i_bin\[6\] dec1._005_ dec1._014_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__1271__A1 _0684_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_333 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_388 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1574__A2 _0294_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1421_ cal_lut\[83\] _0240_ _0246_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1352_ _0509_ _0790_ _0045_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1688__CLK net16 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1283_ _0786_ _0003_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_92_79 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_14_280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0998_ _0522_ _0427_ _0523_ _0524_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_73_288 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1014__A1 _0362_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1565__A2 _0289_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1619_ _0696_ _0347_ _0326_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_1_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xtemp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[0\].vref temp1.dac.parallel_cells\[4\].vdac_batch.en_vref
+ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__invz_3
XFILLER_0_5_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_6_237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_97_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_255 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1830__CLK net17 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1308__A2 _0790_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_39 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0819__A1 ctr\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_28_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0921_ _0400_ _0411_ _0430_ _0448_ _0449_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_0852_ cal_lut\[55\] _0377_ _0379_ cal_lut\[61\] _0380_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_55_299 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1404_ cal_lut\[73\] _0802_ _0239_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1335_ _0808_ _0033_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput2 io_in[2] net2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_94_721 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_61 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1266_ ctr\[7\] _0701_ _0773_ _0774_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1197_ _0357_ _0450_ _0691_ _0451_ _0711_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__1078__A4 _0401_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_325 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_336 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_328 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_403 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1703__CLK net8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_222 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_93 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_417 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_255 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1594__I _0315_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1538__A2 _0294_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1853__CLK clknet_1_1__leaf_io_in[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_347 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_358 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_369 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_96_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_342 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_37_255 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0985__B1 _0408_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_409 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0848__I _0358_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1120_ _0368_ cal_lut\[102\] _0391_ _0413_ _0643_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_73_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_48_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1051_ cal_lut\[16\] _0576_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1726__CLK net15 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_380 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_339 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_52 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_30 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xdec1._109_ dec1._018_ dec1._019_ dec1._048_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_28_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_266 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1217__A1 _0678_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_0904_ _0358_ _0390_ _0363_ _0406_ _0432_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XANTENNA__0976__B1 _0379_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_258 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0835_ dbg3\[2\] _0363_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_12
XFILLER_0_11_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1318_ cal_lut\[26\] _0783_ _0799_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1249_ dec1.i_tens _0682_ _0686_ _0681_ _0759_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__1456__A1 cal_lut\[102\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_78_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_22_323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_255 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_225 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_372 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xseg1._51_ dec1.o_dec\[1\] seg1._03_ seg1._11_ seg1._01_ seg1._21_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_6_160 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_171 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_291 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1749__CLK net10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_103 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_15 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_58 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_63 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1103_ cal_lut\[173\] _0625_ _0626_ cal_lut\[143\] _0627_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XTAP_TAPCELL_ROW_36_404 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1034_ _0557_ _0414_ _0558_ _0559_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_48_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_62 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_158 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_169 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_383 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_236 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1610__A1 _0345_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1798_ _0150_ net9 cal_lut\[151\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_31_239 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_228 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0818_ ctr\[2\] ctr\[3\] _0347_ _0348_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__0964__A3 _0413_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_59_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1141__A3 _0413_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_67_573 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1429__A1 cal_lut\[89\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_103 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_372 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_342 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_217 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xseg1._34_ seg1._00_ seg1._02_ seg1._04_ seg1._07_ seg1.o_segments\[0\] VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
Xtemp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[13\].pupd temp1.dac.parallel_cells\[4\].vdac_batch.en_pupd
+ temp1.dac.parallel_cells\[4\].vdac_batch.npu_pd temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__invz_2
XANTENNA_temp1.dac.parallel_cells\[0\].vdac_batch._5__A1 temp1.dac.i_enable VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_27 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1721_ _0073_ net9 cal_lut\[74\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1652_ _0004_ net11 cal_lut\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_79_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_194 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1583_ cal_lut\[181\] _0294_ _0310_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__0882__A2 _0407_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1017_ _0368_ cal_lut\[136\] _0370_ _0542_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_64_554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_309 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_169 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_82 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_283 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0873__A2 _0363_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_253 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xdec1._090_ dec1.i_bin\[3\] dec1._017_ dec1._029_ dec1._030_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_39_136 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_128 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_364 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtemp1.dac.parallel_cells\[3\].vdac_batch._5_ temp1.dac.i_enable temp1.dac.parallel_cells\[3\].vdac_batch._1_
+ temp1.dac.parallel_cells\[3\].vdac_batch._2_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_35_386 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_17 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_78_635 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0864__A2 _0390_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_15 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_26 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_81_59 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_220 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1704_ _0056_ net8 cal_lut\[57\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_5_269 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1635_ _0674_ _0334_ _0335_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_69_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1566_ cal_lut\[168\] _0294_ _0306_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1497_ _0278_ _0126_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_12_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xfanout13 net2 net13 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_91_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_286 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1280__A2 _0783_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_75_616 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0846__A2 cal_lut\[31\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_83_660 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xdec1._073_ dec1._010_ dec1._012_ dec1._013_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_55_404 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_67_286 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_128 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_323 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_183 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_356 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1023__A2 _0545_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_164 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1420_ _0561_ _0790_ _0082_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1351_ _0465_ _0790_ _0044_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1282_ cal_lut\[3\] _0783_ _0786_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_92_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_242 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1262__A2 _0709_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_418 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_267 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_312 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0997_ _0390_ _0363_ cal_lut\[27\] _0384_ _0523_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__1014__A2 _0357_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1618_ _0347_ _0673_ _0783_ _0200_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_6_238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1549_ _0300_ _0156_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_97_741 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_70 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_dec1._074__A1 dec1.i_bin\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1782__CLK net10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_404 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_64_278 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_289 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_337 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1492__A2 _0240_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_0920_ _0434_ _0438_ _0443_ _0447_ _0448_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_55_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_223 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_418 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_21 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0851_ _0376_ _0378_ _0379_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_23_131 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_259 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1655__CLK net16 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_348 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_18_Right_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1403_ _0238_ _0072_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1334_ cal_lut\[33\] _0805_ _0808_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_3_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1265_ _0681_ _0682_ _0691_ dec1.i_tens _0772_ _0773_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XTAP_TAPCELL_ROW_94_722 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput3 io_in[3] net3 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_36_73 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1196_ temp1.dac.i_data\[1\] _0709_ _0684_ _0710_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_27_Right_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_52_50 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_36_Right_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_10_381 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_45_Right_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1474__A2 _0240_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_25_343 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1678__CLK net11 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_226 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_54_Right_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_29_Left_127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_73_27 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_91_703 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_48_468 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_63_Right_63 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1050_ cal_lut\[172\] _0575_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_28_201 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_38_Left_136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_7_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xdec1._108_ dec1.i_bin\[1\] dec1._047_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XANTENNA__1217__A2 _0684_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_340 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_204 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0903_ cal_lut\[139\] _0431_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_22_86 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0834_ dbg3\[3\] _0362_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_12
XPHY_EDGE_ROW_72_Right_72 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_47_Left_145 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_51_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0900__A1 _0390_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1317_ _0798_ _0025_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_81_Right_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1248_ ctr\[7\] _0697_ _0690_ _0758_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_78_101 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1456__A2 _0255_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_56_Left_154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1179_ _0681_ _0693_ _0694_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_66_307 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_329 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_324 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1820__CLK net14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_384 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_362 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_90_Right_90 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
Xseg1._50_ seg1._00_ seg1._19_ seg1._20_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__0967__A1 _0464_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_65_Left_163 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_97_410 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_74_Left_172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_92_181 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0958__A1 _0376_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_218 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_83_Left_181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_80_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_68_27 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_92_Left_190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch._4__A1 temp1.dac.i_data\[4\] VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1102_ _0360_ _0362_ _0364_ _0382_ _0626_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XTAP_TAPCELL_ROW_36_405 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1843__CLK clknet_1_0__leaf_io_in[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1033_ _0359_ cal_lut\[94\] _0394_ _0558_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
Xtemp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[6\].pupd temp1.dac.parallel_cells\[4\].vdac_batch.en_pupd
+ temp1.dac.parallel_cells\[4\].vdac_batch.npu_pd temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__invz_2
XFILLER_0_75_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1639__B _0783_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1797_ _0149_ net12 cal_lut\[150\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_31_218 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0817_ _0346_ ctr\[1\] _0347_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__0964__A4 _0406_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1141__A4 _0406_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_67_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1429__A2 _0240_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_0_Right_0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_90_91 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_321 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1268__C _0709_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_354 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_365 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xseg1._33_ seg1._05_ seg1._06_ seg1._00_ seg1._07_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_62_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1716__CLK net8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_251 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_284 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1117__A1 cal_lut\[84\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_240 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_41_430 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1720_ _0072_ net11 cal_lut\[73\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_80_151 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1651_ _0003_ net11 cal_lut\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_79_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1582_ _0309_ _0180_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1356__A1 cal_lut\[48\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input6_I io_in[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_96 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1123__A4 _0645_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1016_ cal_lut\[154\] _0452_ _0541_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_64_555 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_273 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_295 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_416 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtemp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[13\].vref temp1.dac.parallel_cells\[4\].vdac_batch.en_vref
+ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__invz_3
XFILLER_0_56_181 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1739__CLK net16 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1849_ _0201_ clknet_1_1__leaf_io_in[0] ctr\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_5_9 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_243 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_310 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_170 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtemp1.dac.parallel_cells\[3\].vdac_batch._4_ temp1.dac.i_data\[3\] temp1.dac.i_data\[5\]
+ temp1.dac.parallel_cells\[3\].vdac_batch._1_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_62_173 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0864__A3 _0363_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_86_680 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_416 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_265 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1026__B1 _0397_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_237 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1703_ _0055_ net8 cal_lut\[56\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_26_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_30_53 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_97 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1634_ ctr\[8\] _0351_ _0334_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_41_368 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1565_ _0610_ _0289_ _0167_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_39_40 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1496_ cal_lut\[126\] _0240_ _0278_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_55_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_49_413 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout14 net2 net14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_17_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_32_368 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[8\].vref_I temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1099__A3 _0378_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_75_617 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0846__A3 _0373_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0906__B _0433_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_221 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_83_661 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xdec1._072_ dec1.i_bin\[6\] dec1._008_ dec1._011_ dec1._012_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_70_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_279 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_290 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_10_Left_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1350_ _0404_ _0790_ _0043_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1281_ _0785_ _0002_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_92_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_25_86 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_202 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0996_ cal_lut\[111\] _0522_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_73_279 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_346 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_176 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1617_ _0346_ _0791_ _0199_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_6_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1548_ cal_lut\[156\] _0294_ _0300_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_97_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_74 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1479_ _0269_ _0117_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_82_81 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_80_642 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_268 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_154 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_62_18 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_29 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_349 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_416 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_33 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0850_ _0362_ _0364_ _0365_ _0356_ _0378_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XTAP_TAPCELL_ROW_11_263 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_44 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_23_154 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1402_ cal_lut\[72\] _0802_ _0238_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1333_ _0807_ _0032_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1264_ _0357_ _0691_ _0772_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_94_723 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput4 io_in[4] net4 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_36_52 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1195_ _0681_ _0703_ _0709_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_0_34_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_205 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0979_ cal_lut\[189\] _0505_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_6_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_96_102 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_349 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_308 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_25_344 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_224 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_192 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_205 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__0985__A2 _0407_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_238 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_102 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_271 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_18 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_39 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_91_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_48_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_224 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xdec1._107_ dec1._045_ dec1._044_ dec1._043_ dec1._046_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_7_129 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_16_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0902_ _0416_ _0420_ _0425_ _0429_ _0430_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_0833_ cal_lut\[151\] _0361_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__0976__A2 _0377_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_249 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_238 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1772__CLK net10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_146 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1316_ cal_lut\[25\] _0783_ _0798_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_47_84 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0900__A2 _0363_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_31 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1247_ _0754_ _0691_ _0756_ _0694_ _0757_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1178_ _0686_ net5 _0693_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_78_124 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_61 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_127 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_22_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_257 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_341 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_205 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_216 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_140 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_238 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0967__A2 _0468_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_411 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_293 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1392__A2 _0805_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1144__A2 _0383_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_179 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_190 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_53_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1795__CLK net13 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1080__A1 _0376_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_355 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_33_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1383__A2 _0805_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch._4__A2 temp1.dac.i_data\[5\] VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1101_ _0376_ _0391_ _0385_ _0625_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__0894__A1 _0390_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1032_ cal_lut\[10\] _0557_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_33_64 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1071__A1 _0360_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_344 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1796_ _0148_ net12 cal_lut\[149\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0816_ ctr\[0\] _0346_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_3_187 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1374__A2 _0805_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_0_net23 net23 clknet_0_net23 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__1668__CLK net17 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_67_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_127 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtemp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[6\].vref temp1.dac.parallel_cells\[4\].vdac_batch.en_vref
+ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__invz_3
XANTENNA__1062__A1 _0368_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xseg1._32_ dec1.o_dec\[1\] seg1._01_ dec1.o_dec\[2\] seg1._06_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_30_241 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_1_1__f_io_in[0] clknet_0_io_in[0] clknet_1_1__leaf_io_in[0] VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_89_219 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_274 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_57_127 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_330 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_149 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_41_431 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_193 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1650_ _0002_ net11 cal_lut\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1581_ cal_lut\[180\] _0294_ _0309_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_21_241 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1356__A2 _0802_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1810__CLK net10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1108__A2 _0392_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_dec1._101__A1 dec1.i_tens VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0867__A1 _0358_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_41 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1015_ _0357_ _0539_ _0540_ dec1.i_bin\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_TAPCELL_ROW_64_556 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_235 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1595__A2 _0780_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1848_ _0200_ clknet_1_1__leaf_io_in[0] ctr\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_1779_ _0131_ net8 cal_lut\[132\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_296 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_285 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0858__A1 _0384_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_92 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_200 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_119 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_182 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtemp1.dac.parallel_cells\[3\].vdac_batch._3_ temp1.dac.i_data\[3\] temp1.dac.parallel_cells\[3\].vdac_batch.npu_pd
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_62_185 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1338__A2 _0802_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1833__CLK net2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0849__A1 _0376_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1510__A2 _0779_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0864__A4 _0391_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_277 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_288 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_5_216 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1702_ _0054_ net8 cal_lut\[55\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_65 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_325 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1577__A2 _0780_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1633_ _0783_ _0333_ _0207_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1564_ _0305_ _0166_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1495_ _0277_ _0125_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_39_63 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1706__CLK net9 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1265__B2 dec1.i_tens VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout15 net2 net15 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_64_417 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_119 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1017__A1 _0368_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1856__CLK clknet_1_0__leaf_io_in[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1568__A2 _0289_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_75_618 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1256__A1 _0670_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_233 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_83_662 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xdec1._071_ dec1.i_bin\[3\] dec1._011_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_3
XFILLER_0_67_255 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_23_303 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1559__A2 _0294_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_347 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1280_ cal_lut\[2\] _0783_ _0785_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__1729__CLK net16 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_65 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_299 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_64 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_314 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_14_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0995_ _0376_ _0519_ _0422_ _0423_ _0520_ _0521_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_0_81_291 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1616_ _0783_ clknet_1_1__leaf__0316_ _0325_ _0198_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_5_53 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1547_ _0299_ _0155_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_97_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1478_ cal_lut\[117\] _0255_ _0269_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_66_94 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_80_643 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_152 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_122 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_72_291 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_temp1.dac.parallel_cells\[3\].vdac_batch._3__I temp1.dac.i_data\[3\] VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xdec1._123_ dec1._003_ dec1._056_ dec1._059_ dec1.i_tens dec1.o_dec\[3\] VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_TAPCELL_ROW_11_264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_188 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1401_ _0237_ _0071_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1332_ cal_lut\[32\] _0805_ _0807_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1263_ temp1.dac.i_enable _0684_ _0770_ _0771_ io_out[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_TAPCELL_ROW_94_724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput5 io_in[5] net5 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_1194_ _0678_ _0684_ _0708_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_34_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1640__A1 _0733_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_269 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0978_ _0500_ _0501_ _0502_ _0503_ _0504_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_14_133 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_171 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1631__A1 _0783_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_217 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_91_705 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_136 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_372 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_33 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xdec1._106_ dec1._042_ dec1._043_ dec1._044_ dec1._045_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_28_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0901_ _0426_ _0427_ _0428_ _0429_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_0832_ _0359_ _0360_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__1138__B1 _0392_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1315_ _0797_ _0024_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1246_ dbg3\[5\] _0755_ _0635_ _0637_ _0691_ _0756_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_1177_ _0356_ _0357_ _0691_ _0692_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_19_203 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_22_326 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_152 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_228 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0967__A3 _0481_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_30_370 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_1_0__f_io_in[0] clknet_0_io_in[0] clknet_1_0__leaf_io_in[0] VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_42_283 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1129__B1 _0377_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_53_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_364 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0958__A3 _0391_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1080__A2 _0362_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_294 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1100_ _0360_ cal_lut\[35\] _0373_ _0624_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_17_55 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__0894__A2 _0363_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1031_ cal_lut\[184\] _0402_ _0403_ cal_lut\[52\] _0555_ _0556_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_56_331 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_375 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_228 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1071__A2 _0394_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1001__B _0433_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_312 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1795_ _0147_ net13 cal_lut\[148\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0815_ ctr\[5\] _0345_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_58_95 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1229_ _0688_ _0739_ _0740_ _0687_ _0741_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_47_364 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1062__A2 _0422_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_323 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xseg1._31_ dec1.o_dec\[1\] seg1._01_ seg1._05_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_62_356 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_294 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_30_275 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_58_521 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1762__CLK net14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_41_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_356 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1580_ _0613_ _0780_ _0179_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_21_286 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__0867__A2 _0394_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_31 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1014_ _0362_ _0357_ _0540_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_64_557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_253 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_88_275 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1292__A2 _0790_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_60_74 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_389 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1847_ _0199_ clknet_1_1__leaf_io_in[0] ctr\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1778_ _0130_ net8 cal_lut\[131\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_69_61 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1785__CLK net12 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_242 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_275 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_128 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_345 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_334 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0849__A2 _0367_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1274__A2 _0780_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_312 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1026__A2 _0395_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1658__CLK net15 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1701_ _0053_ net14 cal_lut\[54\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1632_ _0689_ _0351_ _0333_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1563_ cal_lut\[166\] _0294_ _0305_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1494_ cal_lut\[125\] _0255_ _0277_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_55_96 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_40 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout16 net18 net16 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_29_161 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_197 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_381 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_75_619 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_83_663 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xdec1._070_ dec1.i_bin\[6\] dec1._008_ dec1._009_ dec1._010_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_67_278 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1800__CLK net10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_164 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_186 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_90_292 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtemp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[3\].pupd temp1.dac.parallel_cells\[3\].vdac_batch.en_pupd
+ temp1.dac.parallel_cells\[3\].vdac_batch.npu_pd temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__invz_2
XFILLER_0_26_131 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_14_284 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_304 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_76 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0994_ cal_lut\[87\] _0520_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_41_156 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_dec1._087__I dec1.i_bin\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_220 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_178 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1615_ temp_delay_last _0685_ _0325_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_22_381 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_264 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1546_ cal_lut\[155\] _0294_ _0299_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_5_32 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_97_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0930__A1 _0368_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1477_ _0268_ _0116_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1486__A2 _0240_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_307 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1823__CLK net14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_80_644 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0997__A1 _0390_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_259 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_5_230 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0921__A1 _0400_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xdec1._122_ dec1.i_ones dec1._057_ dec1._058_ dec1._059_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__0988__A1 _0359_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_11_265 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_156 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_68 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1400_ cal_lut\[71\] _0802_ _0237_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__1165__A1 clknet_1_1__leaf_io_in[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1331_ _0806_ _0031_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__0912__A1 _0358_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1262_ clknet_1_0__leaf_temp1.i_precharge_n _0709_ _0684_ _0771_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xinput6 io_in[6] net6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__1846__CLK clknet_1_0__leaf_io_in[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1468__A2 _0791_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_19_310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1193_ _0684_ _0685_ _0707_ io_out[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_78_329 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_226 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_259 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_97 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0977_ cal_lut\[69\] _0383_ _0386_ cal_lut\[75\] _0503_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_58_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1529_ _0292_ _0144_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1459__A2 _0791_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_340 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_92_321 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_14_Right_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_37_259 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_45_270 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1719__CLK net11 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_251 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_273 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[11\].vref_I temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_23_Right_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_91_706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_32_Right_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_68_384 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xdec1._105_ dec1._003_ dec1._044_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_0900_ _0390_ _0363_ cal_lut\[25\] _0384_ _0428_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_43_218 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0831_ _0358_ _0359_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_12
XFILLER_0_3_348 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_41_Right_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1138__B2 cal_lut\[126\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_16_Left_114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1314_ cal_lut\[24\] _0780_ _0797_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__0897__B1 _0423_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1245_ _0357_ _0755_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__0900__A4 _0384_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1176_ _0681_ net6 net5 _0691_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XPHY_EDGE_ROW_50_Right_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_59_373 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_25_Left_123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_6_120 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_218 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_6_164 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_30_371 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_34_Left_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_84_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_43_Left_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_53_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_270 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__0958__A4 _0413_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1368__A1 cal_lut\[54\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_273 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_379 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1691__CLK net17 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_19 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_52_Left_150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_17_23 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__0894__A3 _0365_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_67 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1030_ _0553_ _0407_ _0408_ _0554_ _0555_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_0_56_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0814_ ctr\[7\] _0344_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_24_240 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1794_ _0146_ net13 cal_lut\[147\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_58_30 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1228_ ctr\[3\] _0688_ _0740_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1159_ ctr\[3\] _0672_ _0679_ temp1.dac.i_data\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_66_129 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_313 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_173 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xseg1._30_ dec1.o_dec\[0\] seg1._03_ seg1._04_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_50_477 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_58_522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_416 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_321 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_376 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1013_ _0499_ _0504_ _0538_ _0433_ cal_lut\[3\] _0539_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai32_4
XFILLER_0_48_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_64_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_310 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_321 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_44_313 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_346 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_32 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1846_ _0198_ clknet_1_0__leaf_io_in[0] temp_delay_last VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1777_ _0129_ net8 cal_lut\[130\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_243 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_4_Right_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_12_298 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_85_94 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_254 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_118 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_298 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_302 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_368 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtemp1.dac.parallel_cells\[1\].vdac_batch._8_ temp1.dac.parallel_cells\[1\].vdac_batch._0_
+ temp1.dac.parallel_cells\[1\].vdac_batch._1_ temp1.dac.parallel_cells\[1\].vdac_batch.en_vref
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_85_202 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_24 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_539 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_279 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1700_ _0052_ net17 cal_lut\[53\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_41_349 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1631_ _0783_ _0332_ _0206_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1562_ _0304_ _0165_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1493_ _0276_ _0124_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input4_I io_in[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_405 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout17 net18 net17 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_91_205 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout9_I net13 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1017__A3 _0370_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1829_ _0181_ net17 cal_lut\[182\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1752__CLK net10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_8_Left_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_40_393 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_79_Right_79 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_88_Right_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_23_349 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_168 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_8_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_97_Right_97 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_25_78 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_216 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0993_ cal_lut\[39\] _0519_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1775__CLK net8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1614_ ctr\[7\] clknet_1_0__leaf__0318_ _0324_ _0197_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1545_ _0298_ _0154_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1476_ cal_lut\[116\] _0240_ _0268_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_97_745 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_74 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_80_645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0997__A2 _0363_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_102 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtemp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[3\].vref temp1.dac.parallel_cells\[3\].vdac_batch.en_vref
+ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__invz_3
XFILLER_0_32_146 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0921__A2 _0411_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1648__CLK net8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xdec1._121_ dec1._047_ dec1._039_ dec1._050_ dec1._058_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__1798__CLK net9 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_25 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_260 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_135 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_11_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_18 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1330_ cal_lut\[31\] _0805_ _0806_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__0912__A2 _0391_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1261_ _0346_ _0687_ _0768_ _0769_ _0704_ _0770_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_36_33 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput7 io_in[7] net7 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1192_ _0705_ _0706_ _0684_ _0707_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_19_311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_77 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_238 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_313 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_290 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0976_ cal_lut\[57\] _0377_ _0379_ cal_lut\[63\] _0502_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_1528_ cal_lut\[144\] _0255_ _0292_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_77_95 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1459_ _0462_ _0791_ _0104_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_77_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_92_311 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1092__A1 _0376_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_227 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_52_219 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_263 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_190 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1156__I _0677_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_91_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xdec1._104_ dec1._016_ dec1._025_ dec1._043_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_28_216 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[1\].vref_I temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_208 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0830_ dbg3\[4\] _0358_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_12
XFILLER_0_51_241 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1813__CLK net13 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1313_ _0796_ _0023_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__0897__A1 _0376_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1244_ seg1.o_segments\[5\] _0754_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_47_76 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_39_417 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_45 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_56 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1175_ _0681_ _0686_ net5 _0690_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XANTENNA__1310__A2 _0790_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_47_461 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_341 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_160 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_333 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_22_328 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_208 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_372 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtemp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[1\].pupd temp1.dac.parallel_cells\[4\].vdac_batch.en_pupd
+ temp1.dac.parallel_cells\[4\].vdac_batch.npu_pd temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__invz_2
X_0959_ _0484_ _0436_ _0485_ _0486_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_70_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_382 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_193 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1301__A2 _0790_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_333 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_182 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_53_497 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_325 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1368__A2 _0802_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1836__CLK net10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_308 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__0879__A1 _0359_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1540__A2 _0294_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0894__A4 _0356_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_208 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_185 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0813_ ctr\[10\] _0343_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_71_336 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1793_ _0145_ net13 cal_lut\[146\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_58_64 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1531__A2 _0289_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1227_ _0733_ _0738_ _0690_ _0739_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__1709__CLK net8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1158_ ctr\[2\] _0672_ _0679_ temp1.dac.i_data\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_1089_ cal_lut\[179\] _0613_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_47_333 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_95 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1598__A2 _0780_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1859__CLK clknet_1_0__leaf_io_in[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_50_478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_185 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_255 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_288 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1522__A2 _0289_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_58_523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1589__A2 _0294_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_358 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1210__A1 ctr\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_89_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1012_ _0508_ _0512_ _0525_ _0537_ _0538_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_44_55 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_64_559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_99 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_32 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_325 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_185 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_98 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1845_ _0197_ clknet_1_0__leaf_io_in[0] dbg3\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_8_55 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1776_ _0128_ net8 cal_lut\[129\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_52_380 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_99 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_288 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1504__A2 _0255_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_71_Left_169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_67_417 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1681__CLK net8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_277 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_130 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_314 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_100 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_325 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_80_Left_178 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_7_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xtemp1.dac.parallel_cells\[1\].vdac_batch._7_ temp1.dac.i_enable temp1.dac.parallel_cells\[1\].vdac_batch._0_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_14_47 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_314 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_303 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_291 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_0_temp1.i_precharge_n temp1.i_precharge_n clknet_0_temp1.i_precharge_n VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_1630_ ctr\[7\] _0350_ _0332_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1561_ cal_lut\[165\] _0294_ _0304_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1492_ cal_lut\[124\] _0240_ _0276_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_39_88 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_417 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_225 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_64_409 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout18 net2 net18 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_76_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_258 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_44_111 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_241 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1828_ _0180_ net17 cal_lut\[181\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_20_90 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_296 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1759_ _0111_ net15 cal_lut\[112\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_96_94 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_8_251 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_13 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_74_610 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0992_ _0360_ _0516_ _0378_ _0418_ _0517_ _0518_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_0_26_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_361 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1613_ dbg3\[5\] clknet_1_0__leaf__0318_ _0782_ _0324_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1544_ cal_lut\[154\] _0294_ _0298_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_5_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0930__A3 _0373_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1475_ _0267_ _0115_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_66_42 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_97_746 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_41 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_269 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_100 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_155 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_261 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_199 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0921__A3 _0430_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_356 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xdec1._120_ dec1._039_ dec1._033_ dec1._050_ dec1._057_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_55_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0988__A3 _0394_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_267 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1260_ _0744_ _0701_ _0687_ _0769_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_1191_ temp1.dac.i_data\[0\] _0704_ _0706_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_36_89 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1625__A1 _0345_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1742__CLK net15 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_228 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0975_ _0368_ cal_lut\[129\] _0373_ _0501_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_77_63 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1527_ _0291_ _0143_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1458_ _0398_ _0791_ _0103_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_2_213 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1389_ _0622_ _0791_ _0065_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_93_95 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_dec1._063__B dec1.i_bin\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_301 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1616__A1 _0783_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_130 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_412 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_242 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1765__CLK net12 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xdec1._103_ dec1._004_ dec1._020_ dec1._042_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1607__A1 _0363_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_228 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1312_ cal_lut\[23\] _0780_ _0796_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_47_88 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1243_ _0752_ _0753_ _0731_ io_out[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_39_418 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1174_ ctr\[8\] _0689_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_63_10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_47_462 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_65 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_345 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout18_I net2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0958_ _0376_ cal_lut\[98\] _0391_ _0413_ _0485_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_42_220 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_231 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0889_ cal_lut\[157\] _0417_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_63_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1788__CLK net14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_161 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_53_498 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_345 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_356 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_194 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_294 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_286 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtemp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[1\].vref temp1.dac.parallel_cells\[4\].vdac_batch.en_vref
+ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__invz_3
XANTENNA__0879__A2 _0390_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_312 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_323 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_183 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtemp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[0\].pupd temp1.dac.parallel_cells\[2\].vdac_batch.en_pupd
+ temp1.dac.parallel_cells\[2\].vdac_batch.npu_pd temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__invz_2
XFILLER_0_83_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_367 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_153 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_0812_ dec1.i_ones dec1.i_tens VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XFILLER_0_71_348 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_103 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_231 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1792_ _0144_ net12 cal_lut\[145\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_24_297 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1226_ _0734_ _0736_ _0737_ _0738_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_74_53 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1157_ _0673_ _0678_ _0679_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__1220__1_I clknet_1_1__leaf_io_in[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1295__A2 _0791_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1088_ cal_lut\[59\] _0612_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_90_63 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_356 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_378 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_74_153 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_220 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_50_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_326 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_74_197 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_359 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_275 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_58_524 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1286__A2 _0780_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1803__CLK net12 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_323 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_80_156 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_89_693 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1011_ _0527_ _0530_ _0533_ _0536_ _0537_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_29_345 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_367 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_348 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_197 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_134 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1844_ _0196_ clknet_1_1__leaf_io_in[0] dbg3\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_201 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1775_ _0127_ net8 cal_lut\[128\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_26_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1209_ _0697_ _0721_ _0722_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1826__CLK net13 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_55_505 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_47_186 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_62_123 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtemp1.dac.parallel_cells\[1\].vdac_batch._6_ temp1.dac.parallel_cells\[1\].vdac_batch._2_
+ temp1.dac.parallel_cells\[1\].vdac_batch.en_pupd VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_14_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_120 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_38_164 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1431__A2 _0805_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1560_ _0303_ _0164_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_34_381 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1491_ _0275_ _0123_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_39_67 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1498__A2 _0779_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1849__CLK clknet_1_1__leaf_io_in[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_11 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_77_630 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_88 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_145 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1827_ _0179_ net2 cal_lut\[180\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1758_ _0110_ net15 cal_lut\[111\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1689_ _0041_ net16 cal_lut\[42\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_0_196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref_I temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1413__A2 _0240_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_240 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_251 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_307 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_50_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_295 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_381 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1177__A1 _0356_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0924__A1 _0357_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_384 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_74_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_204 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1101__A1 _0376_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_0991_ cal_lut\[81\] _0517_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1404__A2 _0802_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_123 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_68 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_273 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1612_ ctr\[6\] clknet_1_1__leaf__0318_ _0323_ _0196_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_1_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_395 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1543_ _0297_ _0153_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1671__CLK net15 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_13 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_24 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1474_ cal_lut\[115\] _0240_ _0267_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_97_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_97_736 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtemp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[14\].pupd temp1.dac.parallel_cells\[4\].vdac_batch.en_pupd
+ temp1.dac.parallel_cells\[4\].vdac_batch.npu_pd temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__invz_2
XTAP_TAPCELL_ROW_80_647 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_356 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0997__A4 _0384_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_229 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_72_240 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_295 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1159__A1 ctr\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_170 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_temp1.dac.parallel_cells\[1\].vdac_batch._5__A1 temp1.dac.i_enable VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_233 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_343 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_28_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1634__A2 _0351_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_273 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1694__CLK net18 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1190_ _0356_ _0687_ _0700_ _0702_ _0704_ _0705_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_86_321 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_86_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_0974_ _0360_ cal_lut\[33\] _0373_ _0500_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_1526_ cal_lut\[143\] _0255_ _0291_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_65_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1457_ _0262_ _0102_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1388_ _0231_ _0064_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_2_214 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1092__A3 _0413_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_262 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_192 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1304__A1 cal_lut\[17\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xdec1._102_ dec1._000_ dec1._002_ dec1._041_ dec1.o_dec\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_28_207 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_22_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_26 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_243 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_298 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0897__A3 _0422_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1311_ _0554_ _0791_ _0022_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_10_Right_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1242_ temp1.dac.i_data\[4\] _0709_ _0684_ _0753_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_39_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1173_ _0681_ _0686_ _0682_ _0688_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XTAP_TAPCELL_ROW_47_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_207 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_151 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_413 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_81 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_156 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0957_ cal_lut\[146\] _0484_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_6_189 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_42_243 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0888_ _0412_ _0414_ _0415_ _0416_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_2_384 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_140 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1509_ _0284_ _0132_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1273__I _0779_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_302 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_151 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_143 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_368 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_12_Left_110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1732__CLK net18 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0879__A3 _0363_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_25 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_151 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_335 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1860_ _0212_ clknet_1_0__leaf_io_in[0] dec1.i_ones VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_56_379 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1791_ _0143_ net12 cal_lut\[144\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_58_66 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_99 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1225_ _0345_ _0694_ _0737_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_416 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1156_ _0677_ _0678_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_0_74_98 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1087_ _0360_ _0608_ _0422_ _0609_ _0610_ _0611_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_0_59_151 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_31 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_368 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_305 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1755__CLK net13 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xtemp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[0\].vref temp1.dac.parallel_cells\[2\].vdac_batch.en_vref
+ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__invz_3
XFILLER_0_2_170 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_58_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_89_694 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1010_ _0534_ _0445_ _0535_ _0536_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_76_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1778__CLK net8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_78 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1843_ _0195_ clknet_1_0__leaf_io_in[0] dbg3\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1774_ _0126_ net8 cal_lut\[127\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_213 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_279 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_76 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_85_53 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_85_97 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1208_ seg1.o_segments\[2\] _0691_ _0721_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_55_506 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_246 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1139_ _0657_ _0659_ _0660_ _0661_ _0662_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_67_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_121 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_63_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_290 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_327 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_349 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_157 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_290 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtemp1.dac.parallel_cells\[1\].vdac_batch._5_ temp1.dac.i_enable temp1.dac.parallel_cells\[1\].vdac_batch._1_
+ temp1.dac.parallel_cells\[1\].vdac_batch._2_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_86_675 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_216 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_305 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_26 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_53_146 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_416 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_190 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1490_ cal_lut\[123\] _0255_ _0275_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_49_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_8_Right_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_71_44 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_17_296 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_99 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_349 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_360 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1826_ _0178_ net13 cal_lut\[179\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1757_ _0109_ net15 cal_lut\[110\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_96_41 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1688_ _0040_ net16 cal_lut\[41\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_39_Right_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_67_205 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtemp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[7\].pupd temp1.dac.parallel_cells\[4\].vdac_batch.en_pupd
+ temp1.dac.parallel_cells\[4\].vdac_batch.npu_pd temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__invz_2
XTAP_TAPCELL_ROW_0_197 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_48_Right_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_35_168 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1177__A2 _0357_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_57_Right_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_8_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[14\].vref_I temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_74_612 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1101__A2 _0391_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_66_Right_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_4_Left_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_41_14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1140__B _0384_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_0990_ cal_lut\[159\] _0516_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_41_138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1611_ _0368_ clknet_1_1__leaf__0318_ _0782_ _0323_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_1_224 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_202 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1816__CLK net14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_75_Right_75 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1542_ cal_lut\[153\] _0294_ _0297_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1473_ _0266_ _0114_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__0915__A2 _0401_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_97_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input2_I io_in[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_66 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1340__A2 _0802_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_32 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_84_Right_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_10_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_59_Left_157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_9_346 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0851__A1 _0376_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_260 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_80 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_93_Right_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_32_138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_13_341 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1809_ _0161_ net11 cal_lut\[162\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1276__I _0779_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_68_Left_166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_5_234 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_358 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1095__A1 _0376_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_77_Left_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__0842__A1 _0362_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xtemp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[14\].vref temp1.dac.parallel_cells\[4\].vdac_batch.en_vref
+ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__invz_3
XFILLER_0_63_230 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_39 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1839__CLK net12 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1398__A2 _0802_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_86_Left_184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1570__A2 _0289_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1322__A2 _0780_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_95_Left_193 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_39_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0973_ _0497_ _0498_ _0499_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__1389__A2 _0791_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_263 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_171 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1525_ _0570_ _0289_ _0142_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1561__A2 _0294_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_76 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1456_ cal_lut\[102\] _0255_ _0262_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_93_31 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1387_ cal_lut\[64\] _0802_ _0231_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_93_64 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_2_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1077__B2 cal_lut\[23\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1077__A1 cal_lut\[89\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1092__A4 _0406_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_230 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_187 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_274 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1552__A2 _0289_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1304__A2 _0780_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xdec1._101_ dec1.i_tens dec1._040_ dec1._041_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1661__CLK net17 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1310_ _0510_ _0790_ _0021_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1241_ _0368_ _0687_ _0704_ _0751_ _0752_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_1172_ _0681_ _0686_ _0682_ _0687_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_2_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_23 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_464 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_311 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_322 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_45 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1059__A1 _0368_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_377 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_74_314 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_358 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_124 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_6_168 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0956_ _0482_ _0432_ _0433_ _0483_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__1231__A1 temp1.dac.i_data\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_0887_ _0359_ cal_lut\[91\] _0394_ _0415_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_88_75 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1534__A2 _0289_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_185 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1508_ cal_lut\[132\] _0255_ _0284_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_49_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1439_ cal_lut\[94\] _0805_ _0253_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__1298__A1 cal_lut\[12\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1684__CLK net11 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_21_320 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1222__A1 _0357_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_277 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0981__B1 _0397_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1525__A2 _0289_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0879__A4 _0406_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_44_445 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_314 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_temp1.dac._5__A2 temp1.dac.i_data\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1790_ _0142_ net12 cal_lut\[143\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_24_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_233 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_266 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1516__A2 _0255_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1224_ _0697_ _0735_ _0736_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1155_ dec1.i_tens _0674_ _0675_ _0676_ _0677_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_1086_ cal_lut\[167\] _0610_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_47_325 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_347 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[1\].vref_I temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_65 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1549__I _0300_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_350 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0939_ cal_lut\[20\] _0466_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_30_236 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_58_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_314 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_358 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_147 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_394 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_89_695 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_225 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_269 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_291 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_369 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1842_ _0194_ clknet_1_1__leaf_io_in[0] dbg3\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_56_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_47 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1773_ _0125_ net10 cal_lut\[126\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_52_372 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_31_Left_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_85_21 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_40_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_81 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1207_ _0357_ _0495_ _0691_ _0496_ _0720_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_TAPCELL_ROW_55_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_258 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_40_Left_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1138_ cal_lut\[144\] _0626_ _0392_ cal_lut\[126\] _0661_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1069_ _0360_ _0413_ _0592_ _0593_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XTAP_TAPCELL_ROW_63_551 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1722__CLK net9 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_306 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_103 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_380 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_125 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0936__B1 _0397_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xtemp1.dac.parallel_cells\[1\].vdac_batch._4_ temp1.dac.i_data\[1\] temp1.dac.i_data\[5\]
+ temp1.dac.parallel_cells\[1\].vdac_batch._1_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_86_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_28 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_144 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_155 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_39_36 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_58 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_68 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1745__CLK net12 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_17_297 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_133 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_155 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_291 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_103 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_60_532 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_339 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_222 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1825_ _0177_ net14 cal_lut\[178\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_88_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_372 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1756_ _0108_ net15 cal_lut\[109\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1687_ _0039_ net16 cal_lut\[40\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1646__A1 temp1.dac.i_enable VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_217 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_70 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_0_198 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_253 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_342 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1768__CLK net12 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_74_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1637__A1 _0783_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_49 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1140__C _0390_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xtemp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[7\].vref temp1.dac.parallel_cells\[4\].vdac_batch.en_vref
+ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__invz_3
XANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[4\].vref_I temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_253 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1610_ _0345_ clknet_1_0__leaf__0318_ _0322_ _0195_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1541_ _0296_ _0152_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1472_ cal_lut\[114\] _0240_ _0266_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__0915__A3 _0440_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_97_738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_77 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_314 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__0851__A2 _0378_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_415 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1808_ _0160_ net15 cal_lut\[161\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_79_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_40_150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_40_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1739_ _0091_ net16 cal_lut\[92\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_28_359 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_220 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_264 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_94_719 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0972_ _0368_ cal_lut\[135\] _0370_ _0498_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_6_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_39_294 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_231 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_415 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_312 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1524_ _0526_ _0289_ _0141_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1010__A2 _0445_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_55 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1455_ _0261_ _0101_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_93_10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1386_ _0230_ _0063_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_2_216 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_dec1._070__A1 dec1.i_bin\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_70 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_33_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_267 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_312 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xdec1._100_ dec1._033_ dec1._038_ dec1._039_ dec1._040_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XANTENNA__1068__A2 _0355_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1806__CLK net16 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_39 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_348 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_231 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1240_ _0688_ _0749_ _0750_ _0687_ _0751_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_1171_ net6 _0686_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XANTENNA__1059__A2 _0357_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_47_465 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_345 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_90_700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_348 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_103 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_286 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0955_ cal_lut\[140\] _0482_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_12_83 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0886_ _0359_ _0366_ _0355_ _0413_ _0414_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XANTENNA__1231__A2 _0709_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_32 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_43 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_153 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1507_ _0283_ _0131_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_56_4 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_197 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1438_ _0252_ _0093_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1298__A2 _0780_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1829__CLK net17 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1369_ _0222_ _0054_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_37_80 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_418 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_120 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_77_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_337 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_21_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1470__A2 _0255_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_286 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_131 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_44_446 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_337 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1461__A2 _0791_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_52_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_1_1__f__0318_ clknet_0__0318_ clknet_1_1__leaf__0318_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_3_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0972__A1 _0368_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1223_ seg1.o_segments\[3\] _0691_ _0735_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_74_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_45 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1154_ ctr\[8\] ctr\[10\] ctr\[11\] _0676_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1085_ _0376_ _0362_ _0364_ _0406_ _0609_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_59_131 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_337 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1452__A2 _0255_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout16_I net18 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_189 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0938_ cal_lut\[44\] _0465_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_15_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0869_ _0358_ _0366_ _0355_ _0396_ _0397_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XANTENNA__1651__CLK net11 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_326 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_123 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_38_348 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_89_696 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_59 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_337 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1841_ _0193_ clknet_1_0__leaf_io_in[0] dbg3\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1772_ _0124_ net10 cal_lut\[125\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_52_384 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1674__CLK net15 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_270 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_88 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1206_ _0346_ _0672_ _0708_ _0710_ _0719_ io_out[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_1137_ cal_lut\[174\] _0625_ _0389_ cal_lut\[168\] _0660_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_55_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1068_ _0366_ _0355_ _0592_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_63_552 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_123 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_134 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1425__A2 _0791_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_286 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xtemp1.dac.parallel_cells\[1\].vdac_batch._3_ temp1.dac.i_data\[1\] temp1.dac.parallel_cells\[1\].vdac_batch.npu_pd
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_86_677 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0872__B1 _0392_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_251 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_93_295 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_284 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1697__CLK net18 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0927__A1 _0368_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_373 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_192 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1407__A2 _0240_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_17_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_60_533 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_340 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1824_ _0176_ net2 cal_lut\[177\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_4_234 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1755_ _0107_ net13 cal_lut\[108\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__0918__A1 _0376_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_181 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1040__B1 _0423_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1686_ _0038_ net16 cal_lut\[39\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_24_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_229 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_0_199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_273 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_232 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_148 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_16_373 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0909__A1 _0376_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1031__B1 _0403_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_376 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_17 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_74_614 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_295 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0832__I _0359_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_221 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_265 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_170 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_276 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1540_ cal_lut\[152\] _0294_ _0296_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__1022__B1 _0386_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_226 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_16 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1471_ _0265_ _0113_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1712__CLK net11 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_97_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_207 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_57_295 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1807_ _0159_ net16 cal_lut\[160\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_25_192 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1013__B1 _0433_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1738_ _0090_ net16 cal_lut\[91\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1669_ _0021_ net17 cal_lut\[22\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_95_335 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1095__A3 _0391_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_251 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_381 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_170 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1735__CLK net18 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_173 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0827__I _0355_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_temp1.dac.parallel_cells\[1\].vdac_batch.einvp_batch\[1\].vref_I temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_0971_ cal_lut\[153\] _0452_ _0497_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_14_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_10_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1546__A1 cal_lut\[155\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1523_ _0482_ _0791_ _0140_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1607__B _0782_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_9 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1454_ cal_lut\[101\] _0240_ _0261_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_77_67 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1385_ cal_lut\[63\] _0805_ _0230_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_2_217 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_189 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_33_385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_81 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_33_405 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1758__CLK net15 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_368 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1170_ _0347_ _0677_ _0685_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_63_14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_90_701 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_221 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_148 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0954_ _0471_ _0474_ _0477_ _0480_ _0481_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_12_73 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_235 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0885_ _0396_ _0413_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_82_382 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1519__A1 _0608_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1506_ cal_lut\[131\] _0255_ _0283_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1437_ cal_lut\[93\] _0805_ _0252_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1368_ cal_lut\[54\] _0802_ _0222_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_37_92 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_38_411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1299_ _0793_ _0012_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xtemp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].pupd temp1.dac.parallel_cells\[3\].vdac_batch.en_pupd
+ temp1.dac.parallel_cells\[3\].vdac_batch.npu_pd temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__invz_2
XFILLER_0_53_91 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_243 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_349 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_21_322 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_279 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0981__A2 _0395_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_290 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_44_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_327 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_187 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_146 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_135 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_52_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_308 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_393 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_64_382 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0840__I _0358_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1222_ _0357_ _0539_ _0691_ _0540_ _0734_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1153_ ctr\[12\] _0675_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
X_1084_ cal_lut\[137\] _0608_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_74_102 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_349 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_202 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_179 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0937_ cal_lut\[164\] _0389_ _0392_ cal_lut\[122\] _0463_ _0464_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_15_224 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_279 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_238 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0868_ _0362_ _0363_ _0396_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_23_290 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_151 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_41_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].vref_I temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_249 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1131__A2 _0452_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0890__A1 _0359_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_102 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_349 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_360 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1840_ _0192_ clknet_1_1__leaf_io_in[0] dbg3\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_71_138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1771_ _0123_ net10 cal_lut\[124\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1819__CLK net14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_205 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_49 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_57 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1370__A2 _0805_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1205_ _0365_ _0687_ _0704_ _0718_ _0719_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_2
Xclkbuf_1_0__f_temp1.i_precharge_n clknet_0_temp1.i_precharge_n clknet_1_0__leaf_temp1.i_precharge_n
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_55_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1136_ cal_lut\[180\] _0658_ _0402_ cal_lut\[186\] _0659_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1067_ _0390_ _0363_ cal_lut\[29\] _0384_ _0591_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_TAPCELL_ROW_63_553 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_260 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_360 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_168 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_382 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_190 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0936__A2 _0395_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_86_678 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_102 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_113 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_271 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_146 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_274 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_263 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_157 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_168 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_371 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_182 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1352__A2 _0790_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_15 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0863__A1 _0365_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_146 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_230 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_17_299 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_60_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_263 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_202 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1823_ _0175_ net14 cal_lut\[176\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1754_ _0106_ net9 cal_lut\[107\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1791__CLK net12 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_279 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_333 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1040__A1 _0376_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1685_ _0037_ net16 cal_lut\[38\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1591__A2 _0294_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch._7__I temp1.dac.i_enable VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1343__A2 _0790_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1119_ _0368_ cal_lut\[138\] _0370_ _0642_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__0854__A1 _0365_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_83_659 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_50 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_75_241 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_90_200 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_17_Right_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_90_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_299 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1334__A2 _0805_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_26_Right_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__0845__A1 _0362_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1664__CLK net14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_241 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_35_Right_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_66_285 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_311 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_193 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_377 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1470_ cal_lut\[113\] _0255_ _0265_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__1165__B _0678_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_28 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_44_Right_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1325__A2 _0802_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_19_Left_117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_15_84 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_53_Right_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_57_241 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_414 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_28_Left_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1261__A1 _0346_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_255 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_119 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1806_ _0158_ net16 cal_lut\[159\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1013__A1 _0499_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1737_ _0089_ net16 cal_lut\[90\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_185 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_62_Right_62 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1668_ _0020_ net17 cal_lut\[21\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1599_ _0615_ _0780_ _0191_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_37_Left_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1316__A2 _0783_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1687__CLK net16 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_347 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1095__A4 _0413_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_71_Right_71 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_48_241 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_46_Left_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_16_160 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_266 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_277 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1555__A2 _0294_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_80_Right_80 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_55_Left_153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_86_314 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_64_Left_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_0970_ _0357_ _0495_ _0496_ dec1.i_bin\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_TAPCELL_ROW_10_261 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_185 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_163 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_314 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1546__A2 _0294_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1522_ _0431_ _0289_ _0139_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_73_Left_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1453_ _0260_ _0100_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1384_ _0229_ _0062_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_2_218 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_82_Left_180 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_42_71 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_179 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1234__A1 _0357_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_33_386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_266 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_60_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_314 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_325 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_380 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1702__CLK net8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1225__A1 _0345_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_203 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1852__CLK clknet_1_1__leaf_io_in[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1528__A2 _0255_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0838__I _0365_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_90_702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_369 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_417 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xdec1._089_ dec1._008_ dec1._003_ dec1._029_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_0953_ _0478_ _0427_ _0479_ _0480_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_30_367 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0884_ cal_lut\[7\] _0412_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_42_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1618__B _0783_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1519__A2 _0289_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_67 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_133 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_144 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1505_ _0282_ _0130_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1436_ _0251_ _0092_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1367_ _0221_ _0053_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_38_412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_0_io_in[0]_I io_in[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1298_ cal_lut\[12\] _0780_ _0793_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__1725__CLK net15 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_144 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_155 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_166 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1207__A1 _0357_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_266 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_255 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_309 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_171 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_155 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_44_448 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_52_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_1_1__f__0316_ clknet_0__0316_ clknet_1_1__leaf__0316_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xtemp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].vref temp1.dac.parallel_cells\[3\].vdac_batch.en_vref
+ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__invz_3
XANTENNA__0972__A3 _0370_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1221_ ctr\[11\] _0733_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__1748__CLK net12 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_58 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1152_ ctr\[9\] _0674_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1083_ _0601_ _0603_ _0605_ _0606_ _0607_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_62_309 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_169 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0936_ _0461_ _0395_ _0397_ _0462_ _0463_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_0_30_228 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0867_ _0358_ _0394_ _0395_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_2_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_185 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1419_ _0517_ _0791_ _0081_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1125__B1 _0379_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_3_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_41_429 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_29 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_306 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_125 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_temp1.dac.parallel_cells\[0\].vdac_batch._4__A1 temp1.dac.i_data\[0\] VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_309 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1770_ _0122_ net10 cal_lut\[123\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_52_364 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_261 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_95 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1204_ _0688_ _0716_ _0717_ _0687_ _0718_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_1135_ _0445_ _0658_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_79_228 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1066_ cal_lut\[107\] _0589_ _0590_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_87_272 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_372 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0919_ _0444_ _0445_ _0446_ _0447_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_70_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_272 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_294 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_0__0318_ _0318_ clknet_0__0318_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_86_679 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0872__A2 _0389_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_136 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtemp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[2\].pupd temp1.dac.parallel_cells\[4\].vdac_batch.en_pupd
+ temp1.dac.parallel_cells\[4\].vdac_batch.npu_pd temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__invz_2
XANTENNA__0927__A3 _0370_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1104__A3 _0627_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0863__A2 _0355_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_60_535 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_242 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1822_ _0174_ net14 cal_lut\[175\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1753_ _0105_ net10 cal_lut\[106\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_4_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_40_312 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_74 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1684_ _0036_ net11 cal_lut\[37\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__0918__A3 _0413_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_78 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_96_45 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_50 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1118_ _0639_ _0395_ _0640_ _0641_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__0854__A2 _0355_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1049_ _0572_ _0436_ _0573_ _0574_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_50_109 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_312 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0909__A3 _0391_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1031__A2 _0402_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1809__CLK net11 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_18 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1270__A2 _0684_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_245 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1022__A2 _0383_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xseg1._49_ dec1.o_dec\[2\] seg1._13_ seg1._12_ seg1._19_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_89_345 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_52 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_57_231 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_253 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_286 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_40 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_223 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_84 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_407 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1805_ _0157_ net16 cal_lut\[158\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_120 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1736_ _0088_ net18 cal_lut\[89\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1667_ _0019_ net17 cal_lut\[20\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1598_ _0549_ _0780_ _0190_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_96_730 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_415 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_201 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_256 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_120 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_153 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_29 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_19_307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1781__CLK net8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0818__A2 ctr\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_27_351 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_381 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_286 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_234 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_407 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_10_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1521_ _0290_ _0138_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1452_ cal_lut\[100\] _0255_ _0260_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_77_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1383_ cal_lut\[62\] _0805_ _0229_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_26_62 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_89_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_77_348 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1482__A2 _0255_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_234 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_407 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_186 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1719_ _0071_ net11 cal_lut\[72\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1654__CLK net15 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xtemp1.dac.parallel_cells\[4\].vdac_batch._8_ temp1.dac.parallel_cells\[4\].vdac_batch._0_
+ temp1.dac.parallel_cells\[4\].vdac_batch._1_ temp1.dac.parallel_cells\[4\].vdac_batch.en_vref
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__1105__I cal_lut\[161\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_134 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_223 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_340 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1161__A1 _0345_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_16 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_326 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_337 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1464__A2 _0240_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_348 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0952_ _0390_ _0363_ cal_lut\[26\] _0384_ _0479_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__1216__A2 _0709_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_53 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xdec1._088_ dec1._007_ dec1._013_ dec1._015_ dec1._028_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and3_2
XANTENNA__0975__A1 _0368_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_30_368 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1677__CLK net11 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_0883_ cal_lut\[181\] _0402_ _0403_ cal_lut\[49\] _0410_ _0411_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_82_384 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_301 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_9 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_79 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1504_ cal_lut\[130\] _0255_ _0282_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_2_378 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1435_ cal_lut\[92\] _0240_ _0251_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1366_ cal_lut\[53\] _0802_ _0221_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_37_61 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_38_413 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1297_ _0792_ _0011_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_53_82 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1143__A1 _0368_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_69_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_1_Left_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1446__A2 _0240_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_123 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_44_449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_384 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_281 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1134__A1 cal_lut\[42\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1151_ _0346_ ctr\[1\] _0673_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_74_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1082_ cal_lut\[185\] _0402_ _0403_ cal_lut\[53\] _0606_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__1437__A2 _0805_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_329 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_dec1._060__I dec1.i_bin\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_0935_ cal_lut\[104\] _0462_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_70_310 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0866_ _0362_ _0363_ _0365_ _0355_ _0394_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
XFILLER_0_70_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_2_153 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1418_ _0473_ _0791_ _0080_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1349_ _0214_ _0042_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1842__CLK clknet_1_1__leaf_io_in[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_92 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1428__A2 _0790_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_46_384 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_229 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1419__A2 _0791_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0890__A3 _0355_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_temp1.dac.parallel_cells\[0\].vdac_batch._4__A2 temp1.dac.i_data\[5\] VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_118 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_52_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[7\].vref_I temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1715__CLK net9 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1107__A1 _0360_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1203_ ctr\[1\] _0688_ _0717_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_85_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1134_ cal_lut\[42\] _0586_ _0593_ cal_lut\[18\] _0657_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1065_ _0397_ _0589_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_75_413 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_251 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout14_I net2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_321 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0918_ _0376_ cal_lut\[115\] _0413_ _0406_ _0446_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_0849_ _0376_ _0367_ _0377_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__1346__A1 cal_lut\[41\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_54_500 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_221 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_170 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_416 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtemp1.dcdc temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_ clknet_1_1__leaf_temp1.i_precharge_n
+ temp1.dcdel_capnode_notouch_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__invz_1
XANTENNA__1738__CLK net16 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_17 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtemp1.dac.vdac_single._4__20 net20 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_29_137 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_284 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_273 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_148 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_159 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0862__I _0362_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_60_536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1821_ _0173_ net14 cal_lut\[174\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_25_332 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1752_ _0104_ net10 cal_lut\[105\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_4_226 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_140 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_151 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1683_ _0035_ net11 cal_lut\[36\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__0918__A4 _0406_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1040__A3 _0422_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xtemp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[2\].vref temp1.dac.parallel_cells\[4\].vdac_batch.en_vref
+ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__invz_3
XFILLER_0_0_410 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_61 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1117_ cal_lut\[84\] _0602_ _0640_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1048_ _0358_ cal_lut\[100\] _0391_ _0413_ _0573_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_48_413 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtemp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[1\].pupd temp1.dac.parallel_cells\[2\].vdac_batch.en_pupd
+ temp1.dac.parallel_cells\[2\].vdac_batch.npu_pd temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__invz_2
XTAP_TAPCELL_ROW_16_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_3_Right_3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_63_416 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_321 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__0909__A4 _0413_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_346 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_368 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_8_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0845__A3 _0365_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_170 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_257 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_162 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xseg1._48_ seg1._18_ seg1.o_segments\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_82_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_31 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_86 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1246__B1 _0635_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1804_ _0156_ net16 cal_lut\[157\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1013__A3 _0538_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1735_ _0087_ net18 cal_lut\[88\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_187 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1666_ _0018_ net17 cal_lut\[19\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1597_ _0505_ _0780_ _0189_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_0_240 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_96_731 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_82 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_349 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_70 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_373 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_246 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_279 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_290 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_19_308 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_276 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_298 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1520_ cal_lut\[138\] _0779_ _0290_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1451_ _0259_ _0099_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1382_ _0228_ _0061_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1192__B _0684_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_41 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_26_74 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_246 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1718_ _0070_ net11 cal_lut\[71\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1649_ _0001_ net8 cal_lut\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xtemp1.dac.parallel_cells\[4\].vdac_batch._7_ temp1.dac.i_enable temp1.dac.parallel_cells\[4\].vdac_batch._0_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1170__A2 _0677_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_8_181 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_168 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0951_ cal_lut\[110\] _0478_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xdec1._087_ dec1.i_bin\[2\] dec1._027_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_27_257 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_30_369 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_216 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0882_ _0404_ _0407_ _0408_ _0409_ _0410_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_0_2_313 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_290 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_346 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_50_260 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtemp1.inv1_2 temp1.dcdel_capnode_notouch_ net23 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_10_102 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1503_ _0281_ _0129_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_10_146 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1434_ _0250_ _0091_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1365_ _0220_ _0052_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_38_414 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1296_ cal_lut\[11\] _0780_ _0792_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_53_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_85_190 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1771__CLK net10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xtemp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[15\].pupd temp1.dac.parallel_cells\[4\].vdac_batch.en_pupd
+ temp1.dac.parallel_cells\[4\].vdac_batch.npu_pd temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__invz_2
XTAP_TAPCELL_ROW_69_583 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_102 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_135 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_308 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_127 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_374 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_411 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1150_ ctr\[1\] _0672_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_4
X_1081_ cal_lut\[155\] _0452_ _0604_ cal_lut\[47\] _0605_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_temp1.dac.parallel_cells\[2\].vdac_batch._5__A1 temp1.dac.i_enable VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_146 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_416 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_149 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0934_ cal_lut\[188\] _0461_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1794__CLK net13 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_0865_ cal_lut\[187\] _0393_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1070__B2 cal_lut\[17\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_121 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_260 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1645__B dec1.i_tens VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1417_ _0419_ _0790_ _0079_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1348_ cal_lut\[42\] _0802_ _0214_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1279_ _0784_ _0001_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_58_190 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_208 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1600__A3 _0677_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1364__A2 _0802_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_57_520 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1667__CLK net17 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0875__A1 _0362_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_241 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_127 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_171 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_193 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_230 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_263 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1202_ _0674_ _0715_ _0690_ _0716_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1133_ _0641_ _0646_ _0649_ _0655_ _0656_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
XANTENNA__0866__A1 _0362_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1064_ cal_lut\[41\] _0586_ _0587_ cal_lut\[11\] _0588_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA_dec1._071__I dec1.i_bin\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_41 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_311 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_300 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_119 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_344 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0917_ _0358_ _0366_ _0355_ _0385_ _0445_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_70_152 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0848_ _0358_ _0376_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_70_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1346__A2 _0802_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_263 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_252 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_296 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_0__0316_ _0316_ clknet_0__0316_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_52_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0857__A1 _0362_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_54_501 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_241 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_263 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_266 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_300 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_377 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_130 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1585__A2 _0294_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_77_626 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_85_670 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_241 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xtemp1.dac.vdac_single._4__21 net21 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_TAPCELL_ROW_60_537 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1220__1 clknet_1_1__leaf_io_in[0] net22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_84_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1820_ _0172_ net14 cal_lut\[173\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1751_ _0103_ net10 cal_lut\[104\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_4_238 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1576__A2 _0289_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1682_ _0034_ net11 cal_lut\[35\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_314 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_185 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_98 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1832__CLK net17 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__0839__A1 _0362_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1500__A2 _0779_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1116_ cal_lut\[192\] _0639_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1047_ cal_lut\[148\] _0572_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1264__A1 _0357_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_16_291 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_333 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_171 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_193 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_314 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_8_248 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0845__A4 _0356_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1705__CLK net8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1255__A1 _0346_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_255 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_299 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1855__CLK clknet_1_0__leaf_io_in[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xtemp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[1\].vref temp1.dac.parallel_cells\[2\].vdac_batch.en_vref
+ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__invz_3
XFILLER_0_22_325 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_303 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xseg1._47_ seg1._16_ seg1._17_ seg1._18_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XPHY_EDGE_ROW_13_Right_13 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_89_325 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtemp1.dac.parallel_cells\[0\].vdac_batch.einvp_batch\[0\].pupd temp1.dac.parallel_cells\[0\].vdac_batch.en_pupd
+ temp1.dac.parallel_cells\[0\].vdac_batch.npu_pd temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__invz_2
XFILLER_0_15_76 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_288 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_42 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_299 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_22_Right_22 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_31_64 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1803_ _0155_ net12 cal_lut\[156\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_13_325 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_40_100 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1734_ _0086_ net18 cal_lut\[87\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_166 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1665_ _0017_ net14 cal_lut\[18\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_380 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1596_ _0461_ _0780_ _0188_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_0_274 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_31_Right_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_96_732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1728__CLK net16 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_40_Right_40 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_16_141 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_269 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_185 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_15_Left_113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_31_144 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_24_Left_122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_19_309 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1228__A1 ctr\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_417 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_225 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_33_Left_131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_22_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_155 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_199 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1450_ cal_lut\[99\] _0255_ _0259_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1381_ cal_lut\[61\] _0805_ _0228_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XPHY_EDGE_ROW_42_Left_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_77_306 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_166 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1219__B2 clknet_1_1__leaf_io_in[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_258 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1717_ _0069_ net11 cal_lut\[70\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1648_ _0000_ net8 cal_lut\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_6_30 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1579_ _0578_ _0780_ _0178_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xtemp1.dac.parallel_cells\[4\].vdac_batch._6_ temp1.dac.parallel_cells\[4\].vdac_batch._2_
+ temp1.dac.parallel_cells\[4\].vdac_batch.en_pupd VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_1_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_24_334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_372 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1630__A1 ctr\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].vref_I temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xtemp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[8\].pupd temp1.dac.parallel_cells\[4\].vdac_batch.en_pupd
+ temp1.dac.parallel_cells\[4\].vdac_batch.npu_pd temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__invz_2
XFILLER_0_59_328 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_147 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_225 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0950_ _0376_ _0475_ _0422_ _0423_ _0476_ _0477_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai32_2
Xdec1._086_ dec1._016_ dec1._025_ dec1.i_bin\[2\] dec1._026_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XANTENNA__0975__A3 _0373_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_228 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0881_ cal_lut\[19\] _0409_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_12_99 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_239 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1502_ cal_lut\[129\] _0779_ _0281_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1433_ cal_lut\[91\] _0240_ _0250_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_10_169 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1137__B1 _0389_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_41 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1364_ cal_lut\[52\] _0802_ _0220_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_37_85 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1295_ _0557_ _0791_ _0010_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_38_415 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_136 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_84 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_95 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_58_350 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1143__A3 _0373_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_69_584 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_372 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1603__A1 _0355_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_283 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1080_ _0376_ _0362_ _0364_ _0382_ _0604_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_59_125 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_27 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtemp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[15\].vref temp1.dac.parallel_cells\[4\].vdac_batch.en_vref
+ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__invz_3
XTAP_TAPCELL_ROW_43_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xdec1._069_ dec1.i_bin\[5\] dec1._009_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_0933_ _0456_ _0457_ _0458_ _0459_ _0460_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_82_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0864_ _0376_ _0390_ _0363_ _0391_ _0392_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XANTENNA__1070__A2 _0383_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_334 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_23_272 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_294 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1416_ _0245_ _0078_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1347_ _0213_ _0041_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_3_42 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1278_ cal_lut\[1\] _0783_ _0784_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_66_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_312 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_356 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_401 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_69_Right_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_49_191 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_7_Left_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_52_312 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1052__A2 _0401_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_242 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_78_Right_78 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1201_ _0711_ _0713_ _0714_ _0715_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1107__A3 _0378_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1132_ _0650_ _0651_ _0652_ _0654_ _0655_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__0866__A2 _0363_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_88_690 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1063_ _0360_ _0366_ _0355_ _0413_ _0587_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__1761__CLK net15 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_264 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_87_Right_87 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_87_286 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1291__A2 _0790_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_161 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0916_ cal_lut\[175\] _0444_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_43_356 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_367 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_96_Right_96 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_0847_ _0368_ cal_lut\[127\] _0373_ _0375_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_11_275 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0857__A2 _0363_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_54_502 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_117 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1282__A2 _0783_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_89_Left_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_77_627 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1784__CLK net10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_85_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_267 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1750_ _0102_ net10 cal_lut\[103\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_37_194 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1681_ _0033_ net8 cal_lut\[34\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_96_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_dec1._085__A1 dec1.i_bin\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1115_ _0585_ _0357_ _0638_ dec1.i_bin\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_1046_ _0570_ _0432_ _0433_ _0571_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_16_292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_109 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1016__A2 _0452_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_301 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_367 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_326 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1657__CLK net15 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_249 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_404 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_183 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1007__A2 _0401_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xseg1._46_ dec1.o_dec\[1\] dec1.o_dec\[0\] dec1.o_dec\[2\] seg1._11_ seg1._17_ VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_30_381 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_18 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1191__A1 temp1.dac.i_data\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_28 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1494__A2 _0255_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_245 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_418 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_256 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[10\].vref_I temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_215 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1802_ _0154_ net10 cal_lut\[155\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_72_259 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_87 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1733_ _0085_ net18 cal_lut\[86\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1664_ _0016_ net14 cal_lut\[17\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1595_ _0393_ _0780_ _0187_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_96_733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_4 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_50 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1029_ cal_lut\[22\] _0554_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_36_407 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xtemp1.dac.parallel_cells\[0\].vdac_batch.einvp_batch\[0\].vref temp1.dac.parallel_cells\[0\].vdac_batch.en_vref
+ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__invz_3
XANTENNA__1135__I _0445_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1476__A2 _0240_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_27_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1822__CLK net14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_101 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1400__A2 _0802_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_189 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xseg1._29_ dec1.o_dec\[2\] seg1._03_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
X_1380_ _0227_ _0060_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1164__A1 _0346_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_93_714 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_32 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1467__A2 _0790_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_340 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_226 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_334 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_53_270 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1716_ _0068_ net8 cal_lut\[69\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1647_ _0783_ _0342_ _0212_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1155__A1 dec1.i_tens VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1578_ _0534_ _0780_ _0177_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_67_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xtemp1.dac.parallel_cells\[4\].vdac_batch._5_ temp1.dac.i_enable temp1.dac.parallel_cells\[4\].vdac_batch._1_
+ temp1.dac.parallel_cells\[4\].vdac_batch._2_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__1458__A2 _0791_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_1_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1845__CLK clknet_1_0__leaf_io_in[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_126 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_24_335 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_340 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0969__A1 _0363_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_215 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_384 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_207 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_temp1.dac._4__I temp1.dac.i_enable VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1146__A1 cal_lut\[12\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_19 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_318 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xdec1._085_ dec1.i_bin\[2\] dec1._018_ dec1._019_ dec1._023_ dec1._024_ dec1._025_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai32_4
XANTENNA__1082__B1 _0403_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_0880_ _0359_ _0396_ _0406_ _0408_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_82_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1718__CLK net11 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1501_ _0280_ _0128_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_10_137 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1432_ _0249_ _0090_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1137__B2 cal_lut\[168\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_20 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1363_ _0219_ _0051_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1294_ _0782_ _0791_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_38_416 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_46_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_77_159 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_384 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtemp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[8\].vref temp1.dac.parallel_cells\[4\].vdac_batch.en_vref
+ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__invz_3
XFILLER_0_18_259 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_78_93 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1128__A1 _0360_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_69_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_61_Left_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_68_137 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_159 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_70_Left_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_32_273 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1119__A1 _0368_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_148 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_39 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_43_441 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0932_ cal_lut\[68\] _0383_ _0386_ cal_lut\[74\] _0459_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_2
Xdec1._068_ dec1.i_bin\[4\] dec1._008_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_70_302 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0863_ _0365_ _0355_ _0391_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_2_101 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1690__CLK net17 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_189 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1415_ cal_lut\[78\] _0240_ _0245_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1346_ cal_lut\[41\] _0802_ _0213_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_3_76 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1277_ _0782_ _0783_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_66_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_416 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_181 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_14_273 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0875__A3 _0384_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_287 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_343 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_40_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1052__A3 _0440_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_368 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1200_ ctr\[3\] _0694_ _0714_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_18_77 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1131_ cal_lut\[156\] _0452_ _0653_ cal_lut\[162\] _0654_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__0866__A3 _0365_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_88_691 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1062_ _0368_ _0422_ _0586_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_28_321 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_310 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_31 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_173 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0915_ _0439_ _0401_ _0440_ _0441_ _0442_ _0443_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_0_70_154 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0846_ _0360_ cal_lut\[31\] _0373_ _0374_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_11_265 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1329_ _0782_ _0805_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_54_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_202 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_235 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_365 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_77_628 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_85_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_143 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1680_ _0032_ net8 cal_lut\[33\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_96_49 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1114_ _0635_ _0637_ _0638_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_48_405 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1045_ cal_lut\[142\] _0570_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_0_66 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_44 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_41 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_16_293 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_140 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_85 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout12_I net13 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_335 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_31 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_132 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_290 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_262 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0829_ _0356_ _0357_ dec1.i_bin\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_86_71 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_74_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_82_653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1007__A3 _0440_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_temp1.dac.parallel_cells\[3\].vdac_batch._7__I temp1.dac.i_enable VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xseg1._45_ dec1.o_dec\[2\] seg1._12_ seg1._09_ seg1._00_ seg1._13_ seg1._16_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__1751__CLK net10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_316 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_349 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1801_ _0153_ net10 cal_lut\[154\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_72_227 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_290 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1732_ _0084_ net18 cal_lut\[85\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_13_349 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_198 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1663_ _0015_ net17 cal_lut\[16\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1594_ _0315_ _0186_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_7_Right_7 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_96_734 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[0\].vref_I temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_319 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_48_202 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1028_ cal_lut\[46\] _0553_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_48_235 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_382 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1774__CLK net8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_157 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_97_70 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_27_355 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_290 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xseg1._28_ dec1.o_dec\[1\] seg1._01_ dec1.o_dec\[2\] seg1._02_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_10_308 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_93_715 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_135 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_77 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_308 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_168 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_18_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1797__CLK net12 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_216 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_302 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1227__I0 _0733_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1715_ _0067_ net9 cal_lut\[68\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_53_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_135 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1646_ temp1.dac.i_enable _0341_ _0342_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1577_ _0490_ _0780_ _0176_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xtemp1.dac.parallel_cells\[4\].vdac_batch._4_ temp1.dac.i_data\[4\] temp1.dac.i_data\[5\]
+ temp1.dac.parallel_cells\[4\].vdac_batch._1_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_1_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_308 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_336 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_227 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0969__A2 _0357_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_173 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_380 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1394__A2 _0805_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_171 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_385 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xdec1._084_ dec1.i_bin\[3\] dec1._006_ dec1._024_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_35_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1385__A2 _0805_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1500_ cal_lut\[128\] _0779_ _0280_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1431_ cal_lut\[90\] _0805_ _0249_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1362_ cal_lut\[51\] _0805_ _0219_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1293_ _0513_ _0790_ _0009_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_18_227 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_73_344 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_219 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0820__A1 _0345_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_4 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1376__A2 _0802_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1629_ _0783_ _0331_ _0205_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_68_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1812__CLK net13 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0887__A1 _0359_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_69_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1300__A2 _0790_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_311 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1064__A1 cal_lut\[41\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_43_442 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_119 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0931_ cal_lut\[56\] _0377_ _0379_ cal_lut\[62\] _0458_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_55_311 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_344 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xdec1._067_ dec1._004_ dec1._006_ dec1._007_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_0862_ _0362_ _0390_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_8
XFILLER_0_70_314 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_325 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_185 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1835__CLK net13 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1358__A2 _0805_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1414_ _0244_ _0077_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1345_ _0563_ _0791_ _0040_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__0869__A1 _0358_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1530__A2 _0289_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1276_ _0779_ _0782_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_4
XFILLER_0_64_96 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_66_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_119 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1597__A2 _0780_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_355 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_358 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_296 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_285 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_190 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_233 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_255 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1708__CLK net9 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1037__A1 _0359_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1858__CLK clknet_1_0__leaf_io_in[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_40_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_399 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_314 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_185 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_391 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_18_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_45 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1512__A2 _0255_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1130_ _0360_ _0378_ _0653_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__0866__A4 _0355_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1061_ dbg3\[5\] _0585_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_75_417 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_99 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xdec1._119_ dec1._002_ dec1._054_ dec1._055_ dec1._056_ dec1._017_ dec1.o_dec\[2\]
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai32_4
XANTENNA__1579__A2 _0780_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_0914_ cal_lut\[13\] _0442_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_0845_ _0362_ _0364_ _0365_ _0356_ _0373_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_50_87 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1200__A1 ctr\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_299 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_75_51 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1328_ _0804_ _0030_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1259_ _0766_ _0767_ _0759_ _0768_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_54_504 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1019__A1 _0360_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_314 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_369 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_391 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__0950__B1 _0423_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_77_629 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1258__A1 _0678_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_85_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtemp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[5\].pupd temp1.dac.parallel_cells\[3\].vdac_batch.en_pupd
+ temp1.dac.parallel_cells\[3\].vdac_batch.npu_pd temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__invz_2
XANTENNA__1680__CLK net8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_277 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_299 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_25_336 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1329__I _0782_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_155 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0941__B1 _0403_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0839__A4 _0355_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1113_ _0636_ _0637_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_45_32 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1249__A1 dec1.i_tens VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1044_ _0559_ _0562_ _0565_ _0568_ _0569_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_48_417 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_203 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_325 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_152 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_97 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_380 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0828_ net4 _0357_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__0932__B1 _0386_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_82_654 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_217 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_111 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xseg1._44_ seg1._03_ seg1._00_ seg1._08_ seg1.o_segments\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_15_46 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_68 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1800_ _0152_ net10 cal_lut\[153\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_25_100 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_13_275 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_133 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_45 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1731_ _0083_ net16 cal_lut\[84\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1662_ _0014_ net17 cal_lut\[15\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_372 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1593_ cal_lut\[186\] _0782_ _0315_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_56_31 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_96_735 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1027_ cal_lut\[166\] _0389_ _0392_ cal_lut\[124\] _0551_ _0552_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_48_214 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_111 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_166 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_103 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_294 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_136 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_383 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1633__A1 _0783_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_409 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xseg1._27_ dec1.o_dec\[0\] seg1._01_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_TAPCELL_ROW_93_716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_18_301 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_158 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_55 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1714_ _0066_ net9 cal_lut\[67\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_53_261 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1645_ _0675_ _0339_ dec1.i_tens _0341_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_6_66 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1576_ _0444_ _0289_ _0175_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1155__A3 _0675_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_99 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtemp1.dac.parallel_cells\[4\].vdac_batch._3_ temp1.dac.i_data\[4\] temp1.dac.parallel_cells\[4\].vdac_batch.npu_pd
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_3
XFILLER_0_83_40 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_95 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1741__CLK net15 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_24_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_239 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_32_381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_320 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xdec1._083_ dec1._011_ dec1._021_ dec1._022_ dec1._023_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__1606__A1 ctr\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xtemp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[10\].pupd temp1.dac.parallel_cells\[4\].vdac_batch.en_pupd
+ temp1.dac.parallel_cells\[4\].vdac_batch.npu_pd temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__invz_2
XFILLER_0_94_183 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1082__A2 _0402_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_378 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_294 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_220 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_242 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1430_ _0248_ _0089_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1361_ _0218_ _0050_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_37_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1292_ _0469_ _0790_ _0008_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1764__CLK net14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_87 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_275 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1628_ ctr\[6\] _0330_ _0331_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__1128__A3 _0373_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1559_ cal_lut\[164\] _0294_ _0303_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_91_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_91_197 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_294 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1119__A3 _0370_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1787__CLK net14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_19 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_43_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0930_ _0368_ cal_lut\[128\] _0373_ _0457_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__1055__A2 _0445_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xdec1._066_ dec1.i_bin\[6\] dec1._005_ dec1._006_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_0861_ _0359_ _0381_ _0382_ _0389_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_23_220 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_264 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1413_ cal_lut\[77\] _0240_ _0244_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1344_ _0519_ _0790_ _0039_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1275_ _0781_ _0000_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_3_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_66_568 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_323 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_161 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_183 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_164 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_348 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_14_242 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_29_Right_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_37_356 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_38_Right_38 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_64_197 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_60_370 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_234 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_278 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_47_Right_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[0\].vref_I temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1060_ _0357_ _0583_ _0584_ dec1.i_bin\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_34_45 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_63_549 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1802__CLK net10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xdec1._118_ dec1.i_tens dec1._045_ dec1._056_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_55_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_56_Right_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_71_593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_304 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0913_ _0359_ _0365_ _0356_ _0413_ _0441_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_0844_ _0360_ _0361_ _0367_ _0371_ _0372_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_0_43_348 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_359 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_11_256 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_65_Right_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_3_Left_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1327_ cal_lut\[30\] _0802_ _0804_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1258_ _0678_ _0697_ _0690_ _0767_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1189_ _0681_ _0703_ _0704_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_78_267 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_74_Right_74 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_93_259 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_356 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_326 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_49_Left_147 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_34_359 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_134 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_178 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_83_Right_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__0950__A1 _0376_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_58_Left_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1825__CLK net14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_85_674 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_92_Right_92 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_37_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_67_Left_165 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_clkbuf_1_1__f_io_in[0]_I clknet_0_io_in[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_101 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_348 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_381 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_52_189 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1194__A1 _0678_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_76_Left_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1112_ cal_lut\[5\] _0433_ _0357_ _0636_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1043_ _0566_ _0427_ _0567_ _0568_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_2
XPHY_EDGE_ROW_85_Left_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
Xtemp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[5\].vref temp1.dac.parallel_cells\[3\].vdac_batch.en_vref
+ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__invz_3
XTAP_TAPCELL_ROW_16_295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1421__A2 _0240_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_253 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0827_ _0355_ _0356_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
XPHY_EDGE_ROW_94_Left_192 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_43_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1488__A2 _0255_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1848__CLK clknet_1_1__leaf_io_in[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_82_655 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_164 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_229 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xseg1._43_ seg1._10_ seg1._15_ seg1.o_segments\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_22_329 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_381 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_7_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_395 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__0923__A1 _0365_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_318 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_329 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1100__A1 _0360_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_204 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_229 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_112 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_68 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_270 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_13_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1730_ _0082_ net16 cal_lut\[83\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1661_ _0013_ net17 cal_lut\[14\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1592_ _0314_ _0185_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input7_I io_in[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_43 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_98 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_31 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1026_ _0549_ _0395_ _0397_ _0550_ _0551_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_0_88_384 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_145 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1859_ _0211_ clknet_1_0__leaf_io_in[0] ctr\[12\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1670__CLK net16 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0905__A1 _0384_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1330__A1 cal_lut\[31\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_340 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_259 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_54_229 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_257 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xseg1._26_ dec1.o_dec\[3\] seg1._00_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_62_295 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1149__A1 _0670_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_181 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_93_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_18_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_45 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_218 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtemp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[3\].pupd temp1.dac.parallel_cells\[4\].vdac_batch.en_pupd
+ temp1.dac.parallel_cells\[4\].vdac_batch.npu_pd temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__invz_2
XFILLER_0_53_240 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_251 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1713_ _0065_ net11 cal_lut\[66\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1693__CLK net17 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_137 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1644_ _0783_ _0340_ _0211_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_1_0__f__0318_ clknet_0__0318_ clknet_1_0__leaf__0318_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_6_56 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1575_ _0308_ _0174_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1312__A1 cal_lut\[23\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1009_ _0376_ cal_lut\[117\] _0413_ _0406_ _0535_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XTAP_TAPCELL_ROW_24_338 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_91_324 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_153 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_381 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1443__I _0782_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xdec1._082_ dec1.i_bin\[4\] dec1._003_ dec1._022_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_82_302 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_26 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_346 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1360_ cal_lut\[50\] _0805_ _0218_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_37_45 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1291_ _0412_ _0790_ _0007_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_37_89 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1058__B1 _0433_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_376 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_21_319 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_temp1.dac.parallel_cells\[0\].vdac_batch._3__I temp1.dac.i_data\[0\] VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_251 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xtemp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[10\].vref temp1.dac.parallel_cells\[4\].vdac_batch.en_vref
+ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__invz_3
XFILLER_0_41_232 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_30 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1627_ _0345_ _0349_ _0330_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_68_4 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1558_ _0302_ _0163_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_21_Left_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1489_ _0274_ _0122_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__0887__A3 _0394_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_49_343 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_140 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_30_Left_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_76_184 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_154 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_52_488 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_165 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_32_265 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_416 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_129 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xdec1._065_ dec1.i_bin\[5\] dec1.i_bin\[4\] dec1._005_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_0860_ _0374_ _0375_ _0380_ _0387_ _0388_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_23_276 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1412_ _0243_ _0076_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1731__CLK net16 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1343_ _0475_ _0790_ _0038_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__0869__A3 _0355_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1274_ net3 _0780_ _0781_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_64_10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_32 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_66_569 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_140 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_316 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_73_154 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_176 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_210 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0989_ _0513_ _0414_ _0514_ _0515_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_73_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_95 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_96_213 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_96_257 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_162 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1037__A3 _0378_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_368 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1754__CLK net9 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_382 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0956__B _0433_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_235 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_268 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_302 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xdec1._117_ dec1._047_ dec1._040_ dec1._053_ dec1._055_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_71_594 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0912_ _0358_ _0391_ _0440_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_55_165 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_154 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0843_ _0368_ cal_lut\[133\] _0370_ _0371_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[13\].vref_I temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_65 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_76 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_279 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_268 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1326_ _0803_ _0029_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1257_ seg1.o_segments\[6\] _0691_ _0765_ _0694_ _0766_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_1188_ net6 _0682_ _0703_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_66_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1019__A3 _0373_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1777__CLK net8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_371 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_279 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_238 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_154 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_26 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_19 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1194__A2 _0684_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0941__A2 _0402_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1111_ _0588_ _0598_ _0607_ _0634_ _0635_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XTAP_TAPCELL_ROW_76_620 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1042_ _0390_ _0363_ cal_lut\[28\] _0384_ _0567_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_0_36 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_33 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_121 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_305 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_23 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_308 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_168 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_360 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_319 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0826_ dbg3\[0\] _0355_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_10_70 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0932__A2 _0383_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_41 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_74 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1309_ _0466_ _0790_ _0020_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_82_656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_187 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_74_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xseg1._42_ seg1._11_ seg1._14_ seg1._15_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_34_146 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__0923__A2 _0357_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_216 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_249 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_400 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_72_219 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1660_ _0012_ net14 cal_lut\[13\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1591_ cal_lut\[185\] _0294_ _0314_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1025_ cal_lut\[106\] _0550_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_48_227 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_54 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__0850__A1 _0362_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout10_I net13 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_357 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_71_241 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_91 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1858_ _0210_ clknet_1_0__leaf_io_in[0] ctr\[11\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_31_105 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1815__CLK net13 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1789_ _0141_ net14 cal_lut\[142\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_temp1.dac.parallel_cells\[1\].vdac_batch._4__A2 temp1.dac.i_data\[5\] VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0905__A2 _0413_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1330__A2 _0805_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0841__A1 _0365_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_219 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_93_718 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_127 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_18_303 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1085__A1 _0376_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_79 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1838__CLK net10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1712_ _0064_ net11 cal_lut\[65\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_53_263 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_274 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1643_ ctr\[12\] _0339_ _0340_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1574_ cal_lut\[174\] _0294_ _0308_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_6_68 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0899__A1 _0358_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1312__A2 _0780_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_472 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1076__A1 _0360_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1008_ cal_lut\[177\] _0534_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xtemp1.dac.parallel_cells\[2\].vdac_batch._8_ temp1.dac.parallel_cells\[2\].vdac_batch._0_
+ temp1.dac.parallel_cells\[2\].vdac_batch._1_ temp1.dac.parallel_cells\[2\].vdac_batch.en_vref
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_88_171 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_339 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_143 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_90 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1379__A2 _0802_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xtemp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[3\].vref temp1.dac.parallel_cells\[4\].vdac_batch.en_vref
+ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__invz_3
XANTENNA__1551__A2 _0289_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[0\].vref_I temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1303__A2 _0791_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1067__A1 _0390_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xtemp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[2\].pupd temp1.dac.parallel_cells\[2\].vdac_batch.en_pupd
+ temp1.dac.parallel_cells\[2\].vdac_batch.npu_pd temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__invz_2
XFILLER_0_79_171 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xdec1._081_ dec1._004_ dec1._020_ dec1._006_ dec1._021_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_50_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1542__A2 _0294_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_13 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1290_ _0779_ _0790_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_53_78 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1660__CLK net14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_196 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_124 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_263 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtemp1.dac.vdac_single._8_ temp1.dac.vdac_single._0_ temp1.dac.vdac_single._1_ temp1.dac.vdac_single.en_vref
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1230__A1 _0362_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_41_277 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1626_ _0783_ _0329_ _0204_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1557_ cal_lut\[163\] _0294_ _0302_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__1533__A2 _0289_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1488_ cal_lut\[122\] _0255_ _0274_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA_dec1._080__B dec1.i_bin\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_52_489 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_277 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1524__A2 _0289_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1683__CLK net11 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_119 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_152 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_303 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xdec1._064_ dec1.i_bin\[4\] dec1._003_ dec1.i_bin\[5\] dec1._004_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_55_358 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_200 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_380 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1411_ cal_lut\[76\] _0805_ _0243_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_48_12 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_23 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1342_ _0421_ _0790_ _0037_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1273_ _0779_ _0780_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_46_325 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_152 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_81 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_222 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0988_ _0359_ cal_lut\[93\] _0394_ _0514_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_14_277 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1506__A2 _0255_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1609_ _0362_ clknet_1_0__leaf__0318_ _0782_ _0322_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_69_417 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_152 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_347 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_426 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_214 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_314 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_100 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_208 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xdec1._116_ dec1._047_ dec1._053_ dec1._040_ dec1._054_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_43_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0911_ cal_lut\[169\] _0439_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_70_103 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_71_595 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0842_ _0362_ _0364_ _0369_ _0370_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_43_328 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_36_391 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_70_147 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_11 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1325_ cal_lut\[29\] _0802_ _0803_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_75_32 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_79_640 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1256_ _0670_ _0671_ _0691_ _0765_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[3\].vref_I temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1187_ _0346_ _0701_ _0687_ _0702_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_78_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_93_217 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_111 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_280 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_369 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_158 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_383 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0950__A3 _0422_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_90 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_203 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1721__CLK net9 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_147 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_136 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1110_ _0621_ _0628_ _0631_ _0633_ _0634_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XTAP_TAPCELL_ROW_76_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1041_ cal_lut\[112\] _0566_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_28_100 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_155 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_61_89 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_35 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_125 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_294 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_136 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0825_ _0354_ temp1.dac.i_enable VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_24_372 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_266 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_31 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1308_ _0409_ _0790_ _0019_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_29_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1239_ ctr\[4\] _0688_ _0750_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1645__A1 _0675_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1744__CLK net12 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_82_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_122 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_103 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_261 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xseg1._41_ dec1.o_dec\[2\] seg1._12_ seg1._13_ seg1._14_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA_temp1.dac.parallel_cells\[3\].vdac_batch._5__A1 temp1.dac.i_enable VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_342 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1100__A3 _0373_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_26 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_114 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_13_278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1590_ _0313_ _0184_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_56_23 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1767__CLK net12 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_78 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1024_ cal_lut\[190\] _0549_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_48_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1627__A1 _0345_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_99 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_325 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_63_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_81 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1857_ _0209_ clknet_1_0__leaf_io_in[0] ctr\[10\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_71_286 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_128 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1788_ _0140_ net14 cal_lut\[141\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_4_224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_301 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1231__B _0684_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0841__A2 _0356_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_412 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_294 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_220 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_242 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_10_259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_304 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1609__A1 _0362_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1085__A2 _0362_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_261 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1711_ _0063_ net9 cal_lut\[64\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1642_ ctr\[11\] _0353_ _0339_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_53_286 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_1_0__f__0316_ clknet_0__0316_ clknet_1_0__leaf__0316_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_21_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1573_ _0307_ _0173_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__0899__A2 _0365_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1076__A2 _0413_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1007_ _0531_ _0401_ _0440_ _0441_ _0532_ _0533_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai32_2
Xtemp1.dac.parallel_cells\[2\].vdac_batch._7_ temp1.dac.i_enable temp1.dac.parallel_cells\[2\].vdac_batch._0_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_88_183 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_111 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_348 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1277__I _0782_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_161 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1067__A2 _0363_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_183 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_194 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xdec1._080_ dec1.i_bin\[4\] dec1._003_ dec1.i_bin\[3\] dec1._020_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_12_28 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_381 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_309 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_286 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_68 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1805__CLK net16 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_367 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_73_348 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_136 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_242 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtemp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[2\].vref temp1.dac.parallel_cells\[2\].vdac_batch.en_vref
+ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__invz_3
Xtemp1.dac.vdac_single._7_ temp1.dac._0_ temp1.dac.vdac_single._0_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_5_169 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_234 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_267 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1625_ _0345_ _0349_ _0329_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1556_ _0301_ _0162_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1046__B _0433_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_31 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1487_ _0273_ _0121_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_11_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_37_410 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_345 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_134 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_156 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_253 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_381 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1288__A2 _0780_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1828__CLK net17 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_109 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xdec1._063_ dec1.i_bin\[5\] dec1.i_bin\[4\] dec1.i_bin\[6\] dec1._003_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XANTENNA__1460__A2 _0791_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0814__I ctr\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_348 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_156 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_23_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_329 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1410_ _0242_ _0075_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1341_ _0811_ _0036_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1272_ net1 _0779_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_64_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_164 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_359 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_88 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_73_178 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0987_ cal_lut\[9\] _0513_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_89_31 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1608_ ctr\[4\] clknet_1_1__leaf__0318_ _0321_ _0194_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_59_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1539_ _0295_ _0151_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_38_90 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1290__I _0779_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_57_516 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_65_560 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_164 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_40_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_362 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_384 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_226 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_0_Left_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1650__CLK net11 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_16_Right_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1130__A1 _0360_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xdec1._115_ dec1._026_ dec1._032_ dec1._053_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
X_0910_ _0435_ _0436_ _0437_ _0438_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_55_156 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1433__A2 _0240_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_71_596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0841_ _0365_ _0356_ _0369_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xtemp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[0\].pupd temp1.dac.parallel_cells\[3\].vdac_batch.en_pupd
+ temp1.dac.parallel_cells\[3\].vdac_batch.npu_pd temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__invz_2
XPHY_EDGE_ROW_25_Right_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1197__A1 _0357_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_384 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_259 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1324_ _0779_ _0802_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_79_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtemp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[9\].pupd temp1.dac.parallel_cells\[4\].vdac_batch.en_pupd
+ temp1.dac.parallel_cells\[4\].vdac_batch.npu_pd temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__invz_2
XPHY_EDGE_ROW_34_Right_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1255_ _0346_ ctr\[1\] _0708_ _0763_ _0764_ io_out[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_1186_ _0681_ _0686_ _0682_ _0701_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and3_2
XANTENNA__1121__A1 cal_lut\[54\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1121__B2 cal_lut\[48\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_229 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_304 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_123 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_101 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_292 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_381 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_43_Right_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_18_Left_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_6_297 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1673__CLK net15 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_dec1._086__B dec1.i_bin\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_281 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_292 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_52_Right_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_27_Left_125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__0871__B1 _0397_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_123 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1415__A2 _0240_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_61_Right_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_92_284 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_262 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_18_381 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_36_Left_134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_0_418 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_59 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_70_Right_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_45_Left_143 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_45_36 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_76_622 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1040_ _0376_ _0563_ _0422_ _0423_ _0564_ _0565_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_0_83_240 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_329 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_189 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_54_Left_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1696__CLK net17 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_0824_ dec1.i_ones ctr\[11\] ctr\[12\] _0353_ _0354_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_10_50 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_384 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0917__A1 _0358_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_65 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_temp1.dac.parallel_cells\[1\].vdac_batch.einvp_batch\[0\].vref_I temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_63_Left_161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1307_ _0795_ _0018_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1238_ _0675_ _0748_ _0690_ _0749_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1169_ _0683_ _0684_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_82_658 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_410 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_72_Left_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
Xseg1._40_ dec1.o_dec\[1\] dec1.o_dec\[0\] seg1._13_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__0908__A1 _0358_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1030__B1 _0408_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_376 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_57_218 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_137 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_148 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_310 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_181 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_118 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1021__B1 _0379_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1023_ _0544_ _0545_ _0546_ _0547_ _0548_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_48_229 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_78 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__0850__A3 _0365_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_temp1.dac.parallel_cells\[2\].vdac_batch._7__I temp1.dac.i_enable VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1856_ _0208_ clknet_1_0__leaf_io_in[0] ctr\[9\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_97_31 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_181 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1787_ _0139_ net14 cal_lut\[140\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_71_298 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_343 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1711__CLK net9 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_4_225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_2_Right_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1079__B1 _0386_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_207 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_1_1__f_net23 clknet_0_net23 clknet_1_1__leaf_net23 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_18_305 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_59 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_284 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_232 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1710_ _0062_ net8 cal_lut\[63\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1641_ _0783_ _0338_ _0210_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_6_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1572_ cal_lut\[173\] _0294_ _0307_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__1734__CLK net18 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0899__A3 _0356_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input5_I io_in[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_44 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_49_474 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_71 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1076__A3 _0406_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xtemp1.dac.parallel_cells\[2\].vdac_batch._6_ temp1.dac.parallel_cells\[2\].vdac_batch._2_
+ temp1.dac.parallel_cells\[2\].vdac_batch.en_pupd VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1006_ cal_lut\[15\] _0532_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_76_324 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_44_243 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1839_ _0191_ net12 cal_lut\[192\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_173 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1242__B _0684_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_346 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_187 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_23_330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_18 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_265 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_298 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1757__CLK net15 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[3\].vref_I temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_46_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1058__A3 _0582_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_346 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtemp1.dac.vdac_single._6_ temp1.dac.vdac_single._2_ temp1.dac.vdac_single.en_pupd
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_78_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1624_ _0349_ _0328_ _0783_ _0203_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1555_ cal_lut\[162\] _0294_ _0301_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_68_7 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_77 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_94_10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1486_ cal_lut\[121\] _0240_ _0273_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_94_65 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_94_98 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_80 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_368 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_349 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_265 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_298 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_276 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_213 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_181 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_dec1._108__I dec1.i_bin\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_68_580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xdec1._062_ dec1.i_ones dec1._001_ dec1._002_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_82_102 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_124 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_23_224 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_268 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0971__A2 _0452_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1340_ cal_lut\[36\] _0802_ _0811_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1271_ _0684_ _0777_ _0778_ io_out[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_78_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_198 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_308 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0986_ cal_lut\[183\] _0402_ _0403_ cal_lut\[51\] _0511_ _0512_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_1607_ _0363_ clknet_1_1__leaf__0318_ _0782_ _0321_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__0962__A2 _0401_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1538_ cal_lut\[151\] _0294_ _0295_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1469_ _0566_ _0791_ _0112_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_57_517 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_65_561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_349 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_284 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_262 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_374 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_88_686 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1130__A2 _0378_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xdec1._114_ dec1.i_tens dec1._046_ dec1._052_ dec1.o_dec\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_95_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_308 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_71_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0840_ _0358_ _0368_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_3_416 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_382 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_149 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1605__B _0782_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1323_ _0801_ _0028_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_38_8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1254_ temp1.dac.i_data\[5\] _0709_ _0684_ _0764_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1185_ _0688_ _0699_ _0700_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1121__A2 _0403_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_66 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0880__A1 _0359_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_221 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_243 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_265 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_0969_ _0363_ _0357_ _0496_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_27_393 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_61_138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_92 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1818__CLK net14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtemp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[0\].vref temp1.dac.parallel_cells\[3\].vdac_batch.en_vref
+ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__invz_3
XANTENNA__1360__A2 _0805_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_92 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1112__A2 _0433_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xtemp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[9\].vref temp1.dac.parallel_cells\[4\].vdac_batch.en_vref
+ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__invz_3
XFILLER_0_77_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_37_135 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_341 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0926__A2 _0452_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_16 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_193 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1351__A2 _0790_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_76_623 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_102 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_271 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0823_ _0343_ _0352_ _0353_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_24_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_84 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1342__A2 _0790_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1306_ cal_lut\[18\] _0780_ _0795_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1237_ _0744_ _0697_ _0745_ _0747_ _0748_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_1168_ _0681_ net6 _0682_ _0683_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__0853__A1 _0362_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1099_ _0368_ _0622_ _0378_ _0623_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_15_330 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_127 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0908__A2 _0362_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_160 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1790__CLK net12 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1581__A2 _0294_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_73_604 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0844__A1 _0360_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_208 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1572__A2 _0294_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1022_ cal_lut\[70\] _0383_ _0386_ cal_lut\[76\] _0547_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__1663__CLK net17 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_305 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_241 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0850__A4 _0356_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1855_ _0207_ clknet_1_0__leaf_io_in[0] ctr\[8\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_24_171 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1786_ _0138_ net12 cal_lut\[139\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_333 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1012__A1 _0508_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1563__A2 _0294_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_226 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_80 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_344 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1251__A1 _0345_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_417 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1003__A1 _0376_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1554__A2 _0289_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1306__A2 _0780_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1686__CLK net16 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_18_306 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0817__A1 _0346_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_26_350 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1085__A4 _0406_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_dec1._118__A1 dec1.i_tens VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_266 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1242__A1 temp1.dac.i_data\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1640_ _0733_ _0353_ _0338_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_41_417 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_288 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_91_Left_189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1571_ _0575_ _0289_ _0172_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__0899__A4 _0413_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1613__B _0782_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_92_710 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_49_475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1005_ cal_lut\[171\] _0531_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xtemp1.dac.parallel_cells\[2\].vdac_batch._5_ temp1.dac.i_enable temp1.dac.parallel_cells\[2\].vdac_batch._1_
+ temp1.dac.parallel_cells\[2\].vdac_batch._2_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_76_314 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_157 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_274 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1838_ _0190_ net10 cal_lut\[191\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1769_ _0121_ net10 cal_lut\[122\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_185 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_dec1._094__C dec1.i_bin\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_100 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1067__A4 _0384_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_23_331 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_306 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_222 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_303 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_166 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_328 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_26_233 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1215__A1 _0363_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1701__CLK net14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xtemp1.dac.vdac_single._5_ temp1.dac._0_ temp1.dac.vdac_single._1_ temp1.dac.vdac_single._2_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_26_299 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1623_ ctr\[4\] _0348_ _0328_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1851__CLK clknet_1_1__leaf_io_in[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1554_ _0629_ _0289_ _0161_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1485_ _0272_ _0120_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
.ends

