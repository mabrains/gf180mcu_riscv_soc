VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO peri_top
  CLASS BLOCK ;
  FOREIGN peri_top ;
  ORIGIN 0.000 0.000 ;
  SIZE 450.000 BY 300.000 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 19.940 15.380 26.140 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 119.940 15.380 126.140 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 219.940 15.380 226.140 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 319.940 15.380 326.140 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 419.940 15.380 426.140 282.540 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 69.940 15.380 76.140 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 169.940 15.380 176.140 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 269.940 15.380 276.140 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 369.940 15.380 376.140 282.540 ;
    END
  END VSS
  PIN mclk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 224.000 4.000 224.560 ;
    END
  END mclk
  PIN reg_ack
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 409.920 0.000 410.480 4.000 ;
    END
  END reg_ack
  PIN reg_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 100.800 0.000 101.360 4.000 ;
    END
  END reg_addr[0]
  PIN reg_addr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.898000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 56.000 0.000 56.560 4.000 ;
    END
  END reg_addr[10]
  PIN reg_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 96.320 0.000 96.880 4.000 ;
    END
  END reg_addr[1]
  PIN reg_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 91.840 0.000 92.400 4.000 ;
    END
  END reg_addr[2]
  PIN reg_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 87.360 0.000 87.920 4.000 ;
    END
  END reg_addr[3]
  PIN reg_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 82.880 0.000 83.440 4.000 ;
    END
  END reg_addr[4]
  PIN reg_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 78.400 0.000 78.960 4.000 ;
    END
  END reg_addr[5]
  PIN reg_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 73.920 0.000 74.480 4.000 ;
    END
  END reg_addr[6]
  PIN reg_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.898000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 69.440 0.000 70.000 4.000 ;
    END
  END reg_addr[7]
  PIN reg_addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.652000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 64.960 0.000 65.520 4.000 ;
    END
  END reg_addr[8]
  PIN reg_addr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.652000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 60.480 0.000 61.040 4.000 ;
    END
  END reg_addr[9]
  PIN reg_be[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 118.720 0.000 119.280 4.000 ;
    END
  END reg_be[0]
  PIN reg_be[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 114.240 0.000 114.800 4.000 ;
    END
  END reg_be[1]
  PIN reg_be[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 109.760 0.000 110.320 4.000 ;
    END
  END reg_be[2]
  PIN reg_be[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 105.280 0.000 105.840 4.000 ;
    END
  END reg_be[3]
  PIN reg_cs
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 47.040 0.000 47.600 4.000 ;
    END
  END reg_cs
  PIN reg_rdata[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 405.440 0.000 406.000 4.000 ;
    END
  END reg_rdata[0]
  PIN reg_rdata[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 360.640 0.000 361.200 4.000 ;
    END
  END reg_rdata[10]
  PIN reg_rdata[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 356.160 0.000 356.720 4.000 ;
    END
  END reg_rdata[11]
  PIN reg_rdata[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 351.680 0.000 352.240 4.000 ;
    END
  END reg_rdata[12]
  PIN reg_rdata[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 347.200 0.000 347.760 4.000 ;
    END
  END reg_rdata[13]
  PIN reg_rdata[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 342.720 0.000 343.280 4.000 ;
    END
  END reg_rdata[14]
  PIN reg_rdata[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 338.240 0.000 338.800 4.000 ;
    END
  END reg_rdata[15]
  PIN reg_rdata[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 333.760 0.000 334.320 4.000 ;
    END
  END reg_rdata[16]
  PIN reg_rdata[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 329.280 0.000 329.840 4.000 ;
    END
  END reg_rdata[17]
  PIN reg_rdata[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 324.800 0.000 325.360 4.000 ;
    END
  END reg_rdata[18]
  PIN reg_rdata[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 320.320 0.000 320.880 4.000 ;
    END
  END reg_rdata[19]
  PIN reg_rdata[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 400.960 0.000 401.520 4.000 ;
    END
  END reg_rdata[1]
  PIN reg_rdata[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 315.840 0.000 316.400 4.000 ;
    END
  END reg_rdata[20]
  PIN reg_rdata[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 311.360 0.000 311.920 4.000 ;
    END
  END reg_rdata[21]
  PIN reg_rdata[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 306.880 0.000 307.440 4.000 ;
    END
  END reg_rdata[22]
  PIN reg_rdata[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 302.400 0.000 302.960 4.000 ;
    END
  END reg_rdata[23]
  PIN reg_rdata[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 297.920 0.000 298.480 4.000 ;
    END
  END reg_rdata[24]
  PIN reg_rdata[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 293.440 0.000 294.000 4.000 ;
    END
  END reg_rdata[25]
  PIN reg_rdata[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 288.960 0.000 289.520 4.000 ;
    END
  END reg_rdata[26]
  PIN reg_rdata[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 284.480 0.000 285.040 4.000 ;
    END
  END reg_rdata[27]
  PIN reg_rdata[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 280.000 0.000 280.560 4.000 ;
    END
  END reg_rdata[28]
  PIN reg_rdata[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 275.520 0.000 276.080 4.000 ;
    END
  END reg_rdata[29]
  PIN reg_rdata[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 396.480 0.000 397.040 4.000 ;
    END
  END reg_rdata[2]
  PIN reg_rdata[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 271.040 0.000 271.600 4.000 ;
    END
  END reg_rdata[30]
  PIN reg_rdata[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 266.560 0.000 267.120 4.000 ;
    END
  END reg_rdata[31]
  PIN reg_rdata[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 392.000 0.000 392.560 4.000 ;
    END
  END reg_rdata[3]
  PIN reg_rdata[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 387.520 0.000 388.080 4.000 ;
    END
  END reg_rdata[4]
  PIN reg_rdata[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 383.040 0.000 383.600 4.000 ;
    END
  END reg_rdata[5]
  PIN reg_rdata[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 378.560 0.000 379.120 4.000 ;
    END
  END reg_rdata[6]
  PIN reg_rdata[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 374.080 0.000 374.640 4.000 ;
    END
  END reg_rdata[7]
  PIN reg_rdata[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 369.600 0.000 370.160 4.000 ;
    END
  END reg_rdata[8]
  PIN reg_rdata[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 365.120 0.000 365.680 4.000 ;
    END
  END reg_rdata[9]
  PIN reg_wdata[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 262.080 0.000 262.640 4.000 ;
    END
  END reg_wdata[0]
  PIN reg_wdata[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 217.280 0.000 217.840 4.000 ;
    END
  END reg_wdata[10]
  PIN reg_wdata[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 212.800 0.000 213.360 4.000 ;
    END
  END reg_wdata[11]
  PIN reg_wdata[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 208.320 0.000 208.880 4.000 ;
    END
  END reg_wdata[12]
  PIN reg_wdata[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 203.840 0.000 204.400 4.000 ;
    END
  END reg_wdata[13]
  PIN reg_wdata[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 199.360 0.000 199.920 4.000 ;
    END
  END reg_wdata[14]
  PIN reg_wdata[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 194.880 0.000 195.440 4.000 ;
    END
  END reg_wdata[15]
  PIN reg_wdata[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 190.400 0.000 190.960 4.000 ;
    END
  END reg_wdata[16]
  PIN reg_wdata[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 185.920 0.000 186.480 4.000 ;
    END
  END reg_wdata[17]
  PIN reg_wdata[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 181.440 0.000 182.000 4.000 ;
    END
  END reg_wdata[18]
  PIN reg_wdata[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 176.960 0.000 177.520 4.000 ;
    END
  END reg_wdata[19]
  PIN reg_wdata[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 257.600 0.000 258.160 4.000 ;
    END
  END reg_wdata[1]
  PIN reg_wdata[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 172.480 0.000 173.040 4.000 ;
    END
  END reg_wdata[20]
  PIN reg_wdata[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 168.000 0.000 168.560 4.000 ;
    END
  END reg_wdata[21]
  PIN reg_wdata[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 163.520 0.000 164.080 4.000 ;
    END
  END reg_wdata[22]
  PIN reg_wdata[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 159.040 0.000 159.600 4.000 ;
    END
  END reg_wdata[23]
  PIN reg_wdata[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 154.560 0.000 155.120 4.000 ;
    END
  END reg_wdata[24]
  PIN reg_wdata[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 150.080 0.000 150.640 4.000 ;
    END
  END reg_wdata[25]
  PIN reg_wdata[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 145.600 0.000 146.160 4.000 ;
    END
  END reg_wdata[26]
  PIN reg_wdata[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 141.120 0.000 141.680 4.000 ;
    END
  END reg_wdata[27]
  PIN reg_wdata[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 136.640 0.000 137.200 4.000 ;
    END
  END reg_wdata[28]
  PIN reg_wdata[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 132.160 0.000 132.720 4.000 ;
    END
  END reg_wdata[29]
  PIN reg_wdata[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 253.120 0.000 253.680 4.000 ;
    END
  END reg_wdata[2]
  PIN reg_wdata[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 127.680 0.000 128.240 4.000 ;
    END
  END reg_wdata[30]
  PIN reg_wdata[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 123.200 0.000 123.760 4.000 ;
    END
  END reg_wdata[31]
  PIN reg_wdata[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 248.640 0.000 249.200 4.000 ;
    END
  END reg_wdata[3]
  PIN reg_wdata[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 244.160 0.000 244.720 4.000 ;
    END
  END reg_wdata[4]
  PIN reg_wdata[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 239.680 0.000 240.240 4.000 ;
    END
  END reg_wdata[5]
  PIN reg_wdata[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 235.200 0.000 235.760 4.000 ;
    END
  END reg_wdata[6]
  PIN reg_wdata[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 230.720 0.000 231.280 4.000 ;
    END
  END reg_wdata[7]
  PIN reg_wdata[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 226.240 0.000 226.800 4.000 ;
    END
  END reg_wdata[8]
  PIN reg_wdata[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 221.760 0.000 222.320 4.000 ;
    END
  END reg_wdata[9]
  PIN reg_wr
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 51.520 0.000 52.080 4.000 ;
    END
  END reg_wr
  PIN rtc_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 38.080 0.000 38.640 4.000 ;
    END
  END rtc_clk
  PIN rtc_intr
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 42.560 0.000 43.120 4.000 ;
    END
  END rtc_intr
  PIN s_reset_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.498000 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 73.920 4.000 74.480 ;
    END
  END s_reset_n
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 442.960 282.540 ;
      LAYER Metal2 ;
        RECT 9.100 4.300 441.700 282.430 ;
        RECT 9.100 3.500 37.780 4.300 ;
        RECT 38.940 3.500 42.260 4.300 ;
        RECT 43.420 3.500 46.740 4.300 ;
        RECT 47.900 3.500 51.220 4.300 ;
        RECT 52.380 3.500 55.700 4.300 ;
        RECT 56.860 3.500 60.180 4.300 ;
        RECT 61.340 3.500 64.660 4.300 ;
        RECT 65.820 3.500 69.140 4.300 ;
        RECT 70.300 3.500 73.620 4.300 ;
        RECT 74.780 3.500 78.100 4.300 ;
        RECT 79.260 3.500 82.580 4.300 ;
        RECT 83.740 3.500 87.060 4.300 ;
        RECT 88.220 3.500 91.540 4.300 ;
        RECT 92.700 3.500 96.020 4.300 ;
        RECT 97.180 3.500 100.500 4.300 ;
        RECT 101.660 3.500 104.980 4.300 ;
        RECT 106.140 3.500 109.460 4.300 ;
        RECT 110.620 3.500 113.940 4.300 ;
        RECT 115.100 3.500 118.420 4.300 ;
        RECT 119.580 3.500 122.900 4.300 ;
        RECT 124.060 3.500 127.380 4.300 ;
        RECT 128.540 3.500 131.860 4.300 ;
        RECT 133.020 3.500 136.340 4.300 ;
        RECT 137.500 3.500 140.820 4.300 ;
        RECT 141.980 3.500 145.300 4.300 ;
        RECT 146.460 3.500 149.780 4.300 ;
        RECT 150.940 3.500 154.260 4.300 ;
        RECT 155.420 3.500 158.740 4.300 ;
        RECT 159.900 3.500 163.220 4.300 ;
        RECT 164.380 3.500 167.700 4.300 ;
        RECT 168.860 3.500 172.180 4.300 ;
        RECT 173.340 3.500 176.660 4.300 ;
        RECT 177.820 3.500 181.140 4.300 ;
        RECT 182.300 3.500 185.620 4.300 ;
        RECT 186.780 3.500 190.100 4.300 ;
        RECT 191.260 3.500 194.580 4.300 ;
        RECT 195.740 3.500 199.060 4.300 ;
        RECT 200.220 3.500 203.540 4.300 ;
        RECT 204.700 3.500 208.020 4.300 ;
        RECT 209.180 3.500 212.500 4.300 ;
        RECT 213.660 3.500 216.980 4.300 ;
        RECT 218.140 3.500 221.460 4.300 ;
        RECT 222.620 3.500 225.940 4.300 ;
        RECT 227.100 3.500 230.420 4.300 ;
        RECT 231.580 3.500 234.900 4.300 ;
        RECT 236.060 3.500 239.380 4.300 ;
        RECT 240.540 3.500 243.860 4.300 ;
        RECT 245.020 3.500 248.340 4.300 ;
        RECT 249.500 3.500 252.820 4.300 ;
        RECT 253.980 3.500 257.300 4.300 ;
        RECT 258.460 3.500 261.780 4.300 ;
        RECT 262.940 3.500 266.260 4.300 ;
        RECT 267.420 3.500 270.740 4.300 ;
        RECT 271.900 3.500 275.220 4.300 ;
        RECT 276.380 3.500 279.700 4.300 ;
        RECT 280.860 3.500 284.180 4.300 ;
        RECT 285.340 3.500 288.660 4.300 ;
        RECT 289.820 3.500 293.140 4.300 ;
        RECT 294.300 3.500 297.620 4.300 ;
        RECT 298.780 3.500 302.100 4.300 ;
        RECT 303.260 3.500 306.580 4.300 ;
        RECT 307.740 3.500 311.060 4.300 ;
        RECT 312.220 3.500 315.540 4.300 ;
        RECT 316.700 3.500 320.020 4.300 ;
        RECT 321.180 3.500 324.500 4.300 ;
        RECT 325.660 3.500 328.980 4.300 ;
        RECT 330.140 3.500 333.460 4.300 ;
        RECT 334.620 3.500 337.940 4.300 ;
        RECT 339.100 3.500 342.420 4.300 ;
        RECT 343.580 3.500 346.900 4.300 ;
        RECT 348.060 3.500 351.380 4.300 ;
        RECT 352.540 3.500 355.860 4.300 ;
        RECT 357.020 3.500 360.340 4.300 ;
        RECT 361.500 3.500 364.820 4.300 ;
        RECT 365.980 3.500 369.300 4.300 ;
        RECT 370.460 3.500 373.780 4.300 ;
        RECT 374.940 3.500 378.260 4.300 ;
        RECT 379.420 3.500 382.740 4.300 ;
        RECT 383.900 3.500 387.220 4.300 ;
        RECT 388.380 3.500 391.700 4.300 ;
        RECT 392.860 3.500 396.180 4.300 ;
        RECT 397.340 3.500 400.660 4.300 ;
        RECT 401.820 3.500 405.140 4.300 ;
        RECT 406.300 3.500 409.620 4.300 ;
        RECT 410.780 3.500 441.700 4.300 ;
      LAYER Metal3 ;
        RECT 4.000 224.860 441.750 282.380 ;
        RECT 4.300 223.700 441.750 224.860 ;
        RECT 4.000 74.780 441.750 223.700 ;
        RECT 4.300 73.620 441.750 74.780 ;
        RECT 4.000 14.700 441.750 73.620 ;
      LAYER Metal4 ;
        RECT 26.460 16.890 69.640 269.270 ;
        RECT 76.440 16.890 119.640 269.270 ;
        RECT 126.440 16.890 169.640 269.270 ;
        RECT 176.440 16.890 219.640 269.270 ;
        RECT 226.440 16.890 269.640 269.270 ;
        RECT 276.440 16.890 319.640 269.270 ;
        RECT 326.440 16.890 369.640 269.270 ;
        RECT 376.440 16.890 419.640 269.270 ;
        RECT 426.440 16.890 428.260 269.270 ;
  END
END peri_top
END LIBRARY

