magic
tech gf180mcuD
magscale 1 5
timestamp 1700952138
<< nwell >>
rect 629 172656 254339 173088
rect 629 171872 254339 172304
rect 629 171088 254339 171520
rect 629 170304 254339 170736
rect 629 169520 254339 169952
rect 629 168736 254339 169168
rect 629 167952 254339 168384
rect 629 167168 254339 167600
rect 629 166384 254339 166816
rect 629 165600 254339 166032
rect 629 164816 254339 165248
rect 629 164032 254339 164464
rect 629 163248 254339 163680
rect 629 162464 254339 162896
rect 629 161680 254339 162112
rect 629 160896 254339 161328
rect 629 160112 254339 160544
rect 629 159328 254339 159760
rect 629 158544 254339 158976
rect 629 157760 254339 158192
rect 629 156976 254339 157408
rect 629 156192 254339 156624
rect 629 155408 254339 155840
rect 629 154624 254339 155056
rect 629 153840 254339 154272
rect 629 153056 254339 153488
rect 629 152272 254339 152704
rect 629 151488 254339 151920
rect 629 150704 254339 151136
rect 629 149920 254339 150352
rect 629 149136 254339 149568
rect 629 148352 254339 148784
rect 629 147568 254339 148000
rect 629 146784 254339 147216
rect 629 146000 254339 146432
rect 629 145216 254339 145648
rect 629 144432 254339 144864
rect 629 143648 254339 144080
rect 629 142864 254339 143296
rect 629 142080 254339 142512
rect 629 141296 254339 141728
rect 629 140512 254339 140944
rect 629 139728 254339 140160
rect 629 138944 254339 139376
rect 629 138160 254339 138592
rect 629 137376 254339 137808
rect 629 136592 254339 137024
rect 629 135808 254339 136240
rect 629 135024 254339 135456
rect 629 134240 254339 134672
rect 629 133456 254339 133888
rect 629 132672 254339 133104
rect 629 131888 254339 132320
rect 629 131104 254339 131536
rect 629 130320 254339 130752
rect 629 129536 254339 129968
rect 629 128752 254339 129184
rect 629 127968 254339 128400
rect 629 127184 254339 127616
rect 629 126400 254339 126832
rect 629 125616 254339 126048
rect 629 124832 254339 125264
rect 629 124048 254339 124480
rect 629 123264 254339 123696
rect 629 122480 254339 122912
rect 629 121696 254339 122128
rect 629 120912 254339 121344
rect 629 120128 254339 120560
rect 629 119344 254339 119776
rect 629 118560 254339 118992
rect 629 117776 254339 118208
rect 629 116992 254339 117424
rect 629 116208 254339 116640
rect 629 115424 254339 115856
rect 629 114640 254339 115072
rect 629 113856 254339 114288
rect 629 113072 254339 113504
rect 629 112288 254339 112720
rect 629 111504 254339 111936
rect 629 110720 254339 111152
rect 629 109936 254339 110368
rect 629 109152 254339 109584
rect 629 108368 254339 108800
rect 629 107584 254339 108016
rect 629 106800 254339 107232
rect 629 106016 254339 106448
rect 629 105232 254339 105664
rect 629 104448 254339 104880
rect 629 103664 254339 104096
rect 629 102880 254339 103312
rect 629 102096 254339 102528
rect 629 101312 254339 101744
rect 629 100528 254339 100960
rect 629 99744 254339 100176
rect 629 98960 254339 99392
rect 629 98176 254339 98608
rect 629 97392 254339 97824
rect 629 96608 254339 97040
rect 629 95824 254339 96256
rect 629 95040 254339 95472
rect 629 94256 254339 94688
rect 629 93472 254339 93904
rect 629 92688 254339 93120
rect 629 91904 254339 92336
rect 629 91120 254339 91552
rect 629 90336 254339 90768
rect 629 89552 254339 89984
rect 629 88768 254339 89200
rect 629 87984 254339 88416
rect 629 87200 254339 87632
rect 629 86416 254339 86848
rect 629 85632 254339 86064
rect 629 84848 254339 85280
rect 629 84064 254339 84496
rect 629 83280 254339 83712
rect 629 82496 254339 82928
rect 629 81712 254339 82144
rect 629 80928 254339 81360
rect 629 80144 254339 80576
rect 629 79360 254339 79792
rect 629 78576 254339 79008
rect 629 77792 254339 78224
rect 629 77008 254339 77440
rect 629 76224 254339 76656
rect 629 75440 254339 75872
rect 629 74656 254339 75088
rect 629 73872 254339 74304
rect 629 73088 254339 73520
rect 629 72304 254339 72736
rect 629 71520 254339 71952
rect 629 70736 254339 71168
rect 629 69952 254339 70384
rect 629 69168 254339 69600
rect 629 68384 254339 68816
rect 629 67600 254339 68032
rect 629 66816 254339 67248
rect 629 66032 254339 66464
rect 629 65248 254339 65680
rect 629 64464 254339 64896
rect 629 63680 254339 64112
rect 629 62896 254339 63328
rect 629 62112 254339 62544
rect 629 61328 254339 61760
rect 629 60544 254339 60976
rect 629 59760 254339 60192
rect 629 58976 254339 59408
rect 629 58192 254339 58624
rect 629 57408 254339 57840
rect 629 56624 254339 57056
rect 629 55840 254339 56272
rect 629 55056 254339 55488
rect 629 54272 254339 54704
rect 629 53488 254339 53920
rect 629 52704 254339 53136
rect 629 51920 254339 52352
rect 629 51136 254339 51568
rect 629 50352 254339 50784
rect 629 49568 254339 50000
rect 629 48784 254339 49216
rect 629 48000 254339 48432
rect 629 47216 254339 47648
rect 629 46432 254339 46864
rect 629 45648 254339 46080
rect 629 44864 254339 45296
rect 629 44080 254339 44512
rect 629 43296 254339 43728
rect 629 42512 254339 42944
rect 629 41728 254339 42160
rect 629 40944 254339 41376
rect 629 40160 254339 40592
rect 629 39376 254339 39808
rect 629 38592 254339 39024
rect 629 37808 254339 38240
rect 629 37024 254339 37456
rect 629 36240 254339 36672
rect 629 35456 254339 35888
rect 629 34672 254339 35104
rect 629 33888 254339 34320
rect 629 33104 254339 33536
rect 629 32320 254339 32752
rect 629 31536 254339 31968
rect 629 30752 254339 31184
rect 629 29968 254339 30400
rect 629 29184 254339 29616
rect 629 28400 254339 28832
rect 629 27616 254339 28048
rect 629 26832 254339 27264
rect 629 26048 254339 26480
rect 629 25264 254339 25696
rect 629 24480 254339 24912
rect 629 23696 254339 24128
rect 629 22912 254339 23344
rect 629 22128 254339 22560
rect 629 21344 254339 21776
rect 629 20560 254339 20992
rect 629 19776 254339 20208
rect 629 18992 254339 19424
rect 629 18208 254339 18640
rect 629 17424 254339 17856
rect 629 16640 254339 17072
rect 629 15856 254339 16288
rect 629 15072 254339 15504
rect 629 14288 254339 14720
rect 629 13504 254339 13936
rect 629 12720 254339 13152
rect 629 11936 254339 12368
rect 629 11152 254339 11584
rect 629 10368 254339 10800
rect 629 9584 254339 10016
rect 629 8800 254339 9232
rect 629 8016 254339 8448
rect 629 7232 254339 7664
rect 629 6448 254339 6880
rect 629 5664 254339 6096
rect 629 4880 254339 5312
rect 629 4096 254339 4528
rect 629 3312 254339 3744
rect 629 2528 254339 2960
rect 629 1744 254339 2176
<< pwell >>
rect 629 173088 254339 173307
rect 629 172304 254339 172656
rect 629 171520 254339 171872
rect 629 170736 254339 171088
rect 629 169952 254339 170304
rect 629 169168 254339 169520
rect 629 168384 254339 168736
rect 629 167600 254339 167952
rect 629 166816 254339 167168
rect 629 166032 254339 166384
rect 629 165248 254339 165600
rect 629 164464 254339 164816
rect 629 163680 254339 164032
rect 629 162896 254339 163248
rect 629 162112 254339 162464
rect 629 161328 254339 161680
rect 629 160544 254339 160896
rect 629 159760 254339 160112
rect 629 158976 254339 159328
rect 629 158192 254339 158544
rect 629 157408 254339 157760
rect 629 156624 254339 156976
rect 629 155840 254339 156192
rect 629 155056 254339 155408
rect 629 154272 254339 154624
rect 629 153488 254339 153840
rect 629 152704 254339 153056
rect 629 151920 254339 152272
rect 629 151136 254339 151488
rect 629 150352 254339 150704
rect 629 149568 254339 149920
rect 629 148784 254339 149136
rect 629 148000 254339 148352
rect 629 147216 254339 147568
rect 629 146432 254339 146784
rect 629 145648 254339 146000
rect 629 144864 254339 145216
rect 629 144080 254339 144432
rect 629 143296 254339 143648
rect 629 142512 254339 142864
rect 629 141728 254339 142080
rect 629 140944 254339 141296
rect 629 140160 254339 140512
rect 629 139376 254339 139728
rect 629 138592 254339 138944
rect 629 137808 254339 138160
rect 629 137024 254339 137376
rect 629 136240 254339 136592
rect 629 135456 254339 135808
rect 629 134672 254339 135024
rect 629 133888 254339 134240
rect 629 133104 254339 133456
rect 629 132320 254339 132672
rect 629 131536 254339 131888
rect 629 130752 254339 131104
rect 629 129968 254339 130320
rect 629 129184 254339 129536
rect 629 128400 254339 128752
rect 629 127616 254339 127968
rect 629 126832 254339 127184
rect 629 126048 254339 126400
rect 629 125264 254339 125616
rect 629 124480 254339 124832
rect 629 123696 254339 124048
rect 629 122912 254339 123264
rect 629 122128 254339 122480
rect 629 121344 254339 121696
rect 629 120560 254339 120912
rect 629 119776 254339 120128
rect 629 118992 254339 119344
rect 629 118208 254339 118560
rect 629 117424 254339 117776
rect 629 116640 254339 116992
rect 629 115856 254339 116208
rect 629 115072 254339 115424
rect 629 114288 254339 114640
rect 629 113504 254339 113856
rect 629 112720 254339 113072
rect 629 111936 254339 112288
rect 629 111152 254339 111504
rect 629 110368 254339 110720
rect 629 109584 254339 109936
rect 629 108800 254339 109152
rect 629 108016 254339 108368
rect 629 107232 254339 107584
rect 629 106448 254339 106800
rect 629 105664 254339 106016
rect 629 104880 254339 105232
rect 629 104096 254339 104448
rect 629 103312 254339 103664
rect 629 102528 254339 102880
rect 629 101744 254339 102096
rect 629 100960 254339 101312
rect 629 100176 254339 100528
rect 629 99392 254339 99744
rect 629 98608 254339 98960
rect 629 97824 254339 98176
rect 629 97040 254339 97392
rect 629 96256 254339 96608
rect 629 95472 254339 95824
rect 629 94688 254339 95040
rect 629 93904 254339 94256
rect 629 93120 254339 93472
rect 629 92336 254339 92688
rect 629 91552 254339 91904
rect 629 90768 254339 91120
rect 629 89984 254339 90336
rect 629 89200 254339 89552
rect 629 88416 254339 88768
rect 629 87632 254339 87984
rect 629 86848 254339 87200
rect 629 86064 254339 86416
rect 629 85280 254339 85632
rect 629 84496 254339 84848
rect 629 83712 254339 84064
rect 629 82928 254339 83280
rect 629 82144 254339 82496
rect 629 81360 254339 81712
rect 629 80576 254339 80928
rect 629 79792 254339 80144
rect 629 79008 254339 79360
rect 629 78224 254339 78576
rect 629 77440 254339 77792
rect 629 76656 254339 77008
rect 629 75872 254339 76224
rect 629 75088 254339 75440
rect 629 74304 254339 74656
rect 629 73520 254339 73872
rect 629 72736 254339 73088
rect 629 71952 254339 72304
rect 629 71168 254339 71520
rect 629 70384 254339 70736
rect 629 69600 254339 69952
rect 629 68816 254339 69168
rect 629 68032 254339 68384
rect 629 67248 254339 67600
rect 629 66464 254339 66816
rect 629 65680 254339 66032
rect 629 64896 254339 65248
rect 629 64112 254339 64464
rect 629 63328 254339 63680
rect 629 62544 254339 62896
rect 629 61760 254339 62112
rect 629 60976 254339 61328
rect 629 60192 254339 60544
rect 629 59408 254339 59760
rect 629 58624 254339 58976
rect 629 57840 254339 58192
rect 629 57056 254339 57408
rect 629 56272 254339 56624
rect 629 55488 254339 55840
rect 629 54704 254339 55056
rect 629 53920 254339 54272
rect 629 53136 254339 53488
rect 629 52352 254339 52704
rect 629 51568 254339 51920
rect 629 50784 254339 51136
rect 629 50000 254339 50352
rect 629 49216 254339 49568
rect 629 48432 254339 48784
rect 629 47648 254339 48000
rect 629 46864 254339 47216
rect 629 46080 254339 46432
rect 629 45296 254339 45648
rect 629 44512 254339 44864
rect 629 43728 254339 44080
rect 629 42944 254339 43296
rect 629 42160 254339 42512
rect 629 41376 254339 41728
rect 629 40592 254339 40944
rect 629 39808 254339 40160
rect 629 39024 254339 39376
rect 629 38240 254339 38592
rect 629 37456 254339 37808
rect 629 36672 254339 37024
rect 629 35888 254339 36240
rect 629 35104 254339 35456
rect 629 34320 254339 34672
rect 629 33536 254339 33888
rect 629 32752 254339 33104
rect 629 31968 254339 32320
rect 629 31184 254339 31536
rect 629 30400 254339 30752
rect 629 29616 254339 29968
rect 629 28832 254339 29184
rect 629 28048 254339 28400
rect 629 27264 254339 27616
rect 629 26480 254339 26832
rect 629 25696 254339 26048
rect 629 24912 254339 25264
rect 629 24128 254339 24480
rect 629 23344 254339 23696
rect 629 22560 254339 22912
rect 629 21776 254339 22128
rect 629 20992 254339 21344
rect 629 20208 254339 20560
rect 629 19424 254339 19776
rect 629 18640 254339 18992
rect 629 17856 254339 18208
rect 629 17072 254339 17424
rect 629 16288 254339 16640
rect 629 15504 254339 15856
rect 629 14720 254339 15072
rect 629 13936 254339 14288
rect 629 13152 254339 13504
rect 629 12368 254339 12720
rect 629 11584 254339 11936
rect 629 10800 254339 11152
rect 629 10016 254339 10368
rect 629 9232 254339 9584
rect 629 8448 254339 8800
rect 629 7664 254339 8016
rect 629 6880 254339 7232
rect 629 6096 254339 6448
rect 629 5312 254339 5664
rect 629 4528 254339 4880
rect 629 3744 254339 4096
rect 629 2960 254339 3312
rect 629 2176 254339 2528
rect 629 1525 254339 1744
<< obsm1 >>
rect 672 1538 254296 173294
<< metal2 >>
rect 127344 174600 127400 175000
rect 127008 0 127064 400
rect 127344 0 127400 400
<< obsm2 >>
rect 2004 174570 127314 174600
rect 127430 174570 252604 174600
rect 2004 430 252604 174570
rect 2004 400 126978 430
rect 127094 400 127314 430
rect 127430 400 252604 430
<< obsm3 >>
rect 1999 462 252609 173278
<< metal4 >>
rect 1994 1538 2614 173294
rect 6994 1538 7614 173294
rect 11994 1538 12614 173294
rect 16994 1538 17614 173294
rect 21994 1538 22614 173294
rect 26994 1538 27614 173294
rect 31994 1538 32614 173294
rect 36994 1538 37614 173294
rect 41994 1538 42614 173294
rect 46994 1538 47614 173294
rect 51994 1538 52614 173294
rect 56994 1538 57614 173294
rect 61994 1538 62614 173294
rect 66994 1538 67614 173294
rect 71994 1538 72614 173294
rect 76994 1538 77614 173294
rect 81994 1538 82614 173294
rect 86994 1538 87614 173294
rect 91994 1538 92614 173294
rect 96994 1538 97614 173294
rect 101994 1538 102614 173294
rect 106994 1538 107614 173294
rect 111994 1538 112614 173294
rect 116994 1538 117614 173294
rect 121994 1538 122614 173294
rect 126994 1538 127614 173294
rect 131994 1538 132614 173294
rect 136994 1538 137614 173294
rect 141994 1538 142614 173294
rect 146994 1538 147614 173294
rect 151994 1538 152614 173294
rect 156994 1538 157614 173294
rect 161994 1538 162614 173294
rect 166994 1538 167614 173294
rect 171994 1538 172614 173294
rect 176994 1538 177614 173294
rect 181994 1538 182614 173294
rect 186994 1538 187614 173294
rect 191994 1538 192614 173294
rect 196994 1538 197614 173294
rect 201994 1538 202614 173294
rect 206994 1538 207614 173294
rect 211994 1538 212614 173294
rect 216994 1538 217614 173294
rect 221994 1538 222614 173294
rect 226994 1538 227614 173294
rect 231994 1538 232614 173294
rect 236994 1538 237614 173294
rect 241994 1538 242614 173294
rect 246994 1538 247614 173294
rect 251994 1538 252614 173294
<< labels >>
rlabel metal2 s 127344 0 127400 400 6 in1
port 1 nsew signal input
rlabel metal2 s 127008 0 127064 400 6 in2
port 2 nsew signal input
rlabel metal2 s 127344 174600 127400 175000 6 out
port 3 nsew signal output
rlabel metal4 s 1994 1538 2614 173294 6 vdd
port 4 nsew power bidirectional
rlabel metal4 s 11994 1538 12614 173294 6 vdd
port 4 nsew power bidirectional
rlabel metal4 s 21994 1538 22614 173294 6 vdd
port 4 nsew power bidirectional
rlabel metal4 s 31994 1538 32614 173294 6 vdd
port 4 nsew power bidirectional
rlabel metal4 s 41994 1538 42614 173294 6 vdd
port 4 nsew power bidirectional
rlabel metal4 s 51994 1538 52614 173294 6 vdd
port 4 nsew power bidirectional
rlabel metal4 s 61994 1538 62614 173294 6 vdd
port 4 nsew power bidirectional
rlabel metal4 s 71994 1538 72614 173294 6 vdd
port 4 nsew power bidirectional
rlabel metal4 s 81994 1538 82614 173294 6 vdd
port 4 nsew power bidirectional
rlabel metal4 s 91994 1538 92614 173294 6 vdd
port 4 nsew power bidirectional
rlabel metal4 s 101994 1538 102614 173294 6 vdd
port 4 nsew power bidirectional
rlabel metal4 s 111994 1538 112614 173294 6 vdd
port 4 nsew power bidirectional
rlabel metal4 s 121994 1538 122614 173294 6 vdd
port 4 nsew power bidirectional
rlabel metal4 s 131994 1538 132614 173294 6 vdd
port 4 nsew power bidirectional
rlabel metal4 s 141994 1538 142614 173294 6 vdd
port 4 nsew power bidirectional
rlabel metal4 s 151994 1538 152614 173294 6 vdd
port 4 nsew power bidirectional
rlabel metal4 s 161994 1538 162614 173294 6 vdd
port 4 nsew power bidirectional
rlabel metal4 s 171994 1538 172614 173294 6 vdd
port 4 nsew power bidirectional
rlabel metal4 s 181994 1538 182614 173294 6 vdd
port 4 nsew power bidirectional
rlabel metal4 s 191994 1538 192614 173294 6 vdd
port 4 nsew power bidirectional
rlabel metal4 s 201994 1538 202614 173294 6 vdd
port 4 nsew power bidirectional
rlabel metal4 s 211994 1538 212614 173294 6 vdd
port 4 nsew power bidirectional
rlabel metal4 s 221994 1538 222614 173294 6 vdd
port 4 nsew power bidirectional
rlabel metal4 s 231994 1538 232614 173294 6 vdd
port 4 nsew power bidirectional
rlabel metal4 s 241994 1538 242614 173294 6 vdd
port 4 nsew power bidirectional
rlabel metal4 s 251994 1538 252614 173294 6 vdd
port 4 nsew power bidirectional
rlabel metal4 s 6994 1538 7614 173294 6 vss
port 5 nsew ground bidirectional
rlabel metal4 s 16994 1538 17614 173294 6 vss
port 5 nsew ground bidirectional
rlabel metal4 s 26994 1538 27614 173294 6 vss
port 5 nsew ground bidirectional
rlabel metal4 s 36994 1538 37614 173294 6 vss
port 5 nsew ground bidirectional
rlabel metal4 s 46994 1538 47614 173294 6 vss
port 5 nsew ground bidirectional
rlabel metal4 s 56994 1538 57614 173294 6 vss
port 5 nsew ground bidirectional
rlabel metal4 s 66994 1538 67614 173294 6 vss
port 5 nsew ground bidirectional
rlabel metal4 s 76994 1538 77614 173294 6 vss
port 5 nsew ground bidirectional
rlabel metal4 s 86994 1538 87614 173294 6 vss
port 5 nsew ground bidirectional
rlabel metal4 s 96994 1538 97614 173294 6 vss
port 5 nsew ground bidirectional
rlabel metal4 s 106994 1538 107614 173294 6 vss
port 5 nsew ground bidirectional
rlabel metal4 s 116994 1538 117614 173294 6 vss
port 5 nsew ground bidirectional
rlabel metal4 s 126994 1538 127614 173294 6 vss
port 5 nsew ground bidirectional
rlabel metal4 s 136994 1538 137614 173294 6 vss
port 5 nsew ground bidirectional
rlabel metal4 s 146994 1538 147614 173294 6 vss
port 5 nsew ground bidirectional
rlabel metal4 s 156994 1538 157614 173294 6 vss
port 5 nsew ground bidirectional
rlabel metal4 s 166994 1538 167614 173294 6 vss
port 5 nsew ground bidirectional
rlabel metal4 s 176994 1538 177614 173294 6 vss
port 5 nsew ground bidirectional
rlabel metal4 s 186994 1538 187614 173294 6 vss
port 5 nsew ground bidirectional
rlabel metal4 s 196994 1538 197614 173294 6 vss
port 5 nsew ground bidirectional
rlabel metal4 s 206994 1538 207614 173294 6 vss
port 5 nsew ground bidirectional
rlabel metal4 s 216994 1538 217614 173294 6 vss
port 5 nsew ground bidirectional
rlabel metal4 s 226994 1538 227614 173294 6 vss
port 5 nsew ground bidirectional
rlabel metal4 s 236994 1538 237614 173294 6 vss
port 5 nsew ground bidirectional
rlabel metal4 s 246994 1538 247614 173294 6 vss
port 5 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 255000 175000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 34063102
string GDS_FILE /home/farag/carvel_riscv_soc/gf180mcu_riscv_soc/openlane/analog_wrapper/runs/23_11_26_00_39/results/signoff/analog_wrapper.magic.gds
string GDS_START 49968
<< end >>

