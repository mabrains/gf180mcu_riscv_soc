magic
tech gf180mcuD
magscale 1 5
timestamp 1700131923
<< obsm1 >>
rect 672 1538 89320 98937
<< metal2 >>
rect 2352 99600 2408 100000
rect 2912 99600 2968 100000
rect 3472 99600 3528 100000
rect 4032 99600 4088 100000
rect 4592 99600 4648 100000
rect 5152 99600 5208 100000
rect 5712 99600 5768 100000
rect 6272 99600 6328 100000
rect 6832 99600 6888 100000
rect 7392 99600 7448 100000
rect 7952 99600 8008 100000
rect 8512 99600 8568 100000
rect 9072 99600 9128 100000
rect 9632 99600 9688 100000
rect 10192 99600 10248 100000
rect 10752 99600 10808 100000
rect 11312 99600 11368 100000
rect 11872 99600 11928 100000
rect 12432 99600 12488 100000
rect 12992 99600 13048 100000
rect 13552 99600 13608 100000
rect 14112 99600 14168 100000
rect 14672 99600 14728 100000
rect 15232 99600 15288 100000
rect 15792 99600 15848 100000
rect 16352 99600 16408 100000
rect 16912 99600 16968 100000
rect 17472 99600 17528 100000
rect 18032 99600 18088 100000
rect 18592 99600 18648 100000
rect 19152 99600 19208 100000
rect 19712 99600 19768 100000
rect 20272 99600 20328 100000
rect 20832 99600 20888 100000
rect 21392 99600 21448 100000
rect 21952 99600 22008 100000
rect 22512 99600 22568 100000
rect 23072 99600 23128 100000
rect 23632 99600 23688 100000
rect 24192 99600 24248 100000
rect 24752 99600 24808 100000
rect 25312 99600 25368 100000
rect 25872 99600 25928 100000
rect 26432 99600 26488 100000
rect 26992 99600 27048 100000
rect 27552 99600 27608 100000
rect 28112 99600 28168 100000
rect 28672 99600 28728 100000
rect 29232 99600 29288 100000
rect 29792 99600 29848 100000
rect 30352 99600 30408 100000
rect 30912 99600 30968 100000
rect 31472 99600 31528 100000
rect 32032 99600 32088 100000
rect 32592 99600 32648 100000
rect 33152 99600 33208 100000
rect 33712 99600 33768 100000
rect 34272 99600 34328 100000
rect 34832 99600 34888 100000
rect 35392 99600 35448 100000
rect 35952 99600 36008 100000
rect 36512 99600 36568 100000
rect 37072 99600 37128 100000
rect 37632 99600 37688 100000
rect 38192 99600 38248 100000
rect 38752 99600 38808 100000
rect 39312 99600 39368 100000
rect 39872 99600 39928 100000
rect 40432 99600 40488 100000
rect 40992 99600 41048 100000
rect 41552 99600 41608 100000
rect 42112 99600 42168 100000
rect 42672 99600 42728 100000
rect 43232 99600 43288 100000
rect 43792 99600 43848 100000
rect 44352 99600 44408 100000
rect 44912 99600 44968 100000
rect 45472 99600 45528 100000
rect 46032 99600 46088 100000
rect 46592 99600 46648 100000
rect 47152 99600 47208 100000
rect 47712 99600 47768 100000
rect 48272 99600 48328 100000
rect 48832 99600 48888 100000
rect 49392 99600 49448 100000
rect 49952 99600 50008 100000
rect 50512 99600 50568 100000
rect 51072 99600 51128 100000
rect 51632 99600 51688 100000
rect 52192 99600 52248 100000
rect 52752 99600 52808 100000
rect 53312 99600 53368 100000
rect 53872 99600 53928 100000
rect 54432 99600 54488 100000
rect 54992 99600 55048 100000
rect 55552 99600 55608 100000
rect 56112 99600 56168 100000
rect 56672 99600 56728 100000
rect 57232 99600 57288 100000
rect 57792 99600 57848 100000
rect 58352 99600 58408 100000
rect 58912 99600 58968 100000
rect 59472 99600 59528 100000
rect 60032 99600 60088 100000
rect 60592 99600 60648 100000
rect 61152 99600 61208 100000
rect 61712 99600 61768 100000
rect 62272 99600 62328 100000
rect 62832 99600 62888 100000
rect 63392 99600 63448 100000
rect 63952 99600 64008 100000
rect 64512 99600 64568 100000
rect 65072 99600 65128 100000
rect 65632 99600 65688 100000
rect 66192 99600 66248 100000
rect 66752 99600 66808 100000
rect 67312 99600 67368 100000
rect 67872 99600 67928 100000
rect 68432 99600 68488 100000
rect 68992 99600 69048 100000
rect 69552 99600 69608 100000
rect 70112 99600 70168 100000
rect 70672 99600 70728 100000
rect 71232 99600 71288 100000
rect 71792 99600 71848 100000
rect 72352 99600 72408 100000
rect 72912 99600 72968 100000
rect 73472 99600 73528 100000
rect 74032 99600 74088 100000
rect 74592 99600 74648 100000
rect 75152 99600 75208 100000
rect 75712 99600 75768 100000
rect 76272 99600 76328 100000
rect 76832 99600 76888 100000
rect 77392 99600 77448 100000
rect 77952 99600 78008 100000
rect 78512 99600 78568 100000
rect 79072 99600 79128 100000
rect 79632 99600 79688 100000
rect 80192 99600 80248 100000
rect 80752 99600 80808 100000
rect 81312 99600 81368 100000
rect 81872 99600 81928 100000
rect 82432 99600 82488 100000
rect 82992 99600 83048 100000
rect 83552 99600 83608 100000
rect 84112 99600 84168 100000
rect 84672 99600 84728 100000
rect 85232 99600 85288 100000
rect 85792 99600 85848 100000
rect 86352 99600 86408 100000
rect 86912 99600 86968 100000
rect 87472 99600 87528 100000
rect 1456 0 1512 400
rect 3808 0 3864 400
rect 6160 0 6216 400
rect 8512 0 8568 400
rect 10864 0 10920 400
rect 13216 0 13272 400
rect 15568 0 15624 400
rect 17920 0 17976 400
rect 20272 0 20328 400
rect 22624 0 22680 400
rect 24976 0 25032 400
rect 27328 0 27384 400
rect 29680 0 29736 400
rect 32032 0 32088 400
rect 34384 0 34440 400
rect 36736 0 36792 400
rect 39088 0 39144 400
rect 41440 0 41496 400
rect 43792 0 43848 400
rect 46144 0 46200 400
rect 48496 0 48552 400
rect 50848 0 50904 400
rect 53200 0 53256 400
rect 55552 0 55608 400
rect 57904 0 57960 400
rect 60256 0 60312 400
rect 62608 0 62664 400
rect 64960 0 65016 400
rect 67312 0 67368 400
rect 69664 0 69720 400
rect 72016 0 72072 400
rect 74368 0 74424 400
rect 76720 0 76776 400
rect 79072 0 79128 400
rect 81424 0 81480 400
rect 83776 0 83832 400
rect 86128 0 86184 400
rect 88480 0 88536 400
<< obsm2 >>
rect 798 99570 2322 99666
rect 2438 99570 2882 99666
rect 2998 99570 3442 99666
rect 3558 99570 4002 99666
rect 4118 99570 4562 99666
rect 4678 99570 5122 99666
rect 5238 99570 5682 99666
rect 5798 99570 6242 99666
rect 6358 99570 6802 99666
rect 6918 99570 7362 99666
rect 7478 99570 7922 99666
rect 8038 99570 8482 99666
rect 8598 99570 9042 99666
rect 9158 99570 9602 99666
rect 9718 99570 10162 99666
rect 10278 99570 10722 99666
rect 10838 99570 11282 99666
rect 11398 99570 11842 99666
rect 11958 99570 12402 99666
rect 12518 99570 12962 99666
rect 13078 99570 13522 99666
rect 13638 99570 14082 99666
rect 14198 99570 14642 99666
rect 14758 99570 15202 99666
rect 15318 99570 15762 99666
rect 15878 99570 16322 99666
rect 16438 99570 16882 99666
rect 16998 99570 17442 99666
rect 17558 99570 18002 99666
rect 18118 99570 18562 99666
rect 18678 99570 19122 99666
rect 19238 99570 19682 99666
rect 19798 99570 20242 99666
rect 20358 99570 20802 99666
rect 20918 99570 21362 99666
rect 21478 99570 21922 99666
rect 22038 99570 22482 99666
rect 22598 99570 23042 99666
rect 23158 99570 23602 99666
rect 23718 99570 24162 99666
rect 24278 99570 24722 99666
rect 24838 99570 25282 99666
rect 25398 99570 25842 99666
rect 25958 99570 26402 99666
rect 26518 99570 26962 99666
rect 27078 99570 27522 99666
rect 27638 99570 28082 99666
rect 28198 99570 28642 99666
rect 28758 99570 29202 99666
rect 29318 99570 29762 99666
rect 29878 99570 30322 99666
rect 30438 99570 30882 99666
rect 30998 99570 31442 99666
rect 31558 99570 32002 99666
rect 32118 99570 32562 99666
rect 32678 99570 33122 99666
rect 33238 99570 33682 99666
rect 33798 99570 34242 99666
rect 34358 99570 34802 99666
rect 34918 99570 35362 99666
rect 35478 99570 35922 99666
rect 36038 99570 36482 99666
rect 36598 99570 37042 99666
rect 37158 99570 37602 99666
rect 37718 99570 38162 99666
rect 38278 99570 38722 99666
rect 38838 99570 39282 99666
rect 39398 99570 39842 99666
rect 39958 99570 40402 99666
rect 40518 99570 40962 99666
rect 41078 99570 41522 99666
rect 41638 99570 42082 99666
rect 42198 99570 42642 99666
rect 42758 99570 43202 99666
rect 43318 99570 43762 99666
rect 43878 99570 44322 99666
rect 44438 99570 44882 99666
rect 44998 99570 45442 99666
rect 45558 99570 46002 99666
rect 46118 99570 46562 99666
rect 46678 99570 47122 99666
rect 47238 99570 47682 99666
rect 47798 99570 48242 99666
rect 48358 99570 48802 99666
rect 48918 99570 49362 99666
rect 49478 99570 49922 99666
rect 50038 99570 50482 99666
rect 50598 99570 51042 99666
rect 51158 99570 51602 99666
rect 51718 99570 52162 99666
rect 52278 99570 52722 99666
rect 52838 99570 53282 99666
rect 53398 99570 53842 99666
rect 53958 99570 54402 99666
rect 54518 99570 54962 99666
rect 55078 99570 55522 99666
rect 55638 99570 56082 99666
rect 56198 99570 56642 99666
rect 56758 99570 57202 99666
rect 57318 99570 57762 99666
rect 57878 99570 58322 99666
rect 58438 99570 58882 99666
rect 58998 99570 59442 99666
rect 59558 99570 60002 99666
rect 60118 99570 60562 99666
rect 60678 99570 61122 99666
rect 61238 99570 61682 99666
rect 61798 99570 62242 99666
rect 62358 99570 62802 99666
rect 62918 99570 63362 99666
rect 63478 99570 63922 99666
rect 64038 99570 64482 99666
rect 64598 99570 65042 99666
rect 65158 99570 65602 99666
rect 65718 99570 66162 99666
rect 66278 99570 66722 99666
rect 66838 99570 67282 99666
rect 67398 99570 67842 99666
rect 67958 99570 68402 99666
rect 68518 99570 68962 99666
rect 69078 99570 69522 99666
rect 69638 99570 70082 99666
rect 70198 99570 70642 99666
rect 70758 99570 71202 99666
rect 71318 99570 71762 99666
rect 71878 99570 72322 99666
rect 72438 99570 72882 99666
rect 72998 99570 73442 99666
rect 73558 99570 74002 99666
rect 74118 99570 74562 99666
rect 74678 99570 75122 99666
rect 75238 99570 75682 99666
rect 75798 99570 76242 99666
rect 76358 99570 76802 99666
rect 76918 99570 77362 99666
rect 77478 99570 77922 99666
rect 78038 99570 78482 99666
rect 78598 99570 79042 99666
rect 79158 99570 79602 99666
rect 79718 99570 80162 99666
rect 80278 99570 80722 99666
rect 80838 99570 81282 99666
rect 81398 99570 81842 99666
rect 81958 99570 82402 99666
rect 82518 99570 82962 99666
rect 83078 99570 83522 99666
rect 83638 99570 84082 99666
rect 84198 99570 84642 99666
rect 84758 99570 85202 99666
rect 85318 99570 85762 99666
rect 85878 99570 86322 99666
rect 86438 99570 86882 99666
rect 86998 99570 87442 99666
rect 87558 99570 89250 99666
rect 798 430 89250 99570
rect 798 350 1426 430
rect 1542 350 3778 430
rect 3894 350 6130 430
rect 6246 350 8482 430
rect 8598 350 10834 430
rect 10950 350 13186 430
rect 13302 350 15538 430
rect 15654 350 17890 430
rect 18006 350 20242 430
rect 20358 350 22594 430
rect 22710 350 24946 430
rect 25062 350 27298 430
rect 27414 350 29650 430
rect 29766 350 32002 430
rect 32118 350 34354 430
rect 34470 350 36706 430
rect 36822 350 39058 430
rect 39174 350 41410 430
rect 41526 350 43762 430
rect 43878 350 46114 430
rect 46230 350 48466 430
rect 48582 350 50818 430
rect 50934 350 53170 430
rect 53286 350 55522 430
rect 55638 350 57874 430
rect 57990 350 60226 430
rect 60342 350 62578 430
rect 62694 350 64930 430
rect 65046 350 67282 430
rect 67398 350 69634 430
rect 69750 350 71986 430
rect 72102 350 74338 430
rect 74454 350 76690 430
rect 76806 350 79042 430
rect 79158 350 81394 430
rect 81510 350 83746 430
rect 83862 350 86098 430
rect 86214 350 88450 430
rect 88566 350 89250 430
<< metal3 >>
rect 0 96992 400 97048
rect 89600 96768 90000 96824
rect 0 95872 400 95928
rect 0 94752 400 94808
rect 89600 94640 90000 94696
rect 0 93632 400 93688
rect 0 92512 400 92568
rect 89600 92512 90000 92568
rect 0 91392 400 91448
rect 89600 90384 90000 90440
rect 0 90272 400 90328
rect 0 89152 400 89208
rect 89600 88256 90000 88312
rect 0 88032 400 88088
rect 0 86912 400 86968
rect 89600 86128 90000 86184
rect 0 85792 400 85848
rect 0 84672 400 84728
rect 89600 84000 90000 84056
rect 0 83552 400 83608
rect 0 82432 400 82488
rect 89600 81872 90000 81928
rect 0 81312 400 81368
rect 0 80192 400 80248
rect 89600 79744 90000 79800
rect 0 79072 400 79128
rect 0 77952 400 78008
rect 89600 77616 90000 77672
rect 0 76832 400 76888
rect 0 75712 400 75768
rect 89600 75488 90000 75544
rect 0 74592 400 74648
rect 0 73472 400 73528
rect 89600 73360 90000 73416
rect 0 72352 400 72408
rect 0 71232 400 71288
rect 89600 71232 90000 71288
rect 0 70112 400 70168
rect 89600 69104 90000 69160
rect 0 68992 400 69048
rect 0 67872 400 67928
rect 89600 66976 90000 67032
rect 0 66752 400 66808
rect 0 65632 400 65688
rect 89600 64848 90000 64904
rect 0 64512 400 64568
rect 0 63392 400 63448
rect 89600 62720 90000 62776
rect 0 62272 400 62328
rect 0 61152 400 61208
rect 89600 60592 90000 60648
rect 0 60032 400 60088
rect 0 58912 400 58968
rect 89600 58464 90000 58520
rect 0 57792 400 57848
rect 0 56672 400 56728
rect 89600 56336 90000 56392
rect 0 55552 400 55608
rect 0 54432 400 54488
rect 89600 54208 90000 54264
rect 0 53312 400 53368
rect 0 52192 400 52248
rect 89600 52080 90000 52136
rect 0 51072 400 51128
rect 0 49952 400 50008
rect 89600 49952 90000 50008
rect 0 48832 400 48888
rect 89600 47824 90000 47880
rect 0 47712 400 47768
rect 0 46592 400 46648
rect 89600 45696 90000 45752
rect 0 45472 400 45528
rect 0 44352 400 44408
rect 89600 43568 90000 43624
rect 0 43232 400 43288
rect 0 42112 400 42168
rect 89600 41440 90000 41496
rect 0 40992 400 41048
rect 0 39872 400 39928
rect 89600 39312 90000 39368
rect 0 38752 400 38808
rect 0 37632 400 37688
rect 89600 37184 90000 37240
rect 0 36512 400 36568
rect 0 35392 400 35448
rect 89600 35056 90000 35112
rect 0 34272 400 34328
rect 0 33152 400 33208
rect 89600 32928 90000 32984
rect 0 32032 400 32088
rect 0 30912 400 30968
rect 89600 30800 90000 30856
rect 0 29792 400 29848
rect 0 28672 400 28728
rect 89600 28672 90000 28728
rect 0 27552 400 27608
rect 89600 26544 90000 26600
rect 0 26432 400 26488
rect 0 25312 400 25368
rect 89600 24416 90000 24472
rect 0 24192 400 24248
rect 0 23072 400 23128
rect 89600 22288 90000 22344
rect 0 21952 400 22008
rect 0 20832 400 20888
rect 89600 20160 90000 20216
rect 0 19712 400 19768
rect 0 18592 400 18648
rect 89600 18032 90000 18088
rect 0 17472 400 17528
rect 0 16352 400 16408
rect 89600 15904 90000 15960
rect 0 15232 400 15288
rect 0 14112 400 14168
rect 89600 13776 90000 13832
rect 0 12992 400 13048
rect 0 11872 400 11928
rect 89600 11648 90000 11704
rect 0 10752 400 10808
rect 0 9632 400 9688
rect 89600 9520 90000 9576
rect 0 8512 400 8568
rect 0 7392 400 7448
rect 89600 7392 90000 7448
rect 0 6272 400 6328
rect 89600 5264 90000 5320
rect 0 5152 400 5208
rect 0 4032 400 4088
rect 89600 3136 90000 3192
rect 0 2912 400 2968
<< obsm3 >>
rect 400 97078 89600 98406
rect 430 96962 89600 97078
rect 400 96854 89600 96962
rect 400 96738 89570 96854
rect 400 95958 89600 96738
rect 430 95842 89600 95958
rect 400 94838 89600 95842
rect 430 94726 89600 94838
rect 430 94722 89570 94726
rect 400 94610 89570 94722
rect 400 93718 89600 94610
rect 430 93602 89600 93718
rect 400 92598 89600 93602
rect 430 92482 89570 92598
rect 400 91478 89600 92482
rect 430 91362 89600 91478
rect 400 90470 89600 91362
rect 400 90358 89570 90470
rect 430 90354 89570 90358
rect 430 90242 89600 90354
rect 400 89238 89600 90242
rect 430 89122 89600 89238
rect 400 88342 89600 89122
rect 400 88226 89570 88342
rect 400 88118 89600 88226
rect 430 88002 89600 88118
rect 400 86998 89600 88002
rect 430 86882 89600 86998
rect 400 86214 89600 86882
rect 400 86098 89570 86214
rect 400 85878 89600 86098
rect 430 85762 89600 85878
rect 400 84758 89600 85762
rect 430 84642 89600 84758
rect 400 84086 89600 84642
rect 400 83970 89570 84086
rect 400 83638 89600 83970
rect 430 83522 89600 83638
rect 400 82518 89600 83522
rect 430 82402 89600 82518
rect 400 81958 89600 82402
rect 400 81842 89570 81958
rect 400 81398 89600 81842
rect 430 81282 89600 81398
rect 400 80278 89600 81282
rect 430 80162 89600 80278
rect 400 79830 89600 80162
rect 400 79714 89570 79830
rect 400 79158 89600 79714
rect 430 79042 89600 79158
rect 400 78038 89600 79042
rect 430 77922 89600 78038
rect 400 77702 89600 77922
rect 400 77586 89570 77702
rect 400 76918 89600 77586
rect 430 76802 89600 76918
rect 400 75798 89600 76802
rect 430 75682 89600 75798
rect 400 75574 89600 75682
rect 400 75458 89570 75574
rect 400 74678 89600 75458
rect 430 74562 89600 74678
rect 400 73558 89600 74562
rect 430 73446 89600 73558
rect 430 73442 89570 73446
rect 400 73330 89570 73442
rect 400 72438 89600 73330
rect 430 72322 89600 72438
rect 400 71318 89600 72322
rect 430 71202 89570 71318
rect 400 70198 89600 71202
rect 430 70082 89600 70198
rect 400 69190 89600 70082
rect 400 69078 89570 69190
rect 430 69074 89570 69078
rect 430 68962 89600 69074
rect 400 67958 89600 68962
rect 430 67842 89600 67958
rect 400 67062 89600 67842
rect 400 66946 89570 67062
rect 400 66838 89600 66946
rect 430 66722 89600 66838
rect 400 65718 89600 66722
rect 430 65602 89600 65718
rect 400 64934 89600 65602
rect 400 64818 89570 64934
rect 400 64598 89600 64818
rect 430 64482 89600 64598
rect 400 63478 89600 64482
rect 430 63362 89600 63478
rect 400 62806 89600 63362
rect 400 62690 89570 62806
rect 400 62358 89600 62690
rect 430 62242 89600 62358
rect 400 61238 89600 62242
rect 430 61122 89600 61238
rect 400 60678 89600 61122
rect 400 60562 89570 60678
rect 400 60118 89600 60562
rect 430 60002 89600 60118
rect 400 58998 89600 60002
rect 430 58882 89600 58998
rect 400 58550 89600 58882
rect 400 58434 89570 58550
rect 400 57878 89600 58434
rect 430 57762 89600 57878
rect 400 56758 89600 57762
rect 430 56642 89600 56758
rect 400 56422 89600 56642
rect 400 56306 89570 56422
rect 400 55638 89600 56306
rect 430 55522 89600 55638
rect 400 54518 89600 55522
rect 430 54402 89600 54518
rect 400 54294 89600 54402
rect 400 54178 89570 54294
rect 400 53398 89600 54178
rect 430 53282 89600 53398
rect 400 52278 89600 53282
rect 430 52166 89600 52278
rect 430 52162 89570 52166
rect 400 52050 89570 52162
rect 400 51158 89600 52050
rect 430 51042 89600 51158
rect 400 50038 89600 51042
rect 430 49922 89570 50038
rect 400 48918 89600 49922
rect 430 48802 89600 48918
rect 400 47910 89600 48802
rect 400 47798 89570 47910
rect 430 47794 89570 47798
rect 430 47682 89600 47794
rect 400 46678 89600 47682
rect 430 46562 89600 46678
rect 400 45782 89600 46562
rect 400 45666 89570 45782
rect 400 45558 89600 45666
rect 430 45442 89600 45558
rect 400 44438 89600 45442
rect 430 44322 89600 44438
rect 400 43654 89600 44322
rect 400 43538 89570 43654
rect 400 43318 89600 43538
rect 430 43202 89600 43318
rect 400 42198 89600 43202
rect 430 42082 89600 42198
rect 400 41526 89600 42082
rect 400 41410 89570 41526
rect 400 41078 89600 41410
rect 430 40962 89600 41078
rect 400 39958 89600 40962
rect 430 39842 89600 39958
rect 400 39398 89600 39842
rect 400 39282 89570 39398
rect 400 38838 89600 39282
rect 430 38722 89600 38838
rect 400 37718 89600 38722
rect 430 37602 89600 37718
rect 400 37270 89600 37602
rect 400 37154 89570 37270
rect 400 36598 89600 37154
rect 430 36482 89600 36598
rect 400 35478 89600 36482
rect 430 35362 89600 35478
rect 400 35142 89600 35362
rect 400 35026 89570 35142
rect 400 34358 89600 35026
rect 430 34242 89600 34358
rect 400 33238 89600 34242
rect 430 33122 89600 33238
rect 400 33014 89600 33122
rect 400 32898 89570 33014
rect 400 32118 89600 32898
rect 430 32002 89600 32118
rect 400 30998 89600 32002
rect 430 30886 89600 30998
rect 430 30882 89570 30886
rect 400 30770 89570 30882
rect 400 29878 89600 30770
rect 430 29762 89600 29878
rect 400 28758 89600 29762
rect 430 28642 89570 28758
rect 400 27638 89600 28642
rect 430 27522 89600 27638
rect 400 26630 89600 27522
rect 400 26518 89570 26630
rect 430 26514 89570 26518
rect 430 26402 89600 26514
rect 400 25398 89600 26402
rect 430 25282 89600 25398
rect 400 24502 89600 25282
rect 400 24386 89570 24502
rect 400 24278 89600 24386
rect 430 24162 89600 24278
rect 400 23158 89600 24162
rect 430 23042 89600 23158
rect 400 22374 89600 23042
rect 400 22258 89570 22374
rect 400 22038 89600 22258
rect 430 21922 89600 22038
rect 400 20918 89600 21922
rect 430 20802 89600 20918
rect 400 20246 89600 20802
rect 400 20130 89570 20246
rect 400 19798 89600 20130
rect 430 19682 89600 19798
rect 400 18678 89600 19682
rect 430 18562 89600 18678
rect 400 18118 89600 18562
rect 400 18002 89570 18118
rect 400 17558 89600 18002
rect 430 17442 89600 17558
rect 400 16438 89600 17442
rect 430 16322 89600 16438
rect 400 15990 89600 16322
rect 400 15874 89570 15990
rect 400 15318 89600 15874
rect 430 15202 89600 15318
rect 400 14198 89600 15202
rect 430 14082 89600 14198
rect 400 13862 89600 14082
rect 400 13746 89570 13862
rect 400 13078 89600 13746
rect 430 12962 89600 13078
rect 400 11958 89600 12962
rect 430 11842 89600 11958
rect 400 11734 89600 11842
rect 400 11618 89570 11734
rect 400 10838 89600 11618
rect 430 10722 89600 10838
rect 400 9718 89600 10722
rect 430 9606 89600 9718
rect 430 9602 89570 9606
rect 400 9490 89570 9602
rect 400 8598 89600 9490
rect 430 8482 89600 8598
rect 400 7478 89600 8482
rect 430 7362 89570 7478
rect 400 6358 89600 7362
rect 430 6242 89600 6358
rect 400 5350 89600 6242
rect 400 5238 89570 5350
rect 430 5234 89570 5238
rect 430 5122 89600 5234
rect 400 4118 89600 5122
rect 430 4002 89600 4118
rect 400 3222 89600 4002
rect 400 3106 89570 3222
rect 400 2998 89600 3106
rect 430 2882 89600 2998
rect 400 1554 89600 2882
<< metal4 >>
rect 2224 1538 2384 98422
rect 9904 1538 10064 98422
rect 17584 1538 17744 98422
rect 25264 1538 25424 98422
rect 32944 1538 33104 98422
rect 40624 1538 40784 98422
rect 48304 1538 48464 98422
rect 55984 1538 56144 98422
rect 63664 1538 63824 98422
rect 71344 1538 71504 98422
rect 79024 1538 79184 98422
rect 86704 1538 86864 98422
<< obsm4 >>
rect 1134 1801 2194 98103
rect 2414 1801 9874 98103
rect 10094 1801 17554 98103
rect 17774 1801 25234 98103
rect 25454 1801 32914 98103
rect 33134 1801 40594 98103
rect 40814 1801 48274 98103
rect 48494 1801 55954 98103
rect 56174 1801 63634 98103
rect 63854 1801 71314 98103
rect 71534 1801 78994 98103
rect 79214 1801 86674 98103
rect 86894 1801 88802 98103
<< obsm5 >>
rect 1126 13073 86010 97807
<< labels >>
rlabel metal4 s 2224 1538 2384 98422 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 98422 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 98422 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 98422 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 63664 1538 63824 98422 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 79024 1538 79184 98422 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 98422 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 98422 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 98422 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 98422 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 71344 1538 71504 98422 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 86704 1538 86864 98422 6 VSS
port 2 nsew ground bidirectional
rlabel metal3 s 89600 3136 90000 3192 6 digital_io_in[0]
port 3 nsew signal input
rlabel metal3 s 89600 66976 90000 67032 6 digital_io_in[10]
port 4 nsew signal input
rlabel metal3 s 89600 73360 90000 73416 6 digital_io_in[11]
port 5 nsew signal input
rlabel metal3 s 89600 79744 90000 79800 6 digital_io_in[12]
port 6 nsew signal input
rlabel metal3 s 89600 86128 90000 86184 6 digital_io_in[13]
port 7 nsew signal input
rlabel metal3 s 89600 92512 90000 92568 6 digital_io_in[14]
port 8 nsew signal input
rlabel metal2 s 86352 99600 86408 100000 6 digital_io_in[15]
port 9 nsew signal input
rlabel metal2 s 84672 99600 84728 100000 6 digital_io_in[16]
port 10 nsew signal input
rlabel metal2 s 82992 99600 83048 100000 6 digital_io_in[17]
port 11 nsew signal input
rlabel metal2 s 81312 99600 81368 100000 6 digital_io_in[18]
port 12 nsew signal input
rlabel metal2 s 79632 99600 79688 100000 6 digital_io_in[19]
port 13 nsew signal input
rlabel metal3 s 89600 9520 90000 9576 6 digital_io_in[1]
port 14 nsew signal input
rlabel metal2 s 77952 99600 78008 100000 6 digital_io_in[20]
port 15 nsew signal input
rlabel metal2 s 76272 99600 76328 100000 6 digital_io_in[21]
port 16 nsew signal input
rlabel metal2 s 74592 99600 74648 100000 6 digital_io_in[22]
port 17 nsew signal input
rlabel metal2 s 72912 99600 72968 100000 6 digital_io_in[23]
port 18 nsew signal input
rlabel metal2 s 25312 99600 25368 100000 6 digital_io_in[24]
port 19 nsew signal input
rlabel metal2 s 23632 99600 23688 100000 6 digital_io_in[25]
port 20 nsew signal input
rlabel metal2 s 21952 99600 22008 100000 6 digital_io_in[26]
port 21 nsew signal input
rlabel metal2 s 20272 99600 20328 100000 6 digital_io_in[27]
port 22 nsew signal input
rlabel metal2 s 18592 99600 18648 100000 6 digital_io_in[28]
port 23 nsew signal input
rlabel metal2 s 16912 99600 16968 100000 6 digital_io_in[29]
port 24 nsew signal input
rlabel metal3 s 89600 15904 90000 15960 6 digital_io_in[2]
port 25 nsew signal input
rlabel metal2 s 15232 99600 15288 100000 6 digital_io_in[30]
port 26 nsew signal input
rlabel metal2 s 13552 99600 13608 100000 6 digital_io_in[31]
port 27 nsew signal input
rlabel metal2 s 11872 99600 11928 100000 6 digital_io_in[32]
port 28 nsew signal input
rlabel metal2 s 10192 99600 10248 100000 6 digital_io_in[33]
port 29 nsew signal input
rlabel metal2 s 8512 99600 8568 100000 6 digital_io_in[34]
port 30 nsew signal input
rlabel metal2 s 6832 99600 6888 100000 6 digital_io_in[35]
port 31 nsew signal input
rlabel metal2 s 5152 99600 5208 100000 6 digital_io_in[36]
port 32 nsew signal input
rlabel metal2 s 3472 99600 3528 100000 6 digital_io_in[37]
port 33 nsew signal input
rlabel metal3 s 89600 22288 90000 22344 6 digital_io_in[3]
port 34 nsew signal input
rlabel metal3 s 89600 28672 90000 28728 6 digital_io_in[4]
port 35 nsew signal input
rlabel metal3 s 89600 35056 90000 35112 6 digital_io_in[5]
port 36 nsew signal input
rlabel metal3 s 89600 41440 90000 41496 6 digital_io_in[6]
port 37 nsew signal input
rlabel metal3 s 89600 47824 90000 47880 6 digital_io_in[7]
port 38 nsew signal input
rlabel metal3 s 89600 54208 90000 54264 6 digital_io_in[8]
port 39 nsew signal input
rlabel metal3 s 89600 60592 90000 60648 6 digital_io_in[9]
port 40 nsew signal input
rlabel metal3 s 89600 7392 90000 7448 6 digital_io_oen[0]
port 41 nsew signal output
rlabel metal3 s 89600 71232 90000 71288 6 digital_io_oen[10]
port 42 nsew signal output
rlabel metal3 s 89600 77616 90000 77672 6 digital_io_oen[11]
port 43 nsew signal output
rlabel metal3 s 89600 84000 90000 84056 6 digital_io_oen[12]
port 44 nsew signal output
rlabel metal3 s 89600 90384 90000 90440 6 digital_io_oen[13]
port 45 nsew signal output
rlabel metal3 s 89600 96768 90000 96824 6 digital_io_oen[14]
port 46 nsew signal output
rlabel metal2 s 87472 99600 87528 100000 6 digital_io_oen[15]
port 47 nsew signal output
rlabel metal2 s 85792 99600 85848 100000 6 digital_io_oen[16]
port 48 nsew signal output
rlabel metal2 s 84112 99600 84168 100000 6 digital_io_oen[17]
port 49 nsew signal output
rlabel metal2 s 82432 99600 82488 100000 6 digital_io_oen[18]
port 50 nsew signal output
rlabel metal2 s 80752 99600 80808 100000 6 digital_io_oen[19]
port 51 nsew signal output
rlabel metal3 s 89600 13776 90000 13832 6 digital_io_oen[1]
port 52 nsew signal output
rlabel metal2 s 79072 99600 79128 100000 6 digital_io_oen[20]
port 53 nsew signal output
rlabel metal2 s 77392 99600 77448 100000 6 digital_io_oen[21]
port 54 nsew signal output
rlabel metal2 s 75712 99600 75768 100000 6 digital_io_oen[22]
port 55 nsew signal output
rlabel metal2 s 74032 99600 74088 100000 6 digital_io_oen[23]
port 56 nsew signal output
rlabel metal2 s 24192 99600 24248 100000 6 digital_io_oen[24]
port 57 nsew signal output
rlabel metal2 s 22512 99600 22568 100000 6 digital_io_oen[25]
port 58 nsew signal output
rlabel metal2 s 20832 99600 20888 100000 6 digital_io_oen[26]
port 59 nsew signal output
rlabel metal2 s 19152 99600 19208 100000 6 digital_io_oen[27]
port 60 nsew signal output
rlabel metal2 s 17472 99600 17528 100000 6 digital_io_oen[28]
port 61 nsew signal output
rlabel metal2 s 15792 99600 15848 100000 6 digital_io_oen[29]
port 62 nsew signal output
rlabel metal3 s 89600 20160 90000 20216 6 digital_io_oen[2]
port 63 nsew signal output
rlabel metal2 s 14112 99600 14168 100000 6 digital_io_oen[30]
port 64 nsew signal output
rlabel metal2 s 12432 99600 12488 100000 6 digital_io_oen[31]
port 65 nsew signal output
rlabel metal2 s 10752 99600 10808 100000 6 digital_io_oen[32]
port 66 nsew signal output
rlabel metal2 s 9072 99600 9128 100000 6 digital_io_oen[33]
port 67 nsew signal output
rlabel metal2 s 7392 99600 7448 100000 6 digital_io_oen[34]
port 68 nsew signal output
rlabel metal2 s 5712 99600 5768 100000 6 digital_io_oen[35]
port 69 nsew signal output
rlabel metal2 s 4032 99600 4088 100000 6 digital_io_oen[36]
port 70 nsew signal output
rlabel metal2 s 2352 99600 2408 100000 6 digital_io_oen[37]
port 71 nsew signal output
rlabel metal3 s 89600 26544 90000 26600 6 digital_io_oen[3]
port 72 nsew signal output
rlabel metal3 s 89600 32928 90000 32984 6 digital_io_oen[4]
port 73 nsew signal output
rlabel metal3 s 89600 39312 90000 39368 6 digital_io_oen[5]
port 74 nsew signal output
rlabel metal3 s 89600 45696 90000 45752 6 digital_io_oen[6]
port 75 nsew signal output
rlabel metal3 s 89600 52080 90000 52136 6 digital_io_oen[7]
port 76 nsew signal output
rlabel metal3 s 89600 58464 90000 58520 6 digital_io_oen[8]
port 77 nsew signal output
rlabel metal3 s 89600 64848 90000 64904 6 digital_io_oen[9]
port 78 nsew signal output
rlabel metal3 s 89600 5264 90000 5320 6 digital_io_out[0]
port 79 nsew signal output
rlabel metal3 s 89600 69104 90000 69160 6 digital_io_out[10]
port 80 nsew signal output
rlabel metal3 s 89600 75488 90000 75544 6 digital_io_out[11]
port 81 nsew signal output
rlabel metal3 s 89600 81872 90000 81928 6 digital_io_out[12]
port 82 nsew signal output
rlabel metal3 s 89600 88256 90000 88312 6 digital_io_out[13]
port 83 nsew signal output
rlabel metal3 s 89600 94640 90000 94696 6 digital_io_out[14]
port 84 nsew signal output
rlabel metal2 s 86912 99600 86968 100000 6 digital_io_out[15]
port 85 nsew signal output
rlabel metal2 s 85232 99600 85288 100000 6 digital_io_out[16]
port 86 nsew signal output
rlabel metal2 s 83552 99600 83608 100000 6 digital_io_out[17]
port 87 nsew signal output
rlabel metal2 s 81872 99600 81928 100000 6 digital_io_out[18]
port 88 nsew signal output
rlabel metal2 s 80192 99600 80248 100000 6 digital_io_out[19]
port 89 nsew signal output
rlabel metal3 s 89600 11648 90000 11704 6 digital_io_out[1]
port 90 nsew signal output
rlabel metal2 s 78512 99600 78568 100000 6 digital_io_out[20]
port 91 nsew signal output
rlabel metal2 s 76832 99600 76888 100000 6 digital_io_out[21]
port 92 nsew signal output
rlabel metal2 s 75152 99600 75208 100000 6 digital_io_out[22]
port 93 nsew signal output
rlabel metal2 s 73472 99600 73528 100000 6 digital_io_out[23]
port 94 nsew signal output
rlabel metal2 s 24752 99600 24808 100000 6 digital_io_out[24]
port 95 nsew signal output
rlabel metal2 s 23072 99600 23128 100000 6 digital_io_out[25]
port 96 nsew signal output
rlabel metal2 s 21392 99600 21448 100000 6 digital_io_out[26]
port 97 nsew signal output
rlabel metal2 s 19712 99600 19768 100000 6 digital_io_out[27]
port 98 nsew signal output
rlabel metal2 s 18032 99600 18088 100000 6 digital_io_out[28]
port 99 nsew signal output
rlabel metal2 s 16352 99600 16408 100000 6 digital_io_out[29]
port 100 nsew signal output
rlabel metal3 s 89600 18032 90000 18088 6 digital_io_out[2]
port 101 nsew signal output
rlabel metal2 s 14672 99600 14728 100000 6 digital_io_out[30]
port 102 nsew signal output
rlabel metal2 s 12992 99600 13048 100000 6 digital_io_out[31]
port 103 nsew signal output
rlabel metal2 s 11312 99600 11368 100000 6 digital_io_out[32]
port 104 nsew signal output
rlabel metal2 s 9632 99600 9688 100000 6 digital_io_out[33]
port 105 nsew signal output
rlabel metal2 s 7952 99600 8008 100000 6 digital_io_out[34]
port 106 nsew signal output
rlabel metal2 s 6272 99600 6328 100000 6 digital_io_out[35]
port 107 nsew signal output
rlabel metal2 s 4592 99600 4648 100000 6 digital_io_out[36]
port 108 nsew signal output
rlabel metal2 s 2912 99600 2968 100000 6 digital_io_out[37]
port 109 nsew signal output
rlabel metal3 s 89600 24416 90000 24472 6 digital_io_out[3]
port 110 nsew signal output
rlabel metal3 s 89600 30800 90000 30856 6 digital_io_out[4]
port 111 nsew signal output
rlabel metal3 s 89600 37184 90000 37240 6 digital_io_out[5]
port 112 nsew signal output
rlabel metal3 s 89600 43568 90000 43624 6 digital_io_out[6]
port 113 nsew signal output
rlabel metal3 s 89600 49952 90000 50008 6 digital_io_out[7]
port 114 nsew signal output
rlabel metal3 s 89600 56336 90000 56392 6 digital_io_out[8]
port 115 nsew signal output
rlabel metal3 s 89600 62720 90000 62776 6 digital_io_out[9]
port 116 nsew signal output
rlabel metal3 s 0 4032 400 4088 6 e_reset_n
port 117 nsew signal input
rlabel metal2 s 43792 0 43848 400 6 i2cm_clk_i
port 118 nsew signal output
rlabel metal2 s 41440 0 41496 400 6 i2cm_clk_o
port 119 nsew signal input
rlabel metal2 s 46144 0 46200 400 6 i2cm_clk_oen
port 120 nsew signal input
rlabel metal2 s 53200 0 53256 400 6 i2cm_data_i
port 121 nsew signal output
rlabel metal2 s 50848 0 50904 400 6 i2cm_data_o
port 122 nsew signal input
rlabel metal2 s 48496 0 48552 400 6 i2cm_data_oen
port 123 nsew signal input
rlabel metal2 s 74368 0 74424 400 6 i2cm_intr
port 124 nsew signal input
rlabel metal2 s 8512 0 8568 400 6 i2cm_rst_n
port 125 nsew signal output
rlabel metal3 s 0 5152 400 5208 6 mclk
port 126 nsew signal input
rlabel metal3 s 0 2912 400 2968 6 p_reset_n
port 127 nsew signal input
rlabel metal2 s 72016 0 72072 400 6 pulse1m_mclk
port 128 nsew signal output
rlabel metal3 s 0 96992 400 97048 6 reg_ack
port 129 nsew signal output
rlabel metal3 s 0 19712 400 19768 6 reg_addr[0]
port 130 nsew signal input
rlabel metal3 s 0 8512 400 8568 6 reg_addr[10]
port 131 nsew signal input
rlabel metal3 s 0 18592 400 18648 6 reg_addr[1]
port 132 nsew signal input
rlabel metal3 s 0 17472 400 17528 6 reg_addr[2]
port 133 nsew signal input
rlabel metal3 s 0 16352 400 16408 6 reg_addr[3]
port 134 nsew signal input
rlabel metal3 s 0 15232 400 15288 6 reg_addr[4]
port 135 nsew signal input
rlabel metal3 s 0 14112 400 14168 6 reg_addr[5]
port 136 nsew signal input
rlabel metal3 s 0 12992 400 13048 6 reg_addr[6]
port 137 nsew signal input
rlabel metal3 s 0 11872 400 11928 6 reg_addr[7]
port 138 nsew signal input
rlabel metal3 s 0 10752 400 10808 6 reg_addr[8]
port 139 nsew signal input
rlabel metal3 s 0 9632 400 9688 6 reg_addr[9]
port 140 nsew signal input
rlabel metal3 s 0 24192 400 24248 6 reg_be[0]
port 141 nsew signal input
rlabel metal3 s 0 23072 400 23128 6 reg_be[1]
port 142 nsew signal input
rlabel metal3 s 0 21952 400 22008 6 reg_be[2]
port 143 nsew signal input
rlabel metal3 s 0 20832 400 20888 6 reg_be[3]
port 144 nsew signal input
rlabel metal3 s 0 6272 400 6328 6 reg_cs
port 145 nsew signal input
rlabel metal2 s 72352 99600 72408 100000 6 reg_peri_ack
port 146 nsew signal input
rlabel metal2 s 33712 99600 33768 100000 6 reg_peri_addr[0]
port 147 nsew signal output
rlabel metal2 s 28112 99600 28168 100000 6 reg_peri_addr[10]
port 148 nsew signal output
rlabel metal2 s 33152 99600 33208 100000 6 reg_peri_addr[1]
port 149 nsew signal output
rlabel metal2 s 32592 99600 32648 100000 6 reg_peri_addr[2]
port 150 nsew signal output
rlabel metal2 s 32032 99600 32088 100000 6 reg_peri_addr[3]
port 151 nsew signal output
rlabel metal2 s 31472 99600 31528 100000 6 reg_peri_addr[4]
port 152 nsew signal output
rlabel metal2 s 30912 99600 30968 100000 6 reg_peri_addr[5]
port 153 nsew signal output
rlabel metal2 s 30352 99600 30408 100000 6 reg_peri_addr[6]
port 154 nsew signal output
rlabel metal2 s 29792 99600 29848 100000 6 reg_peri_addr[7]
port 155 nsew signal output
rlabel metal2 s 29232 99600 29288 100000 6 reg_peri_addr[8]
port 156 nsew signal output
rlabel metal2 s 28672 99600 28728 100000 6 reg_peri_addr[9]
port 157 nsew signal output
rlabel metal2 s 35952 99600 36008 100000 6 reg_peri_be[0]
port 158 nsew signal output
rlabel metal2 s 35392 99600 35448 100000 6 reg_peri_be[1]
port 159 nsew signal output
rlabel metal2 s 34832 99600 34888 100000 6 reg_peri_be[2]
port 160 nsew signal output
rlabel metal2 s 34272 99600 34328 100000 6 reg_peri_be[3]
port 161 nsew signal output
rlabel metal2 s 26992 99600 27048 100000 6 reg_peri_cs
port 162 nsew signal output
rlabel metal2 s 71792 99600 71848 100000 6 reg_peri_rdata[0]
port 163 nsew signal input
rlabel metal2 s 66192 99600 66248 100000 6 reg_peri_rdata[10]
port 164 nsew signal input
rlabel metal2 s 65632 99600 65688 100000 6 reg_peri_rdata[11]
port 165 nsew signal input
rlabel metal2 s 65072 99600 65128 100000 6 reg_peri_rdata[12]
port 166 nsew signal input
rlabel metal2 s 64512 99600 64568 100000 6 reg_peri_rdata[13]
port 167 nsew signal input
rlabel metal2 s 63952 99600 64008 100000 6 reg_peri_rdata[14]
port 168 nsew signal input
rlabel metal2 s 63392 99600 63448 100000 6 reg_peri_rdata[15]
port 169 nsew signal input
rlabel metal2 s 62832 99600 62888 100000 6 reg_peri_rdata[16]
port 170 nsew signal input
rlabel metal2 s 62272 99600 62328 100000 6 reg_peri_rdata[17]
port 171 nsew signal input
rlabel metal2 s 61712 99600 61768 100000 6 reg_peri_rdata[18]
port 172 nsew signal input
rlabel metal2 s 61152 99600 61208 100000 6 reg_peri_rdata[19]
port 173 nsew signal input
rlabel metal2 s 71232 99600 71288 100000 6 reg_peri_rdata[1]
port 174 nsew signal input
rlabel metal2 s 60592 99600 60648 100000 6 reg_peri_rdata[20]
port 175 nsew signal input
rlabel metal2 s 60032 99600 60088 100000 6 reg_peri_rdata[21]
port 176 nsew signal input
rlabel metal2 s 59472 99600 59528 100000 6 reg_peri_rdata[22]
port 177 nsew signal input
rlabel metal2 s 58912 99600 58968 100000 6 reg_peri_rdata[23]
port 178 nsew signal input
rlabel metal2 s 58352 99600 58408 100000 6 reg_peri_rdata[24]
port 179 nsew signal input
rlabel metal2 s 57792 99600 57848 100000 6 reg_peri_rdata[25]
port 180 nsew signal input
rlabel metal2 s 57232 99600 57288 100000 6 reg_peri_rdata[26]
port 181 nsew signal input
rlabel metal2 s 56672 99600 56728 100000 6 reg_peri_rdata[27]
port 182 nsew signal input
rlabel metal2 s 56112 99600 56168 100000 6 reg_peri_rdata[28]
port 183 nsew signal input
rlabel metal2 s 55552 99600 55608 100000 6 reg_peri_rdata[29]
port 184 nsew signal input
rlabel metal2 s 70672 99600 70728 100000 6 reg_peri_rdata[2]
port 185 nsew signal input
rlabel metal2 s 54992 99600 55048 100000 6 reg_peri_rdata[30]
port 186 nsew signal input
rlabel metal2 s 54432 99600 54488 100000 6 reg_peri_rdata[31]
port 187 nsew signal input
rlabel metal2 s 70112 99600 70168 100000 6 reg_peri_rdata[3]
port 188 nsew signal input
rlabel metal2 s 69552 99600 69608 100000 6 reg_peri_rdata[4]
port 189 nsew signal input
rlabel metal2 s 68992 99600 69048 100000 6 reg_peri_rdata[5]
port 190 nsew signal input
rlabel metal2 s 68432 99600 68488 100000 6 reg_peri_rdata[6]
port 191 nsew signal input
rlabel metal2 s 67872 99600 67928 100000 6 reg_peri_rdata[7]
port 192 nsew signal input
rlabel metal2 s 67312 99600 67368 100000 6 reg_peri_rdata[8]
port 193 nsew signal input
rlabel metal2 s 66752 99600 66808 100000 6 reg_peri_rdata[9]
port 194 nsew signal input
rlabel metal2 s 53872 99600 53928 100000 6 reg_peri_wdata[0]
port 195 nsew signal output
rlabel metal2 s 48272 99600 48328 100000 6 reg_peri_wdata[10]
port 196 nsew signal output
rlabel metal2 s 47712 99600 47768 100000 6 reg_peri_wdata[11]
port 197 nsew signal output
rlabel metal2 s 47152 99600 47208 100000 6 reg_peri_wdata[12]
port 198 nsew signal output
rlabel metal2 s 46592 99600 46648 100000 6 reg_peri_wdata[13]
port 199 nsew signal output
rlabel metal2 s 46032 99600 46088 100000 6 reg_peri_wdata[14]
port 200 nsew signal output
rlabel metal2 s 45472 99600 45528 100000 6 reg_peri_wdata[15]
port 201 nsew signal output
rlabel metal2 s 44912 99600 44968 100000 6 reg_peri_wdata[16]
port 202 nsew signal output
rlabel metal2 s 44352 99600 44408 100000 6 reg_peri_wdata[17]
port 203 nsew signal output
rlabel metal2 s 43792 99600 43848 100000 6 reg_peri_wdata[18]
port 204 nsew signal output
rlabel metal2 s 43232 99600 43288 100000 6 reg_peri_wdata[19]
port 205 nsew signal output
rlabel metal2 s 53312 99600 53368 100000 6 reg_peri_wdata[1]
port 206 nsew signal output
rlabel metal2 s 42672 99600 42728 100000 6 reg_peri_wdata[20]
port 207 nsew signal output
rlabel metal2 s 42112 99600 42168 100000 6 reg_peri_wdata[21]
port 208 nsew signal output
rlabel metal2 s 41552 99600 41608 100000 6 reg_peri_wdata[22]
port 209 nsew signal output
rlabel metal2 s 40992 99600 41048 100000 6 reg_peri_wdata[23]
port 210 nsew signal output
rlabel metal2 s 40432 99600 40488 100000 6 reg_peri_wdata[24]
port 211 nsew signal output
rlabel metal2 s 39872 99600 39928 100000 6 reg_peri_wdata[25]
port 212 nsew signal output
rlabel metal2 s 39312 99600 39368 100000 6 reg_peri_wdata[26]
port 213 nsew signal output
rlabel metal2 s 38752 99600 38808 100000 6 reg_peri_wdata[27]
port 214 nsew signal output
rlabel metal2 s 38192 99600 38248 100000 6 reg_peri_wdata[28]
port 215 nsew signal output
rlabel metal2 s 37632 99600 37688 100000 6 reg_peri_wdata[29]
port 216 nsew signal output
rlabel metal2 s 52752 99600 52808 100000 6 reg_peri_wdata[2]
port 217 nsew signal output
rlabel metal2 s 37072 99600 37128 100000 6 reg_peri_wdata[30]
port 218 nsew signal output
rlabel metal2 s 36512 99600 36568 100000 6 reg_peri_wdata[31]
port 219 nsew signal output
rlabel metal2 s 52192 99600 52248 100000 6 reg_peri_wdata[3]
port 220 nsew signal output
rlabel metal2 s 51632 99600 51688 100000 6 reg_peri_wdata[4]
port 221 nsew signal output
rlabel metal2 s 51072 99600 51128 100000 6 reg_peri_wdata[5]
port 222 nsew signal output
rlabel metal2 s 50512 99600 50568 100000 6 reg_peri_wdata[6]
port 223 nsew signal output
rlabel metal2 s 49952 99600 50008 100000 6 reg_peri_wdata[7]
port 224 nsew signal output
rlabel metal2 s 49392 99600 49448 100000 6 reg_peri_wdata[8]
port 225 nsew signal output
rlabel metal2 s 48832 99600 48888 100000 6 reg_peri_wdata[9]
port 226 nsew signal output
rlabel metal2 s 27552 99600 27608 100000 6 reg_peri_wr
port 227 nsew signal output
rlabel metal3 s 0 95872 400 95928 6 reg_rdata[0]
port 228 nsew signal output
rlabel metal3 s 0 84672 400 84728 6 reg_rdata[10]
port 229 nsew signal output
rlabel metal3 s 0 83552 400 83608 6 reg_rdata[11]
port 230 nsew signal output
rlabel metal3 s 0 82432 400 82488 6 reg_rdata[12]
port 231 nsew signal output
rlabel metal3 s 0 81312 400 81368 6 reg_rdata[13]
port 232 nsew signal output
rlabel metal3 s 0 80192 400 80248 6 reg_rdata[14]
port 233 nsew signal output
rlabel metal3 s 0 79072 400 79128 6 reg_rdata[15]
port 234 nsew signal output
rlabel metal3 s 0 77952 400 78008 6 reg_rdata[16]
port 235 nsew signal output
rlabel metal3 s 0 76832 400 76888 6 reg_rdata[17]
port 236 nsew signal output
rlabel metal3 s 0 75712 400 75768 6 reg_rdata[18]
port 237 nsew signal output
rlabel metal3 s 0 74592 400 74648 6 reg_rdata[19]
port 238 nsew signal output
rlabel metal3 s 0 94752 400 94808 6 reg_rdata[1]
port 239 nsew signal output
rlabel metal3 s 0 73472 400 73528 6 reg_rdata[20]
port 240 nsew signal output
rlabel metal3 s 0 72352 400 72408 6 reg_rdata[21]
port 241 nsew signal output
rlabel metal3 s 0 71232 400 71288 6 reg_rdata[22]
port 242 nsew signal output
rlabel metal3 s 0 70112 400 70168 6 reg_rdata[23]
port 243 nsew signal output
rlabel metal3 s 0 68992 400 69048 6 reg_rdata[24]
port 244 nsew signal output
rlabel metal3 s 0 67872 400 67928 6 reg_rdata[25]
port 245 nsew signal output
rlabel metal3 s 0 66752 400 66808 6 reg_rdata[26]
port 246 nsew signal output
rlabel metal3 s 0 65632 400 65688 6 reg_rdata[27]
port 247 nsew signal output
rlabel metal3 s 0 64512 400 64568 6 reg_rdata[28]
port 248 nsew signal output
rlabel metal3 s 0 63392 400 63448 6 reg_rdata[29]
port 249 nsew signal output
rlabel metal3 s 0 93632 400 93688 6 reg_rdata[2]
port 250 nsew signal output
rlabel metal3 s 0 62272 400 62328 6 reg_rdata[30]
port 251 nsew signal output
rlabel metal3 s 0 61152 400 61208 6 reg_rdata[31]
port 252 nsew signal output
rlabel metal3 s 0 92512 400 92568 6 reg_rdata[3]
port 253 nsew signal output
rlabel metal3 s 0 91392 400 91448 6 reg_rdata[4]
port 254 nsew signal output
rlabel metal3 s 0 90272 400 90328 6 reg_rdata[5]
port 255 nsew signal output
rlabel metal3 s 0 89152 400 89208 6 reg_rdata[6]
port 256 nsew signal output
rlabel metal3 s 0 88032 400 88088 6 reg_rdata[7]
port 257 nsew signal output
rlabel metal3 s 0 86912 400 86968 6 reg_rdata[8]
port 258 nsew signal output
rlabel metal3 s 0 85792 400 85848 6 reg_rdata[9]
port 259 nsew signal output
rlabel metal3 s 0 60032 400 60088 6 reg_wdata[0]
port 260 nsew signal input
rlabel metal3 s 0 48832 400 48888 6 reg_wdata[10]
port 261 nsew signal input
rlabel metal3 s 0 47712 400 47768 6 reg_wdata[11]
port 262 nsew signal input
rlabel metal3 s 0 46592 400 46648 6 reg_wdata[12]
port 263 nsew signal input
rlabel metal3 s 0 45472 400 45528 6 reg_wdata[13]
port 264 nsew signal input
rlabel metal3 s 0 44352 400 44408 6 reg_wdata[14]
port 265 nsew signal input
rlabel metal3 s 0 43232 400 43288 6 reg_wdata[15]
port 266 nsew signal input
rlabel metal3 s 0 42112 400 42168 6 reg_wdata[16]
port 267 nsew signal input
rlabel metal3 s 0 40992 400 41048 6 reg_wdata[17]
port 268 nsew signal input
rlabel metal3 s 0 39872 400 39928 6 reg_wdata[18]
port 269 nsew signal input
rlabel metal3 s 0 38752 400 38808 6 reg_wdata[19]
port 270 nsew signal input
rlabel metal3 s 0 58912 400 58968 6 reg_wdata[1]
port 271 nsew signal input
rlabel metal3 s 0 37632 400 37688 6 reg_wdata[20]
port 272 nsew signal input
rlabel metal3 s 0 36512 400 36568 6 reg_wdata[21]
port 273 nsew signal input
rlabel metal3 s 0 35392 400 35448 6 reg_wdata[22]
port 274 nsew signal input
rlabel metal3 s 0 34272 400 34328 6 reg_wdata[23]
port 275 nsew signal input
rlabel metal3 s 0 33152 400 33208 6 reg_wdata[24]
port 276 nsew signal input
rlabel metal3 s 0 32032 400 32088 6 reg_wdata[25]
port 277 nsew signal input
rlabel metal3 s 0 30912 400 30968 6 reg_wdata[26]
port 278 nsew signal input
rlabel metal3 s 0 29792 400 29848 6 reg_wdata[27]
port 279 nsew signal input
rlabel metal3 s 0 28672 400 28728 6 reg_wdata[28]
port 280 nsew signal input
rlabel metal3 s 0 27552 400 27608 6 reg_wdata[29]
port 281 nsew signal input
rlabel metal3 s 0 57792 400 57848 6 reg_wdata[2]
port 282 nsew signal input
rlabel metal3 s 0 26432 400 26488 6 reg_wdata[30]
port 283 nsew signal input
rlabel metal3 s 0 25312 400 25368 6 reg_wdata[31]
port 284 nsew signal input
rlabel metal3 s 0 56672 400 56728 6 reg_wdata[3]
port 285 nsew signal input
rlabel metal3 s 0 55552 400 55608 6 reg_wdata[4]
port 286 nsew signal input
rlabel metal3 s 0 54432 400 54488 6 reg_wdata[5]
port 287 nsew signal input
rlabel metal3 s 0 53312 400 53368 6 reg_wdata[6]
port 288 nsew signal input
rlabel metal3 s 0 52192 400 52248 6 reg_wdata[7]
port 289 nsew signal input
rlabel metal3 s 0 51072 400 51128 6 reg_wdata[8]
port 290 nsew signal input
rlabel metal3 s 0 49952 400 50008 6 reg_wdata[9]
port 291 nsew signal input
rlabel metal3 s 0 7392 400 7448 6 reg_wr
port 292 nsew signal input
rlabel metal2 s 25872 99600 25928 100000 6 rtc_clk
port 293 nsew signal output
rlabel metal2 s 26432 99600 26488 100000 6 rtc_intr
port 294 nsew signal input
rlabel metal2 s 86128 0 86184 400 6 s_reset_n
port 295 nsew signal input
rlabel metal2 s 67312 0 67368 400 6 spim_miso
port 296 nsew signal input
rlabel metal2 s 69664 0 69720 400 6 spim_mosi
port 297 nsew signal output
rlabel metal2 s 55552 0 55608 400 6 spim_sck
port 298 nsew signal input
rlabel metal2 s 64960 0 65016 400 6 spim_ssn[0]
port 299 nsew signal input
rlabel metal2 s 62608 0 62664 400 6 spim_ssn[1]
port 300 nsew signal input
rlabel metal2 s 60256 0 60312 400 6 spim_ssn[2]
port 301 nsew signal input
rlabel metal2 s 57904 0 57960 400 6 spim_ssn[3]
port 302 nsew signal input
rlabel metal2 s 1456 0 1512 400 6 sspim_rst_n
port 303 nsew signal output
rlabel metal2 s 6160 0 6216 400 6 uart_rst_n[0]
port 304 nsew signal output
rlabel metal2 s 3808 0 3864 400 6 uart_rst_n[1]
port 305 nsew signal output
rlabel metal2 s 39088 0 39144 400 6 uart_rxd[0]
port 306 nsew signal output
rlabel metal2 s 34384 0 34440 400 6 uart_rxd[1]
port 307 nsew signal output
rlabel metal2 s 36736 0 36792 400 6 uart_txd[0]
port 308 nsew signal input
rlabel metal2 s 32032 0 32088 400 6 uart_txd[1]
port 309 nsew signal input
rlabel metal2 s 88480 0 88536 400 6 usb_clk
port 310 nsew signal output
rlabel metal2 s 29680 0 29736 400 6 usb_dn_i
port 311 nsew signal output
rlabel metal2 s 22624 0 22680 400 6 usb_dn_o
port 312 nsew signal input
rlabel metal2 s 27328 0 27384 400 6 usb_dp_i
port 313 nsew signal output
rlabel metal2 s 20272 0 20328 400 6 usb_dp_o
port 314 nsew signal input
rlabel metal2 s 76720 0 76776 400 6 usb_intr
port 315 nsew signal input
rlabel metal2 s 24976 0 25032 400 6 usb_oen
port 316 nsew signal input
rlabel metal2 s 10864 0 10920 400 6 usb_rst_n
port 317 nsew signal output
rlabel metal2 s 79072 0 79128 400 6 user_clock1
port 318 nsew signal input
rlabel metal2 s 81424 0 81480 400 6 user_clock2
port 319 nsew signal input
rlabel metal2 s 13216 0 13272 400 6 user_irq[0]
port 320 nsew signal output
rlabel metal2 s 15568 0 15624 400 6 user_irq[1]
port 321 nsew signal output
rlabel metal2 s 17920 0 17976 400 6 user_irq[2]
port 322 nsew signal output
rlabel metal2 s 83776 0 83832 400 6 xtal_clk
port 323 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 90000 100000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 28543122
string GDS_FILE /home/farag/carvel_riscv_soc/gf180mcu_riscv_soc/openlane/pinmux_top/runs/23_11_16_12_30/results/signoff/pinmux_top.magic.gds
string GDS_START 585258
<< end >>

