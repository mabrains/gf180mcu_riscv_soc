magic
tech gf180mcuD
magscale 1 5
timestamp 1698594342
<< obsm1 >>
rect 672 1538 19320 48246
<< metal2 >>
rect 1680 49600 1736 50000
rect 1344 0 1400 400
<< obsm2 >>
rect 854 49570 1650 49600
rect 1766 49570 19138 49600
rect 854 430 19138 49570
rect 854 400 1314 430
rect 1430 400 19138 430
<< metal3 >>
rect 0 33936 400 33992
rect 0 33600 400 33656
rect 0 33264 400 33320
rect 0 32256 400 32312
rect 0 31920 400 31976
rect 19600 31920 20000 31976
rect 0 31584 400 31640
rect 0 31248 400 31304
rect 0 29568 400 29624
rect 0 28896 400 28952
rect 0 28560 400 28616
rect 0 28224 400 28280
rect 0 27888 400 27944
rect 0 27552 400 27608
rect 0 26544 400 26600
rect 19600 26544 20000 26600
rect 0 25872 400 25928
rect 0 25536 400 25592
rect 0 25200 400 25256
rect 0 24864 400 24920
rect 19600 24864 20000 24920
rect 0 24528 400 24584
rect 0 24192 400 24248
rect 0 23856 400 23912
rect 19600 23520 20000 23576
rect 19600 23184 20000 23240
rect 0 22176 400 22232
rect 0 21840 400 21896
rect 19600 21168 20000 21224
rect 19600 20832 20000 20888
rect 0 20160 400 20216
rect 0 19824 400 19880
rect 0 19488 400 19544
rect 19600 19488 20000 19544
rect 19600 18144 20000 18200
rect 0 16464 400 16520
rect 19600 15456 20000 15512
rect 19600 15120 20000 15176
rect 19600 11424 20000 11480
<< obsm3 >>
rect 400 34022 19600 48230
rect 430 33906 19600 34022
rect 400 33686 19600 33906
rect 430 33570 19600 33686
rect 400 33350 19600 33570
rect 430 33234 19600 33350
rect 400 32342 19600 33234
rect 430 32226 19600 32342
rect 400 32006 19600 32226
rect 430 31890 19570 32006
rect 400 31670 19600 31890
rect 430 31554 19600 31670
rect 400 31334 19600 31554
rect 430 31218 19600 31334
rect 400 29654 19600 31218
rect 430 29538 19600 29654
rect 400 28982 19600 29538
rect 430 28866 19600 28982
rect 400 28646 19600 28866
rect 430 28530 19600 28646
rect 400 28310 19600 28530
rect 430 28194 19600 28310
rect 400 27974 19600 28194
rect 430 27858 19600 27974
rect 400 27638 19600 27858
rect 430 27522 19600 27638
rect 400 26630 19600 27522
rect 430 26514 19570 26630
rect 400 25958 19600 26514
rect 430 25842 19600 25958
rect 400 25622 19600 25842
rect 430 25506 19600 25622
rect 400 25286 19600 25506
rect 430 25170 19600 25286
rect 400 24950 19600 25170
rect 430 24834 19570 24950
rect 400 24614 19600 24834
rect 430 24498 19600 24614
rect 400 24278 19600 24498
rect 430 24162 19600 24278
rect 400 23942 19600 24162
rect 430 23826 19600 23942
rect 400 23606 19600 23826
rect 400 23490 19570 23606
rect 400 23270 19600 23490
rect 400 23154 19570 23270
rect 400 22262 19600 23154
rect 430 22146 19600 22262
rect 400 21926 19600 22146
rect 430 21810 19600 21926
rect 400 21254 19600 21810
rect 400 21138 19570 21254
rect 400 20918 19600 21138
rect 400 20802 19570 20918
rect 400 20246 19600 20802
rect 430 20130 19600 20246
rect 400 19910 19600 20130
rect 430 19794 19600 19910
rect 400 19574 19600 19794
rect 430 19458 19570 19574
rect 400 18230 19600 19458
rect 400 18114 19570 18230
rect 400 16550 19600 18114
rect 430 16434 19600 16550
rect 400 15542 19600 16434
rect 400 15426 19570 15542
rect 400 15206 19600 15426
rect 400 15090 19570 15206
rect 400 11510 19600 15090
rect 400 11394 19570 11510
rect 400 1554 19600 11394
<< metal4 >>
rect 2224 1538 2384 48246
rect 9904 1538 10064 48246
rect 17584 1538 17744 48246
<< obsm4 >>
rect 9310 16977 9874 31183
rect 10094 16977 17458 31183
<< labels >>
rlabel metal3 s 19600 15456 20000 15512 6 clk
port 1 nsew signal input
rlabel metal3 s 0 31920 400 31976 6 compare_in[0]
port 2 nsew signal input
rlabel metal3 s 0 24528 400 24584 6 compare_in[10]
port 3 nsew signal input
rlabel metal3 s 0 28224 400 28280 6 compare_in[11]
port 4 nsew signal input
rlabel metal3 s 0 25872 400 25928 6 compare_in[12]
port 5 nsew signal input
rlabel metal3 s 0 24192 400 24248 6 compare_in[13]
port 6 nsew signal input
rlabel metal3 s 0 27888 400 27944 6 compare_in[14]
port 7 nsew signal input
rlabel metal3 s 0 25536 400 25592 6 compare_in[15]
port 8 nsew signal input
rlabel metal3 s 0 25200 400 25256 6 compare_in[16]
port 9 nsew signal input
rlabel metal3 s 0 24864 400 24920 6 compare_in[17]
port 10 nsew signal input
rlabel metal3 s 0 22176 400 22232 6 compare_in[18]
port 11 nsew signal input
rlabel metal3 s 0 23856 400 23912 6 compare_in[19]
port 12 nsew signal input
rlabel metal3 s 0 33264 400 33320 6 compare_in[1]
port 13 nsew signal input
rlabel metal3 s 0 19488 400 19544 6 compare_in[20]
port 14 nsew signal input
rlabel metal3 s 0 19824 400 19880 6 compare_in[21]
port 15 nsew signal input
rlabel metal3 s 0 20160 400 20216 6 compare_in[22]
port 16 nsew signal input
rlabel metal3 s 0 21840 400 21896 6 compare_in[23]
port 17 nsew signal input
rlabel metal3 s 0 33936 400 33992 6 compare_in[2]
port 18 nsew signal input
rlabel metal3 s 0 33600 400 33656 6 compare_in[3]
port 19 nsew signal input
rlabel metal3 s 0 32256 400 32312 6 compare_in[4]
port 20 nsew signal input
rlabel metal3 s 0 31248 400 31304 6 compare_in[5]
port 21 nsew signal input
rlabel metal3 s 0 31584 400 31640 6 compare_in[6]
port 22 nsew signal input
rlabel metal3 s 0 29568 400 29624 6 compare_in[7]
port 23 nsew signal input
rlabel metal3 s 0 28560 400 28616 6 compare_in[8]
port 24 nsew signal input
rlabel metal3 s 0 28896 400 28952 6 compare_in[9]
port 25 nsew signal input
rlabel metal3 s 19600 15120 20000 15176 6 io_oeb[0]
port 26 nsew signal output
rlabel metal2 s 1344 0 1400 400 6 io_oeb[1]
port 27 nsew signal output
rlabel metal3 s 19600 31920 20000 31976 6 io_oeb[2]
port 28 nsew signal output
rlabel metal3 s 19600 18144 20000 18200 6 io_oeb[3]
port 29 nsew signal output
rlabel metal3 s 19600 11424 20000 11480 6 io_oeb[4]
port 30 nsew signal output
rlabel metal2 s 1680 49600 1736 50000 6 io_oeb[5]
port 31 nsew signal output
rlabel metal3 s 0 16464 400 16520 6 io_oeb[6]
port 32 nsew signal output
rlabel metal3 s 19600 19488 20000 19544 6 led_out[0]
port 33 nsew signal output
rlabel metal3 s 19600 26544 20000 26600 6 led_out[1]
port 34 nsew signal output
rlabel metal3 s 19600 20832 20000 20888 6 led_out[2]
port 35 nsew signal output
rlabel metal3 s 19600 21168 20000 21224 6 led_out[3]
port 36 nsew signal output
rlabel metal3 s 19600 23184 20000 23240 6 led_out[4]
port 37 nsew signal output
rlabel metal3 s 19600 23520 20000 23576 6 led_out[5]
port 38 nsew signal output
rlabel metal3 s 19600 24864 20000 24920 6 led_out[6]
port 39 nsew signal output
rlabel metal3 s 0 27552 400 27608 6 reset
port 40 nsew signal input
rlabel metal3 s 0 26544 400 26600 6 update_compare
port 41 nsew signal input
rlabel metal4 s 2224 1538 2384 48246 6 vdd
port 42 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 48246 6 vdd
port 42 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 48246 6 vss
port 43 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 20000 50000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1337790
string GDS_FILE /home/farag/carvel_riscv_soc/gf180mcu_riscv_soc/openlane/riscv_top/runs/23_10_29_17_42/results/signoff/riscv_top.magic.gds
string GDS_START 336542
<< end >>

