VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO serv_rf_top
  CLASS BLOCK ;
  FOREIGN serv_rf_top ;
  ORIGIN 0.000 0.000 ;
  SIZE 755.700 BY 773.620 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 756.860 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 756.860 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 15.380 331.040 756.860 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 483.040 15.380 484.640 756.860 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 636.640 15.380 638.240 756.860 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 756.860 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 756.860 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 406.240 15.380 407.840 756.860 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 559.840 15.380 561.440 756.860 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 713.440 15.380 715.040 756.860 ;
    END
  END VSS
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.738000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 554.400 755.700 554.960 ;
    END
  END clk
  PIN i_dbus_ack
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 147.840 755.700 148.400 ;
    END
  END i_dbus_ack
  PIN i_dbus_rdt[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 131.040 755.700 131.600 ;
    END
  END i_dbus_rdt[0]
  PIN i_dbus_rdt[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 551.040 755.700 551.600 ;
    END
  END i_dbus_rdt[10]
  PIN i_dbus_rdt[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 473.760 755.700 474.320 ;
    END
  END i_dbus_rdt[11]
  PIN i_dbus_rdt[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 504.000 755.700 504.560 ;
    END
  END i_dbus_rdt[12]
  PIN i_dbus_rdt[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 436.800 755.700 437.360 ;
    END
  END i_dbus_rdt[13]
  PIN i_dbus_rdt[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 426.720 755.700 427.280 ;
    END
  END i_dbus_rdt[14]
  PIN i_dbus_rdt[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 352.800 755.700 353.360 ;
    END
  END i_dbus_rdt[15]
  PIN i_dbus_rdt[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 403.200 755.700 403.760 ;
    END
  END i_dbus_rdt[16]
  PIN i_dbus_rdt[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 396.480 755.700 397.040 ;
    END
  END i_dbus_rdt[17]
  PIN i_dbus_rdt[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 430.080 755.700 430.640 ;
    END
  END i_dbus_rdt[18]
  PIN i_dbus_rdt[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 477.120 755.700 477.680 ;
    END
  END i_dbus_rdt[19]
  PIN i_dbus_rdt[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 258.720 755.700 259.280 ;
    END
  END i_dbus_rdt[1]
  PIN i_dbus_rdt[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 547.680 755.700 548.240 ;
    END
  END i_dbus_rdt[20]
  PIN i_dbus_rdt[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 416.640 755.700 417.200 ;
    END
  END i_dbus_rdt[21]
  PIN i_dbus_rdt[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 453.600 755.700 454.160 ;
    END
  END i_dbus_rdt[22]
  PIN i_dbus_rdt[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 342.720 755.700 343.280 ;
    END
  END i_dbus_rdt[23]
  PIN i_dbus_rdt[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 510.720 755.700 511.280 ;
    END
  END i_dbus_rdt[24]
  PIN i_dbus_rdt[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 356.160 755.700 356.720 ;
    END
  END i_dbus_rdt[25]
  PIN i_dbus_rdt[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 514.080 755.700 514.640 ;
    END
  END i_dbus_rdt[26]
  PIN i_dbus_rdt[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 383.040 755.700 383.600 ;
    END
  END i_dbus_rdt[27]
  PIN i_dbus_rdt[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 295.680 755.700 296.240 ;
    END
  END i_dbus_rdt[28]
  PIN i_dbus_rdt[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 544.320 755.700 544.880 ;
    END
  END i_dbus_rdt[29]
  PIN i_dbus_rdt[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 120.960 755.700 121.520 ;
    END
  END i_dbus_rdt[2]
  PIN i_dbus_rdt[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 524.160 755.700 524.720 ;
    END
  END i_dbus_rdt[30]
  PIN i_dbus_rdt[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 292.320 755.700 292.880 ;
    END
  END i_dbus_rdt[31]
  PIN i_dbus_rdt[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 238.560 755.700 239.120 ;
    END
  END i_dbus_rdt[3]
  PIN i_dbus_rdt[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 228.480 755.700 229.040 ;
    END
  END i_dbus_rdt[4]
  PIN i_dbus_rdt[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 225.120 755.700 225.680 ;
    END
  END i_dbus_rdt[5]
  PIN i_dbus_rdt[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 520.800 755.700 521.360 ;
    END
  END i_dbus_rdt[6]
  PIN i_dbus_rdt[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 336.000 755.700 336.560 ;
    END
  END i_dbus_rdt[7]
  PIN i_dbus_rdt[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 312.480 755.700 313.040 ;
    END
  END i_dbus_rdt[8]
  PIN i_dbus_rdt[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 346.080 755.700 346.640 ;
    END
  END i_dbus_rdt[9]
  PIN i_ext_rd[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 0.000 0.560 4.000 ;
    END
  END i_ext_rd[0]
  PIN i_ext_rd[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3.360 0.000 3.920 4.000 ;
    END
  END i_ext_rd[10]
  PIN i_ext_rd[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 6.720 0.000 7.280 4.000 ;
    END
  END i_ext_rd[11]
  PIN i_ext_rd[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 10.080 0.000 10.640 4.000 ;
    END
  END i_ext_rd[12]
  PIN i_ext_rd[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 13.440 0.000 14.000 4.000 ;
    END
  END i_ext_rd[13]
  PIN i_ext_rd[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 16.800 0.000 17.360 4.000 ;
    END
  END i_ext_rd[14]
  PIN i_ext_rd[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 20.160 0.000 20.720 4.000 ;
    END
  END i_ext_rd[15]
  PIN i_ext_rd[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 23.520 0.000 24.080 4.000 ;
    END
  END i_ext_rd[16]
  PIN i_ext_rd[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 26.880 0.000 27.440 4.000 ;
    END
  END i_ext_rd[17]
  PIN i_ext_rd[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 30.240 0.000 30.800 4.000 ;
    END
  END i_ext_rd[18]
  PIN i_ext_rd[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 33.600 0.000 34.160 4.000 ;
    END
  END i_ext_rd[19]
  PIN i_ext_rd[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 36.960 0.000 37.520 4.000 ;
    END
  END i_ext_rd[1]
  PIN i_ext_rd[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 40.320 0.000 40.880 4.000 ;
    END
  END i_ext_rd[20]
  PIN i_ext_rd[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 43.680 0.000 44.240 4.000 ;
    END
  END i_ext_rd[21]
  PIN i_ext_rd[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 47.040 0.000 47.600 4.000 ;
    END
  END i_ext_rd[22]
  PIN i_ext_rd[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 50.400 0.000 50.960 4.000 ;
    END
  END i_ext_rd[23]
  PIN i_ext_rd[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 53.760 0.000 54.320 4.000 ;
    END
  END i_ext_rd[24]
  PIN i_ext_rd[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 57.120 0.000 57.680 4.000 ;
    END
  END i_ext_rd[25]
  PIN i_ext_rd[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 60.480 0.000 61.040 4.000 ;
    END
  END i_ext_rd[26]
  PIN i_ext_rd[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 63.840 0.000 64.400 4.000 ;
    END
  END i_ext_rd[27]
  PIN i_ext_rd[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 67.200 0.000 67.760 4.000 ;
    END
  END i_ext_rd[28]
  PIN i_ext_rd[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 70.560 0.000 71.120 4.000 ;
    END
  END i_ext_rd[29]
  PIN i_ext_rd[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 73.920 0.000 74.480 4.000 ;
    END
  END i_ext_rd[2]
  PIN i_ext_rd[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 77.280 0.000 77.840 4.000 ;
    END
  END i_ext_rd[30]
  PIN i_ext_rd[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 80.640 0.000 81.200 4.000 ;
    END
  END i_ext_rd[31]
  PIN i_ext_rd[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 84.000 0.000 84.560 4.000 ;
    END
  END i_ext_rd[3]
  PIN i_ext_rd[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 87.360 0.000 87.920 4.000 ;
    END
  END i_ext_rd[4]
  PIN i_ext_rd[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 90.720 0.000 91.280 4.000 ;
    END
  END i_ext_rd[5]
  PIN i_ext_rd[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 94.080 0.000 94.640 4.000 ;
    END
  END i_ext_rd[6]
  PIN i_ext_rd[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 97.440 0.000 98.000 4.000 ;
    END
  END i_ext_rd[7]
  PIN i_ext_rd[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 100.800 0.000 101.360 4.000 ;
    END
  END i_ext_rd[8]
  PIN i_ext_rd[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 104.160 0.000 104.720 4.000 ;
    END
  END i_ext_rd[9]
  PIN i_ext_ready
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 107.520 0.000 108.080 4.000 ;
    END
  END i_ext_ready
  PIN i_ibus_ack
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 181.440 755.700 182.000 ;
    END
  END i_ibus_ack
  PIN i_ibus_rdt[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 110.880 0.000 111.440 4.000 ;
    END
  END i_ibus_rdt[0]
  PIN i_ibus_rdt[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 208.320 755.700 208.880 ;
    END
  END i_ibus_rdt[10]
  PIN i_ibus_rdt[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 191.520 755.700 192.080 ;
    END
  END i_ibus_rdt[11]
  PIN i_ibus_rdt[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 278.880 755.700 279.440 ;
    END
  END i_ibus_rdt[12]
  PIN i_ibus_rdt[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 268.800 755.700 269.360 ;
    END
  END i_ibus_rdt[13]
  PIN i_ibus_rdt[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 262.080 755.700 262.640 ;
    END
  END i_ibus_rdt[14]
  PIN i_ibus_rdt[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 285.600 755.700 286.160 ;
    END
  END i_ibus_rdt[15]
  PIN i_ibus_rdt[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 325.920 755.700 326.480 ;
    END
  END i_ibus_rdt[16]
  PIN i_ibus_rdt[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 255.360 755.700 255.920 ;
    END
  END i_ibus_rdt[17]
  PIN i_ibus_rdt[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 124.320 755.700 124.880 ;
    END
  END i_ibus_rdt[18]
  PIN i_ibus_rdt[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 134.400 755.700 134.960 ;
    END
  END i_ibus_rdt[19]
  PIN i_ibus_rdt[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 114.240 0.000 114.800 4.000 ;
    END
  END i_ibus_rdt[1]
  PIN i_ibus_rdt[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 688.800 0.000 689.360 4.000 ;
    END
  END i_ibus_rdt[20]
  PIN i_ibus_rdt[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 194.880 755.700 195.440 ;
    END
  END i_ibus_rdt[21]
  PIN i_ibus_rdt[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 745.920 0.000 746.480 4.000 ;
    END
  END i_ibus_rdt[22]
  PIN i_ibus_rdt[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 161.280 755.700 161.840 ;
    END
  END i_ibus_rdt[23]
  PIN i_ibus_rdt[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 171.360 755.700 171.920 ;
    END
  END i_ibus_rdt[24]
  PIN i_ibus_rdt[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 749.280 0.000 749.840 4.000 ;
    END
  END i_ibus_rdt[25]
  PIN i_ibus_rdt[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 678.720 0.000 679.280 4.000 ;
    END
  END i_ibus_rdt[26]
  PIN i_ibus_rdt[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 729.120 0.000 729.680 4.000 ;
    END
  END i_ibus_rdt[27]
  PIN i_ibus_rdt[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 735.840 0.000 736.400 4.000 ;
    END
  END i_ibus_rdt[28]
  PIN i_ibus_rdt[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 739.200 0.000 739.760 4.000 ;
    END
  END i_ibus_rdt[29]
  PIN i_ibus_rdt[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 685.440 0.000 686.000 4.000 ;
    END
  END i_ibus_rdt[2]
  PIN i_ibus_rdt[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 732.480 0.000 733.040 4.000 ;
    END
  END i_ibus_rdt[30]
  PIN i_ibus_rdt[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 164.640 755.700 165.200 ;
    END
  END i_ibus_rdt[31]
  PIN i_ibus_rdt[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 288.960 755.700 289.520 ;
    END
  END i_ibus_rdt[3]
  PIN i_ibus_rdt[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 218.400 755.700 218.960 ;
    END
  END i_ibus_rdt[4]
  PIN i_ibus_rdt[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 188.160 755.700 188.720 ;
    END
  END i_ibus_rdt[5]
  PIN i_ibus_rdt[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 231.840 755.700 232.400 ;
    END
  END i_ibus_rdt[6]
  PIN i_ibus_rdt[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 201.600 755.700 202.160 ;
    END
  END i_ibus_rdt[7]
  PIN i_ibus_rdt[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 198.240 755.700 198.800 ;
    END
  END i_ibus_rdt[8]
  PIN i_ibus_rdt[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 211.680 755.700 212.240 ;
    END
  END i_ibus_rdt[9]
  PIN i_rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 752.640 0.000 753.200 4.000 ;
    END
  END i_rst
  PIN i_timer_irq
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 712.320 0.000 712.880 4.000 ;
    END
  END i_timer_irq
  PIN o_dbus_adr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 305.760 4.000 306.320 ;
    END
  END o_dbus_adr[0]
  PIN o_dbus_adr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 722.400 0.000 722.960 4.000 ;
    END
  END o_dbus_adr[10]
  PIN o_dbus_adr[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 698.880 0.000 699.440 4.000 ;
    END
  END o_dbus_adr[11]
  PIN o_dbus_adr[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 719.040 0.000 719.600 4.000 ;
    END
  END o_dbus_adr[12]
  PIN o_dbus_adr[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 695.520 0.000 696.080 4.000 ;
    END
  END o_dbus_adr[13]
  PIN o_dbus_adr[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 708.960 0.000 709.520 4.000 ;
    END
  END o_dbus_adr[14]
  PIN o_dbus_adr[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 705.600 0.000 706.160 4.000 ;
    END
  END o_dbus_adr[15]
  PIN o_dbus_adr[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 692.160 0.000 692.720 4.000 ;
    END
  END o_dbus_adr[16]
  PIN o_dbus_adr[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 715.680 0.000 716.240 4.000 ;
    END
  END o_dbus_adr[17]
  PIN o_dbus_adr[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 725.760 0.000 726.320 4.000 ;
    END
  END o_dbus_adr[18]
  PIN o_dbus_adr[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 702.240 0.000 702.800 4.000 ;
    END
  END o_dbus_adr[19]
  PIN o_dbus_adr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 446.880 755.700 447.440 ;
    END
  END o_dbus_adr[1]
  PIN o_dbus_adr[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 682.080 0.000 682.640 4.000 ;
    END
  END o_dbus_adr[20]
  PIN o_dbus_adr[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 742.560 0.000 743.120 4.000 ;
    END
  END o_dbus_adr[21]
  PIN o_dbus_adr[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 524.160 0.000 524.720 4.000 ;
    END
  END o_dbus_adr[22]
  PIN o_dbus_adr[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 500.640 0.000 501.200 4.000 ;
    END
  END o_dbus_adr[23]
  PIN o_dbus_adr[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 504.000 0.000 504.560 4.000 ;
    END
  END o_dbus_adr[24]
  PIN o_dbus_adr[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 517.440 0.000 518.000 4.000 ;
    END
  END o_dbus_adr[25]
  PIN o_dbus_adr[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 672.000 0.000 672.560 4.000 ;
    END
  END o_dbus_adr[26]
  PIN o_dbus_adr[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 675.360 0.000 675.920 4.000 ;
    END
  END o_dbus_adr[27]
  PIN o_dbus_adr[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 551.040 0.000 551.600 4.000 ;
    END
  END o_dbus_adr[28]
  PIN o_dbus_adr[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 567.840 0.000 568.400 4.000 ;
    END
  END o_dbus_adr[29]
  PIN o_dbus_adr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 0.000 755.700 0.560 ;
    END
  END o_dbus_adr[2]
  PIN o_dbus_adr[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 574.560 0.000 575.120 4.000 ;
    END
  END o_dbus_adr[30]
  PIN o_dbus_adr[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 588.000 0.000 588.560 4.000 ;
    END
  END o_dbus_adr[31]
  PIN o_dbus_adr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 13.440 755.700 14.000 ;
    END
  END o_dbus_adr[3]
  PIN o_dbus_adr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 618.240 0.000 618.800 4.000 ;
    END
  END o_dbus_adr[4]
  PIN o_dbus_adr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 598.080 0.000 598.640 4.000 ;
    END
  END o_dbus_adr[5]
  PIN o_dbus_adr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 611.520 0.000 612.080 4.000 ;
    END
  END o_dbus_adr[6]
  PIN o_dbus_adr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 638.400 0.000 638.960 4.000 ;
    END
  END o_dbus_adr[7]
  PIN o_dbus_adr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 635.040 0.000 635.600 4.000 ;
    END
  END o_dbus_adr[8]
  PIN o_dbus_adr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 621.600 0.000 622.160 4.000 ;
    END
  END o_dbus_adr[9]
  PIN o_dbus_cyc
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 204.960 755.700 205.520 ;
    END
  END o_dbus_cyc
  PIN o_dbus_dat[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 137.760 755.700 138.320 ;
    END
  END o_dbus_dat[0]
  PIN o_dbus_dat[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 480.480 755.700 481.040 ;
    END
  END o_dbus_dat[10]
  PIN o_dbus_dat[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 322.560 755.700 323.120 ;
    END
  END o_dbus_dat[11]
  PIN o_dbus_dat[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 393.120 755.700 393.680 ;
    END
  END o_dbus_dat[12]
  PIN o_dbus_dat[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 359.520 755.700 360.080 ;
    END
  END o_dbus_dat[13]
  PIN o_dbus_dat[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 409.920 755.700 410.480 ;
    END
  END o_dbus_dat[14]
  PIN o_dbus_dat[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 470.400 755.700 470.960 ;
    END
  END o_dbus_dat[15]
  PIN o_dbus_dat[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 487.200 755.700 487.760 ;
    END
  END o_dbus_dat[16]
  PIN o_dbus_dat[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 386.400 755.700 386.960 ;
    END
  END o_dbus_dat[17]
  PIN o_dbus_dat[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 467.040 755.700 467.600 ;
    END
  END o_dbus_dat[18]
  PIN o_dbus_dat[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 420.000 755.700 420.560 ;
    END
  END o_dbus_dat[19]
  PIN o_dbus_dat[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 275.520 755.700 276.080 ;
    END
  END o_dbus_dat[1]
  PIN o_dbus_dat[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 369.600 755.700 370.160 ;
    END
  END o_dbus_dat[20]
  PIN o_dbus_dat[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 379.680 755.700 380.240 ;
    END
  END o_dbus_dat[21]
  PIN o_dbus_dat[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 349.440 755.700 350.000 ;
    END
  END o_dbus_dat[22]
  PIN o_dbus_dat[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 362.880 755.700 363.440 ;
    END
  END o_dbus_dat[23]
  PIN o_dbus_dat[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 433.440 755.700 434.000 ;
    END
  END o_dbus_dat[24]
  PIN o_dbus_dat[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 376.320 755.700 376.880 ;
    END
  END o_dbus_dat[25]
  PIN o_dbus_dat[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 389.760 755.700 390.320 ;
    END
  END o_dbus_dat[26]
  PIN o_dbus_dat[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 329.280 755.700 329.840 ;
    END
  END o_dbus_dat[27]
  PIN o_dbus_dat[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 537.600 755.700 538.160 ;
    END
  END o_dbus_dat[28]
  PIN o_dbus_dat[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 413.280 755.700 413.840 ;
    END
  END o_dbus_dat[29]
  PIN o_dbus_dat[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 144.480 755.700 145.040 ;
    END
  END o_dbus_dat[2]
  PIN o_dbus_dat[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 315.840 755.700 316.400 ;
    END
  END o_dbus_dat[30]
  PIN o_dbus_dat[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 302.400 755.700 302.960 ;
    END
  END o_dbus_dat[31]
  PIN o_dbus_dat[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 235.200 755.700 235.760 ;
    END
  END o_dbus_dat[3]
  PIN o_dbus_dat[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 174.720 755.700 175.280 ;
    END
  END o_dbus_dat[4]
  PIN o_dbus_dat[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 215.040 755.700 215.600 ;
    END
  END o_dbus_dat[5]
  PIN o_dbus_dat[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 221.760 755.700 222.320 ;
    END
  END o_dbus_dat[6]
  PIN o_dbus_dat[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 319.200 755.700 319.760 ;
    END
  END o_dbus_dat[7]
  PIN o_dbus_dat[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 507.360 755.700 507.920 ;
    END
  END o_dbus_dat[8]
  PIN o_dbus_dat[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 332.640 755.700 333.200 ;
    END
  END o_dbus_dat[9]
  PIN o_dbus_sel[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 141.120 755.700 141.680 ;
    END
  END o_dbus_sel[0]
  PIN o_dbus_sel[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 245.280 755.700 245.840 ;
    END
  END o_dbus_sel[1]
  PIN o_dbus_sel[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 157.920 755.700 158.480 ;
    END
  END o_dbus_sel[2]
  PIN o_dbus_sel[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 154.560 755.700 155.120 ;
    END
  END o_dbus_sel[3]
  PIN o_dbus_we
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 184.800 755.700 185.360 ;
    END
  END o_dbus_we
  PIN o_ext_funct3[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 252.000 755.700 252.560 ;
    END
  END o_ext_funct3[0]
  PIN o_ext_funct3[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 241.920 755.700 242.480 ;
    END
  END o_ext_funct3[1]
  PIN o_ext_funct3[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 248.640 755.700 249.200 ;
    END
  END o_ext_funct3[2]
  PIN o_ext_rs1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 114.240 755.700 114.800 ;
    END
  END o_ext_rs1[0]
  PIN o_ext_rs1[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 604.800 0.000 605.360 4.000 ;
    END
  END o_ext_rs1[10]
  PIN o_ext_rs1[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 591.360 0.000 591.920 4.000 ;
    END
  END o_ext_rs1[11]
  PIN o_ext_rs1[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 577.920 0.000 578.480 4.000 ;
    END
  END o_ext_rs1[12]
  PIN o_ext_rs1[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 584.640 0.000 585.200 4.000 ;
    END
  END o_ext_rs1[13]
  PIN o_ext_rs1[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 571.200 0.000 571.760 4.000 ;
    END
  END o_ext_rs1[14]
  PIN o_ext_rs1[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 561.120 0.000 561.680 4.000 ;
    END
  END o_ext_rs1[15]
  PIN o_ext_rs1[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 554.400 0.000 554.960 4.000 ;
    END
  END o_ext_rs1[16]
  PIN o_ext_rs1[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 544.320 0.000 544.880 4.000 ;
    END
  END o_ext_rs1[17]
  PIN o_ext_rs1[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 527.520 0.000 528.080 4.000 ;
    END
  END o_ext_rs1[18]
  PIN o_ext_rs1[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 534.240 0.000 534.800 4.000 ;
    END
  END o_ext_rs1[19]
  PIN o_ext_rs1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 110.880 755.700 111.440 ;
    END
  END o_ext_rs1[1]
  PIN o_ext_rs1[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 540.960 0.000 541.520 4.000 ;
    END
  END o_ext_rs1[20]
  PIN o_ext_rs1[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 537.600 0.000 538.160 4.000 ;
    END
  END o_ext_rs1[21]
  PIN o_ext_rs1[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 520.800 0.000 521.360 4.000 ;
    END
  END o_ext_rs1[22]
  PIN o_ext_rs1[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 510.720 0.000 511.280 4.000 ;
    END
  END o_ext_rs1[23]
  PIN o_ext_rs1[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 507.360 0.000 507.920 4.000 ;
    END
  END o_ext_rs1[24]
  PIN o_ext_rs1[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 514.080 0.000 514.640 4.000 ;
    END
  END o_ext_rs1[25]
  PIN o_ext_rs1[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 530.880 0.000 531.440 4.000 ;
    END
  END o_ext_rs1[26]
  PIN o_ext_rs1[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 547.680 0.000 548.240 4.000 ;
    END
  END o_ext_rs1[27]
  PIN o_ext_rs1[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 557.760 0.000 558.320 4.000 ;
    END
  END o_ext_rs1[28]
  PIN o_ext_rs1[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 564.480 0.000 565.040 4.000 ;
    END
  END o_ext_rs1[29]
  PIN o_ext_rs1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 6.720 755.700 7.280 ;
    END
  END o_ext_rs1[2]
  PIN o_ext_rs1[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 581.280 0.000 581.840 4.000 ;
    END
  END o_ext_rs1[30]
  PIN o_ext_rs1[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 594.720 0.000 595.280 4.000 ;
    END
  END o_ext_rs1[31]
  PIN o_ext_rs1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 80.640 755.700 81.200 ;
    END
  END o_ext_rs1[3]
  PIN o_ext_rs1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 614.880 0.000 615.440 4.000 ;
    END
  END o_ext_rs1[4]
  PIN o_ext_rs1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 601.440 0.000 602.000 4.000 ;
    END
  END o_ext_rs1[5]
  PIN o_ext_rs1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 608.160 0.000 608.720 4.000 ;
    END
  END o_ext_rs1[6]
  PIN o_ext_rs1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 628.320 0.000 628.880 4.000 ;
    END
  END o_ext_rs1[7]
  PIN o_ext_rs1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 631.680 0.000 632.240 4.000 ;
    END
  END o_ext_rs1[8]
  PIN o_ext_rs1[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 624.960 0.000 625.520 4.000 ;
    END
  END o_ext_rs1[9]
  PIN o_ext_rs2[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 127.680 755.700 128.240 ;
    END
  END o_ext_rs2[0]
  PIN o_ext_rs2[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 339.360 755.700 339.920 ;
    END
  END o_ext_rs2[10]
  PIN o_ext_rs2[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 500.640 755.700 501.200 ;
    END
  END o_ext_rs2[11]
  PIN o_ext_rs2[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 406.560 755.700 407.120 ;
    END
  END o_ext_rs2[12]
  PIN o_ext_rs2[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 366.240 755.700 366.800 ;
    END
  END o_ext_rs2[13]
  PIN o_ext_rs2[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 450.240 755.700 450.800 ;
    END
  END o_ext_rs2[14]
  PIN o_ext_rs2[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 456.960 755.700 457.520 ;
    END
  END o_ext_rs2[15]
  PIN o_ext_rs2[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 265.440 755.700 266.000 ;
    END
  END o_ext_rs2[16]
  PIN o_ext_rs2[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 463.680 755.700 464.240 ;
    END
  END o_ext_rs2[17]
  PIN o_ext_rs2[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 493.920 755.700 494.480 ;
    END
  END o_ext_rs2[18]
  PIN o_ext_rs2[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 423.360 755.700 423.920 ;
    END
  END o_ext_rs2[19]
  PIN o_ext_rs2[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 272.160 755.700 272.720 ;
    END
  END o_ext_rs2[1]
  PIN o_ext_rs2[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 399.840 755.700 400.400 ;
    END
  END o_ext_rs2[20]
  PIN o_ext_rs2[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 517.440 755.700 518.000 ;
    END
  END o_ext_rs2[21]
  PIN o_ext_rs2[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 440.160 755.700 440.720 ;
    END
  END o_ext_rs2[22]
  PIN o_ext_rs2[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 443.520 755.700 444.080 ;
    END
  END o_ext_rs2[23]
  PIN o_ext_rs2[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 490.560 755.700 491.120 ;
    END
  END o_ext_rs2[24]
  PIN o_ext_rs2[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 460.320 755.700 460.880 ;
    END
  END o_ext_rs2[25]
  PIN o_ext_rs2[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 530.880 755.700 531.440 ;
    END
  END o_ext_rs2[26]
  PIN o_ext_rs2[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 540.960 755.700 541.520 ;
    END
  END o_ext_rs2[27]
  PIN o_ext_rs2[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 527.520 755.700 528.080 ;
    END
  END o_ext_rs2[28]
  PIN o_ext_rs2[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 282.240 755.700 282.800 ;
    END
  END o_ext_rs2[29]
  PIN o_ext_rs2[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 497.280 755.700 497.840 ;
    END
  END o_ext_rs2[2]
  PIN o_ext_rs2[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 372.960 755.700 373.520 ;
    END
  END o_ext_rs2[30]
  PIN o_ext_rs2[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 534.240 755.700 534.800 ;
    END
  END o_ext_rs2[31]
  PIN o_ext_rs2[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 151.200 755.700 151.760 ;
    END
  END o_ext_rs2[3]
  PIN o_ext_rs2[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 168.000 755.700 168.560 ;
    END
  END o_ext_rs2[4]
  PIN o_ext_rs2[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 178.080 755.700 178.640 ;
    END
  END o_ext_rs2[5]
  PIN o_ext_rs2[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 305.760 755.700 306.320 ;
    END
  END o_ext_rs2[6]
  PIN o_ext_rs2[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 483.840 755.700 484.400 ;
    END
  END o_ext_rs2[7]
  PIN o_ext_rs2[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 299.040 755.700 299.600 ;
    END
  END o_ext_rs2[8]
  PIN o_ext_rs2[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 309.120 755.700 309.680 ;
    END
  END o_ext_rs2[9]
  PIN o_ibus_adr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 94.080 755.700 94.640 ;
    END
  END o_ibus_adr[0]
  PIN o_ibus_adr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 23.520 755.700 24.080 ;
    END
  END o_ibus_adr[10]
  PIN o_ibus_adr[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 26.880 755.700 27.440 ;
    END
  END o_ibus_adr[11]
  PIN o_ibus_adr[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 30.240 755.700 30.800 ;
    END
  END o_ibus_adr[12]
  PIN o_ibus_adr[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 33.600 755.700 34.160 ;
    END
  END o_ibus_adr[13]
  PIN o_ibus_adr[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 36.960 755.700 37.520 ;
    END
  END o_ibus_adr[14]
  PIN o_ibus_adr[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 40.320 755.700 40.880 ;
    END
  END o_ibus_adr[15]
  PIN o_ibus_adr[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 47.040 755.700 47.600 ;
    END
  END o_ibus_adr[16]
  PIN o_ibus_adr[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 53.760 755.700 54.320 ;
    END
  END o_ibus_adr[17]
  PIN o_ibus_adr[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 63.840 755.700 64.400 ;
    END
  END o_ibus_adr[18]
  PIN o_ibus_adr[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 73.920 755.700 74.480 ;
    END
  END o_ibus_adr[19]
  PIN o_ibus_adr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 77.280 755.700 77.840 ;
    END
  END o_ibus_adr[1]
  PIN o_ibus_adr[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 20.160 755.700 20.720 ;
    END
  END o_ibus_adr[20]
  PIN o_ibus_adr[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 70.560 755.700 71.120 ;
    END
  END o_ibus_adr[21]
  PIN o_ibus_adr[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 16.800 755.700 17.360 ;
    END
  END o_ibus_adr[22]
  PIN o_ibus_adr[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 84.000 755.700 84.560 ;
    END
  END o_ibus_adr[23]
  PIN o_ibus_adr[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 97.440 755.700 98.000 ;
    END
  END o_ibus_adr[24]
  PIN o_ibus_adr[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 3.360 755.700 3.920 ;
    END
  END o_ibus_adr[25]
  PIN o_ibus_adr[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 107.520 755.700 108.080 ;
    END
  END o_ibus_adr[26]
  PIN o_ibus_adr[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 104.160 755.700 104.720 ;
    END
  END o_ibus_adr[27]
  PIN o_ibus_adr[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 100.800 755.700 101.360 ;
    END
  END o_ibus_adr[28]
  PIN o_ibus_adr[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 10.080 755.700 10.640 ;
    END
  END o_ibus_adr[29]
  PIN o_ibus_adr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 67.200 755.700 67.760 ;
    END
  END o_ibus_adr[2]
  PIN o_ibus_adr[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 90.720 755.700 91.280 ;
    END
  END o_ibus_adr[30]
  PIN o_ibus_adr[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 87.360 755.700 87.920 ;
    END
  END o_ibus_adr[31]
  PIN o_ibus_adr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 57.120 755.700 57.680 ;
    END
  END o_ibus_adr[3]
  PIN o_ibus_adr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 648.480 0.000 649.040 4.000 ;
    END
  END o_ibus_adr[4]
  PIN o_ibus_adr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 651.840 0.000 652.400 4.000 ;
    END
  END o_ibus_adr[5]
  PIN o_ibus_adr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 655.200 0.000 655.760 4.000 ;
    END
  END o_ibus_adr[6]
  PIN o_ibus_adr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 43.680 755.700 44.240 ;
    END
  END o_ibus_adr[7]
  PIN o_ibus_adr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 50.400 755.700 50.960 ;
    END
  END o_ibus_adr[8]
  PIN o_ibus_adr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 60.480 755.700 61.040 ;
    END
  END o_ibus_adr[9]
  PIN o_ibus_cyc
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 751.700 117.600 755.700 118.160 ;
    END
  END o_ibus_cyc
  PIN o_mdu_valid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 571.200 769.620 571.760 773.620 ;
    END
  END o_mdu_valid
  OBS
      LAYER Metal1 ;
        RECT 6.720 4.630 748.720 756.860 ;
      LAYER Metal2 ;
        RECT 8.540 769.320 570.900 769.620 ;
        RECT 572.060 769.320 753.060 769.620 ;
        RECT 8.540 4.300 753.060 769.320 ;
        RECT 8.540 0.090 9.780 4.300 ;
        RECT 10.940 0.090 13.140 4.300 ;
        RECT 14.300 0.090 16.500 4.300 ;
        RECT 17.660 0.090 19.860 4.300 ;
        RECT 21.020 0.090 23.220 4.300 ;
        RECT 24.380 0.090 26.580 4.300 ;
        RECT 27.740 0.090 29.940 4.300 ;
        RECT 31.100 0.090 33.300 4.300 ;
        RECT 34.460 0.090 36.660 4.300 ;
        RECT 37.820 0.090 40.020 4.300 ;
        RECT 41.180 0.090 43.380 4.300 ;
        RECT 44.540 0.090 46.740 4.300 ;
        RECT 47.900 0.090 50.100 4.300 ;
        RECT 51.260 0.090 53.460 4.300 ;
        RECT 54.620 0.090 56.820 4.300 ;
        RECT 57.980 0.090 60.180 4.300 ;
        RECT 61.340 0.090 63.540 4.300 ;
        RECT 64.700 0.090 66.900 4.300 ;
        RECT 68.060 0.090 70.260 4.300 ;
        RECT 71.420 0.090 73.620 4.300 ;
        RECT 74.780 0.090 76.980 4.300 ;
        RECT 78.140 0.090 80.340 4.300 ;
        RECT 81.500 0.090 83.700 4.300 ;
        RECT 84.860 0.090 87.060 4.300 ;
        RECT 88.220 0.090 90.420 4.300 ;
        RECT 91.580 0.090 93.780 4.300 ;
        RECT 94.940 0.090 97.140 4.300 ;
        RECT 98.300 0.090 100.500 4.300 ;
        RECT 101.660 0.090 103.860 4.300 ;
        RECT 105.020 0.090 107.220 4.300 ;
        RECT 108.380 0.090 110.580 4.300 ;
        RECT 111.740 0.090 113.940 4.300 ;
        RECT 115.100 0.090 500.340 4.300 ;
        RECT 501.500 0.090 503.700 4.300 ;
        RECT 504.860 0.090 507.060 4.300 ;
        RECT 508.220 0.090 510.420 4.300 ;
        RECT 511.580 0.090 513.780 4.300 ;
        RECT 514.940 0.090 517.140 4.300 ;
        RECT 518.300 0.090 520.500 4.300 ;
        RECT 521.660 0.090 523.860 4.300 ;
        RECT 525.020 0.090 527.220 4.300 ;
        RECT 528.380 0.090 530.580 4.300 ;
        RECT 531.740 0.090 533.940 4.300 ;
        RECT 535.100 0.090 537.300 4.300 ;
        RECT 538.460 0.090 540.660 4.300 ;
        RECT 541.820 0.090 544.020 4.300 ;
        RECT 545.180 0.090 547.380 4.300 ;
        RECT 548.540 0.090 550.740 4.300 ;
        RECT 551.900 0.090 554.100 4.300 ;
        RECT 555.260 0.090 557.460 4.300 ;
        RECT 558.620 0.090 560.820 4.300 ;
        RECT 561.980 0.090 564.180 4.300 ;
        RECT 565.340 0.090 567.540 4.300 ;
        RECT 568.700 0.090 570.900 4.300 ;
        RECT 572.060 0.090 574.260 4.300 ;
        RECT 575.420 0.090 577.620 4.300 ;
        RECT 578.780 0.090 580.980 4.300 ;
        RECT 582.140 0.090 584.340 4.300 ;
        RECT 585.500 0.090 587.700 4.300 ;
        RECT 588.860 0.090 591.060 4.300 ;
        RECT 592.220 0.090 594.420 4.300 ;
        RECT 595.580 0.090 597.780 4.300 ;
        RECT 598.940 0.090 601.140 4.300 ;
        RECT 602.300 0.090 604.500 4.300 ;
        RECT 605.660 0.090 607.860 4.300 ;
        RECT 609.020 0.090 611.220 4.300 ;
        RECT 612.380 0.090 614.580 4.300 ;
        RECT 615.740 0.090 617.940 4.300 ;
        RECT 619.100 0.090 621.300 4.300 ;
        RECT 622.460 0.090 624.660 4.300 ;
        RECT 625.820 0.090 628.020 4.300 ;
        RECT 629.180 0.090 631.380 4.300 ;
        RECT 632.540 0.090 634.740 4.300 ;
        RECT 635.900 0.090 638.100 4.300 ;
        RECT 639.260 0.090 648.180 4.300 ;
        RECT 649.340 0.090 651.540 4.300 ;
        RECT 652.700 0.090 654.900 4.300 ;
        RECT 656.060 0.090 671.700 4.300 ;
        RECT 672.860 0.090 675.060 4.300 ;
        RECT 676.220 0.090 678.420 4.300 ;
        RECT 679.580 0.090 681.780 4.300 ;
        RECT 682.940 0.090 685.140 4.300 ;
        RECT 686.300 0.090 688.500 4.300 ;
        RECT 689.660 0.090 691.860 4.300 ;
        RECT 693.020 0.090 695.220 4.300 ;
        RECT 696.380 0.090 698.580 4.300 ;
        RECT 699.740 0.090 701.940 4.300 ;
        RECT 703.100 0.090 705.300 4.300 ;
        RECT 706.460 0.090 708.660 4.300 ;
        RECT 709.820 0.090 712.020 4.300 ;
        RECT 713.180 0.090 715.380 4.300 ;
        RECT 716.540 0.090 718.740 4.300 ;
        RECT 719.900 0.090 722.100 4.300 ;
        RECT 723.260 0.090 725.460 4.300 ;
        RECT 726.620 0.090 728.820 4.300 ;
        RECT 729.980 0.090 732.180 4.300 ;
        RECT 733.340 0.090 735.540 4.300 ;
        RECT 736.700 0.090 738.900 4.300 ;
        RECT 740.060 0.090 742.260 4.300 ;
        RECT 743.420 0.090 745.620 4.300 ;
        RECT 746.780 0.090 748.980 4.300 ;
        RECT 750.140 0.090 752.340 4.300 ;
      LAYER Metal3 ;
        RECT 4.000 555.260 753.110 756.700 ;
        RECT 4.000 554.100 751.400 555.260 ;
        RECT 4.000 551.900 753.110 554.100 ;
        RECT 4.000 550.740 751.400 551.900 ;
        RECT 4.000 548.540 753.110 550.740 ;
        RECT 4.000 547.380 751.400 548.540 ;
        RECT 4.000 545.180 753.110 547.380 ;
        RECT 4.000 544.020 751.400 545.180 ;
        RECT 4.000 541.820 753.110 544.020 ;
        RECT 4.000 540.660 751.400 541.820 ;
        RECT 4.000 538.460 753.110 540.660 ;
        RECT 4.000 537.300 751.400 538.460 ;
        RECT 4.000 535.100 753.110 537.300 ;
        RECT 4.000 533.940 751.400 535.100 ;
        RECT 4.000 531.740 753.110 533.940 ;
        RECT 4.000 530.580 751.400 531.740 ;
        RECT 4.000 528.380 753.110 530.580 ;
        RECT 4.000 527.220 751.400 528.380 ;
        RECT 4.000 525.020 753.110 527.220 ;
        RECT 4.000 523.860 751.400 525.020 ;
        RECT 4.000 521.660 753.110 523.860 ;
        RECT 4.000 520.500 751.400 521.660 ;
        RECT 4.000 518.300 753.110 520.500 ;
        RECT 4.000 517.140 751.400 518.300 ;
        RECT 4.000 514.940 753.110 517.140 ;
        RECT 4.000 513.780 751.400 514.940 ;
        RECT 4.000 511.580 753.110 513.780 ;
        RECT 4.000 510.420 751.400 511.580 ;
        RECT 4.000 508.220 753.110 510.420 ;
        RECT 4.000 507.060 751.400 508.220 ;
        RECT 4.000 504.860 753.110 507.060 ;
        RECT 4.000 503.700 751.400 504.860 ;
        RECT 4.000 501.500 753.110 503.700 ;
        RECT 4.000 500.340 751.400 501.500 ;
        RECT 4.000 498.140 753.110 500.340 ;
        RECT 4.000 496.980 751.400 498.140 ;
        RECT 4.000 494.780 753.110 496.980 ;
        RECT 4.000 493.620 751.400 494.780 ;
        RECT 4.000 491.420 753.110 493.620 ;
        RECT 4.000 490.260 751.400 491.420 ;
        RECT 4.000 488.060 753.110 490.260 ;
        RECT 4.000 486.900 751.400 488.060 ;
        RECT 4.000 484.700 753.110 486.900 ;
        RECT 4.000 483.540 751.400 484.700 ;
        RECT 4.000 481.340 753.110 483.540 ;
        RECT 4.000 480.180 751.400 481.340 ;
        RECT 4.000 477.980 753.110 480.180 ;
        RECT 4.000 476.820 751.400 477.980 ;
        RECT 4.000 474.620 753.110 476.820 ;
        RECT 4.000 473.460 751.400 474.620 ;
        RECT 4.000 471.260 753.110 473.460 ;
        RECT 4.000 470.100 751.400 471.260 ;
        RECT 4.000 467.900 753.110 470.100 ;
        RECT 4.000 466.740 751.400 467.900 ;
        RECT 4.000 464.540 753.110 466.740 ;
        RECT 4.000 463.380 751.400 464.540 ;
        RECT 4.000 461.180 753.110 463.380 ;
        RECT 4.000 460.020 751.400 461.180 ;
        RECT 4.000 457.820 753.110 460.020 ;
        RECT 4.000 456.660 751.400 457.820 ;
        RECT 4.000 454.460 753.110 456.660 ;
        RECT 4.000 453.300 751.400 454.460 ;
        RECT 4.000 451.100 753.110 453.300 ;
        RECT 4.000 449.940 751.400 451.100 ;
        RECT 4.000 447.740 753.110 449.940 ;
        RECT 4.000 446.580 751.400 447.740 ;
        RECT 4.000 444.380 753.110 446.580 ;
        RECT 4.000 443.220 751.400 444.380 ;
        RECT 4.000 441.020 753.110 443.220 ;
        RECT 4.000 439.860 751.400 441.020 ;
        RECT 4.000 437.660 753.110 439.860 ;
        RECT 4.000 436.500 751.400 437.660 ;
        RECT 4.000 434.300 753.110 436.500 ;
        RECT 4.000 433.140 751.400 434.300 ;
        RECT 4.000 430.940 753.110 433.140 ;
        RECT 4.000 429.780 751.400 430.940 ;
        RECT 4.000 427.580 753.110 429.780 ;
        RECT 4.000 426.420 751.400 427.580 ;
        RECT 4.000 424.220 753.110 426.420 ;
        RECT 4.000 423.060 751.400 424.220 ;
        RECT 4.000 420.860 753.110 423.060 ;
        RECT 4.000 419.700 751.400 420.860 ;
        RECT 4.000 417.500 753.110 419.700 ;
        RECT 4.000 416.340 751.400 417.500 ;
        RECT 4.000 414.140 753.110 416.340 ;
        RECT 4.000 412.980 751.400 414.140 ;
        RECT 4.000 410.780 753.110 412.980 ;
        RECT 4.000 409.620 751.400 410.780 ;
        RECT 4.000 407.420 753.110 409.620 ;
        RECT 4.000 406.260 751.400 407.420 ;
        RECT 4.000 404.060 753.110 406.260 ;
        RECT 4.000 402.900 751.400 404.060 ;
        RECT 4.000 400.700 753.110 402.900 ;
        RECT 4.000 399.540 751.400 400.700 ;
        RECT 4.000 397.340 753.110 399.540 ;
        RECT 4.000 396.180 751.400 397.340 ;
        RECT 4.000 393.980 753.110 396.180 ;
        RECT 4.000 392.820 751.400 393.980 ;
        RECT 4.000 390.620 753.110 392.820 ;
        RECT 4.000 389.460 751.400 390.620 ;
        RECT 4.000 387.260 753.110 389.460 ;
        RECT 4.000 386.100 751.400 387.260 ;
        RECT 4.000 383.900 753.110 386.100 ;
        RECT 4.000 382.740 751.400 383.900 ;
        RECT 4.000 380.540 753.110 382.740 ;
        RECT 4.000 379.380 751.400 380.540 ;
        RECT 4.000 377.180 753.110 379.380 ;
        RECT 4.000 376.020 751.400 377.180 ;
        RECT 4.000 373.820 753.110 376.020 ;
        RECT 4.000 372.660 751.400 373.820 ;
        RECT 4.000 370.460 753.110 372.660 ;
        RECT 4.000 369.300 751.400 370.460 ;
        RECT 4.000 367.100 753.110 369.300 ;
        RECT 4.000 365.940 751.400 367.100 ;
        RECT 4.000 363.740 753.110 365.940 ;
        RECT 4.000 362.580 751.400 363.740 ;
        RECT 4.000 360.380 753.110 362.580 ;
        RECT 4.000 359.220 751.400 360.380 ;
        RECT 4.000 357.020 753.110 359.220 ;
        RECT 4.000 355.860 751.400 357.020 ;
        RECT 4.000 353.660 753.110 355.860 ;
        RECT 4.000 352.500 751.400 353.660 ;
        RECT 4.000 350.300 753.110 352.500 ;
        RECT 4.000 349.140 751.400 350.300 ;
        RECT 4.000 346.940 753.110 349.140 ;
        RECT 4.000 345.780 751.400 346.940 ;
        RECT 4.000 343.580 753.110 345.780 ;
        RECT 4.000 342.420 751.400 343.580 ;
        RECT 4.000 340.220 753.110 342.420 ;
        RECT 4.000 339.060 751.400 340.220 ;
        RECT 4.000 336.860 753.110 339.060 ;
        RECT 4.000 335.700 751.400 336.860 ;
        RECT 4.000 333.500 753.110 335.700 ;
        RECT 4.000 332.340 751.400 333.500 ;
        RECT 4.000 330.140 753.110 332.340 ;
        RECT 4.000 328.980 751.400 330.140 ;
        RECT 4.000 326.780 753.110 328.980 ;
        RECT 4.000 325.620 751.400 326.780 ;
        RECT 4.000 323.420 753.110 325.620 ;
        RECT 4.000 322.260 751.400 323.420 ;
        RECT 4.000 320.060 753.110 322.260 ;
        RECT 4.000 318.900 751.400 320.060 ;
        RECT 4.000 316.700 753.110 318.900 ;
        RECT 4.000 315.540 751.400 316.700 ;
        RECT 4.000 313.340 753.110 315.540 ;
        RECT 4.000 312.180 751.400 313.340 ;
        RECT 4.000 309.980 753.110 312.180 ;
        RECT 4.000 308.820 751.400 309.980 ;
        RECT 4.000 306.620 753.110 308.820 ;
        RECT 4.300 305.460 751.400 306.620 ;
        RECT 4.000 303.260 753.110 305.460 ;
        RECT 4.000 302.100 751.400 303.260 ;
        RECT 4.000 299.900 753.110 302.100 ;
        RECT 4.000 298.740 751.400 299.900 ;
        RECT 4.000 296.540 753.110 298.740 ;
        RECT 4.000 295.380 751.400 296.540 ;
        RECT 4.000 293.180 753.110 295.380 ;
        RECT 4.000 292.020 751.400 293.180 ;
        RECT 4.000 289.820 753.110 292.020 ;
        RECT 4.000 288.660 751.400 289.820 ;
        RECT 4.000 286.460 753.110 288.660 ;
        RECT 4.000 285.300 751.400 286.460 ;
        RECT 4.000 283.100 753.110 285.300 ;
        RECT 4.000 281.940 751.400 283.100 ;
        RECT 4.000 279.740 753.110 281.940 ;
        RECT 4.000 278.580 751.400 279.740 ;
        RECT 4.000 276.380 753.110 278.580 ;
        RECT 4.000 275.220 751.400 276.380 ;
        RECT 4.000 273.020 753.110 275.220 ;
        RECT 4.000 271.860 751.400 273.020 ;
        RECT 4.000 269.660 753.110 271.860 ;
        RECT 4.000 268.500 751.400 269.660 ;
        RECT 4.000 266.300 753.110 268.500 ;
        RECT 4.000 265.140 751.400 266.300 ;
        RECT 4.000 262.940 753.110 265.140 ;
        RECT 4.000 261.780 751.400 262.940 ;
        RECT 4.000 259.580 753.110 261.780 ;
        RECT 4.000 258.420 751.400 259.580 ;
        RECT 4.000 256.220 753.110 258.420 ;
        RECT 4.000 255.060 751.400 256.220 ;
        RECT 4.000 252.860 753.110 255.060 ;
        RECT 4.000 251.700 751.400 252.860 ;
        RECT 4.000 249.500 753.110 251.700 ;
        RECT 4.000 248.340 751.400 249.500 ;
        RECT 4.000 246.140 753.110 248.340 ;
        RECT 4.000 244.980 751.400 246.140 ;
        RECT 4.000 242.780 753.110 244.980 ;
        RECT 4.000 241.620 751.400 242.780 ;
        RECT 4.000 239.420 753.110 241.620 ;
        RECT 4.000 238.260 751.400 239.420 ;
        RECT 4.000 236.060 753.110 238.260 ;
        RECT 4.000 234.900 751.400 236.060 ;
        RECT 4.000 232.700 753.110 234.900 ;
        RECT 4.000 231.540 751.400 232.700 ;
        RECT 4.000 229.340 753.110 231.540 ;
        RECT 4.000 228.180 751.400 229.340 ;
        RECT 4.000 225.980 753.110 228.180 ;
        RECT 4.000 224.820 751.400 225.980 ;
        RECT 4.000 222.620 753.110 224.820 ;
        RECT 4.000 221.460 751.400 222.620 ;
        RECT 4.000 219.260 753.110 221.460 ;
        RECT 4.000 218.100 751.400 219.260 ;
        RECT 4.000 215.900 753.110 218.100 ;
        RECT 4.000 214.740 751.400 215.900 ;
        RECT 4.000 212.540 753.110 214.740 ;
        RECT 4.000 211.380 751.400 212.540 ;
        RECT 4.000 209.180 753.110 211.380 ;
        RECT 4.000 208.020 751.400 209.180 ;
        RECT 4.000 205.820 753.110 208.020 ;
        RECT 4.000 204.660 751.400 205.820 ;
        RECT 4.000 202.460 753.110 204.660 ;
        RECT 4.000 201.300 751.400 202.460 ;
        RECT 4.000 199.100 753.110 201.300 ;
        RECT 4.000 197.940 751.400 199.100 ;
        RECT 4.000 195.740 753.110 197.940 ;
        RECT 4.000 194.580 751.400 195.740 ;
        RECT 4.000 192.380 753.110 194.580 ;
        RECT 4.000 191.220 751.400 192.380 ;
        RECT 4.000 189.020 753.110 191.220 ;
        RECT 4.000 187.860 751.400 189.020 ;
        RECT 4.000 185.660 753.110 187.860 ;
        RECT 4.000 184.500 751.400 185.660 ;
        RECT 4.000 182.300 753.110 184.500 ;
        RECT 4.000 181.140 751.400 182.300 ;
        RECT 4.000 178.940 753.110 181.140 ;
        RECT 4.000 177.780 751.400 178.940 ;
        RECT 4.000 175.580 753.110 177.780 ;
        RECT 4.000 174.420 751.400 175.580 ;
        RECT 4.000 172.220 753.110 174.420 ;
        RECT 4.000 171.060 751.400 172.220 ;
        RECT 4.000 168.860 753.110 171.060 ;
        RECT 4.000 167.700 751.400 168.860 ;
        RECT 4.000 165.500 753.110 167.700 ;
        RECT 4.000 164.340 751.400 165.500 ;
        RECT 4.000 162.140 753.110 164.340 ;
        RECT 4.000 160.980 751.400 162.140 ;
        RECT 4.000 158.780 753.110 160.980 ;
        RECT 4.000 157.620 751.400 158.780 ;
        RECT 4.000 155.420 753.110 157.620 ;
        RECT 4.000 154.260 751.400 155.420 ;
        RECT 4.000 152.060 753.110 154.260 ;
        RECT 4.000 150.900 751.400 152.060 ;
        RECT 4.000 148.700 753.110 150.900 ;
        RECT 4.000 147.540 751.400 148.700 ;
        RECT 4.000 145.340 753.110 147.540 ;
        RECT 4.000 144.180 751.400 145.340 ;
        RECT 4.000 141.980 753.110 144.180 ;
        RECT 4.000 140.820 751.400 141.980 ;
        RECT 4.000 138.620 753.110 140.820 ;
        RECT 4.000 137.460 751.400 138.620 ;
        RECT 4.000 135.260 753.110 137.460 ;
        RECT 4.000 134.100 751.400 135.260 ;
        RECT 4.000 131.900 753.110 134.100 ;
        RECT 4.000 130.740 751.400 131.900 ;
        RECT 4.000 128.540 753.110 130.740 ;
        RECT 4.000 127.380 751.400 128.540 ;
        RECT 4.000 125.180 753.110 127.380 ;
        RECT 4.000 124.020 751.400 125.180 ;
        RECT 4.000 121.820 753.110 124.020 ;
        RECT 4.000 120.660 751.400 121.820 ;
        RECT 4.000 118.460 753.110 120.660 ;
        RECT 4.000 117.300 751.400 118.460 ;
        RECT 4.000 115.100 753.110 117.300 ;
        RECT 4.000 113.940 751.400 115.100 ;
        RECT 4.000 111.740 753.110 113.940 ;
        RECT 4.000 110.580 751.400 111.740 ;
        RECT 4.000 108.380 753.110 110.580 ;
        RECT 4.000 107.220 751.400 108.380 ;
        RECT 4.000 105.020 753.110 107.220 ;
        RECT 4.000 103.860 751.400 105.020 ;
        RECT 4.000 101.660 753.110 103.860 ;
        RECT 4.000 100.500 751.400 101.660 ;
        RECT 4.000 98.300 753.110 100.500 ;
        RECT 4.000 97.140 751.400 98.300 ;
        RECT 4.000 94.940 753.110 97.140 ;
        RECT 4.000 93.780 751.400 94.940 ;
        RECT 4.000 91.580 753.110 93.780 ;
        RECT 4.000 90.420 751.400 91.580 ;
        RECT 4.000 88.220 753.110 90.420 ;
        RECT 4.000 87.060 751.400 88.220 ;
        RECT 4.000 84.860 753.110 87.060 ;
        RECT 4.000 83.700 751.400 84.860 ;
        RECT 4.000 81.500 753.110 83.700 ;
        RECT 4.000 80.340 751.400 81.500 ;
        RECT 4.000 78.140 753.110 80.340 ;
        RECT 4.000 76.980 751.400 78.140 ;
        RECT 4.000 74.780 753.110 76.980 ;
        RECT 4.000 73.620 751.400 74.780 ;
        RECT 4.000 71.420 753.110 73.620 ;
        RECT 4.000 70.260 751.400 71.420 ;
        RECT 4.000 68.060 753.110 70.260 ;
        RECT 4.000 66.900 751.400 68.060 ;
        RECT 4.000 64.700 753.110 66.900 ;
        RECT 4.000 63.540 751.400 64.700 ;
        RECT 4.000 61.340 753.110 63.540 ;
        RECT 4.000 60.180 751.400 61.340 ;
        RECT 4.000 57.980 753.110 60.180 ;
        RECT 4.000 56.820 751.400 57.980 ;
        RECT 4.000 54.620 753.110 56.820 ;
        RECT 4.000 53.460 751.400 54.620 ;
        RECT 4.000 51.260 753.110 53.460 ;
        RECT 4.000 50.100 751.400 51.260 ;
        RECT 4.000 47.900 753.110 50.100 ;
        RECT 4.000 46.740 751.400 47.900 ;
        RECT 4.000 44.540 753.110 46.740 ;
        RECT 4.000 43.380 751.400 44.540 ;
        RECT 4.000 41.180 753.110 43.380 ;
        RECT 4.000 40.020 751.400 41.180 ;
        RECT 4.000 37.820 753.110 40.020 ;
        RECT 4.000 36.660 751.400 37.820 ;
        RECT 4.000 34.460 753.110 36.660 ;
        RECT 4.000 33.300 751.400 34.460 ;
        RECT 4.000 31.100 753.110 33.300 ;
        RECT 4.000 29.940 751.400 31.100 ;
        RECT 4.000 27.740 753.110 29.940 ;
        RECT 4.000 26.580 751.400 27.740 ;
        RECT 4.000 24.380 753.110 26.580 ;
        RECT 4.000 23.220 751.400 24.380 ;
        RECT 4.000 21.020 753.110 23.220 ;
        RECT 4.000 19.860 751.400 21.020 ;
        RECT 4.000 17.660 753.110 19.860 ;
        RECT 4.000 16.500 751.400 17.660 ;
        RECT 4.000 14.300 753.110 16.500 ;
        RECT 4.000 13.140 751.400 14.300 ;
        RECT 4.000 10.940 753.110 13.140 ;
        RECT 4.000 9.780 751.400 10.940 ;
        RECT 4.000 7.580 753.110 9.780 ;
        RECT 4.000 6.420 751.400 7.580 ;
        RECT 4.000 4.220 753.110 6.420 ;
        RECT 4.000 3.060 751.400 4.220 ;
        RECT 4.000 0.860 753.110 3.060 ;
        RECT 4.000 0.140 751.400 0.860 ;
      LAYER Metal4 ;
        RECT 58.380 16.890 98.740 734.630 ;
        RECT 100.940 16.890 175.540 734.630 ;
        RECT 177.740 16.890 252.340 734.630 ;
        RECT 254.540 16.890 329.140 734.630 ;
        RECT 331.340 16.890 405.940 734.630 ;
        RECT 408.140 16.890 482.740 734.630 ;
        RECT 484.940 16.890 559.540 734.630 ;
        RECT 561.740 16.890 636.340 734.630 ;
        RECT 638.540 16.890 713.140 734.630 ;
        RECT 715.340 16.890 745.220 734.630 ;
      LAYER Metal5 ;
        RECT 84.060 108.230 745.300 555.070 ;
  END
END serv_rf_top
END LIBRARY

