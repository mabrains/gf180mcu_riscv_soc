VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO analog_wrapper
  CLASS BLOCK ;
  FOREIGN analog_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2550.000 BY 1370.000 ;
  OBS
      LAYER Metal1 ;
        RECT 0.000 0.000 2550.000 1370.000 ;
      LAYER Metal2 ;
        RECT 0.000 0.000 2550.000 1370.000 ;          
      LAYER Metal3 ;
        RECT 0.000 0.000 2550.000 1370.000 ;  
      LAYER Metal4 ;
        RECT 0.000 0.000 2550.000 1370.000 ;
      LAYER Metal5 ;
        RECT 0.000 0.000 2550.000 1370.000 ;
      LAYER via1 ;
        RECT 0.000 0.000 2550.000 1370.000 ;
      LAYER via2 ;
        RECT 0.000 0.000 2550.000 1370.000 ;          
      LAYER via3 ;
        RECT 0.000 0.000 2550.000 1370.000 ;  
      LAYER via4 ;
        RECT 0.000 0.000 2550.000 1370.000 ;
      LAYER contact ;
        RECT 0.000 0.000 2550.000 1370.000 ;                   
  END
END analog_wrapper
END LIBRARY
