magic
tech gf180mcuD
magscale 1 5
timestamp 1700584330
<< obsm1 >>
rect 672 1359 9735 6369
<< metal2 >>
rect 1232 7600 1288 8000
rect 3696 7600 3752 8000
rect 6160 7600 6216 8000
rect 8624 7600 8680 8000
rect 672 0 728 400
rect 896 0 952 400
rect 1120 0 1176 400
rect 1344 0 1400 400
rect 1568 0 1624 400
rect 1792 0 1848 400
rect 2016 0 2072 400
rect 2240 0 2296 400
rect 2464 0 2520 400
rect 2688 0 2744 400
rect 2912 0 2968 400
rect 3136 0 3192 400
rect 3360 0 3416 400
rect 3584 0 3640 400
rect 3808 0 3864 400
rect 4032 0 4088 400
rect 4256 0 4312 400
rect 4480 0 4536 400
rect 4704 0 4760 400
rect 4928 0 4984 400
rect 5152 0 5208 400
rect 5376 0 5432 400
rect 5600 0 5656 400
rect 5824 0 5880 400
rect 6048 0 6104 400
rect 6272 0 6328 400
rect 6496 0 6552 400
rect 6720 0 6776 400
rect 6944 0 7000 400
rect 7168 0 7224 400
rect 7392 0 7448 400
rect 7616 0 7672 400
rect 7840 0 7896 400
rect 8064 0 8120 400
rect 8288 0 8344 400
rect 8512 0 8568 400
rect 8736 0 8792 400
rect 8960 0 9016 400
rect 9184 0 9240 400
<< obsm2 >>
rect 630 7570 1202 7663
rect 1318 7570 3666 7663
rect 3782 7570 6130 7663
rect 6246 7570 8594 7663
rect 8710 7570 9730 7663
rect 630 430 9730 7570
rect 630 400 642 430
rect 758 400 866 430
rect 982 400 1090 430
rect 1206 400 1314 430
rect 1430 400 1538 430
rect 1654 400 1762 430
rect 1878 400 1986 430
rect 2102 400 2210 430
rect 2326 400 2434 430
rect 2550 400 2658 430
rect 2774 400 2882 430
rect 2998 400 3106 430
rect 3222 400 3330 430
rect 3446 400 3554 430
rect 3670 400 3778 430
rect 3894 400 4002 430
rect 4118 400 4226 430
rect 4342 400 4450 430
rect 4566 400 4674 430
rect 4790 400 4898 430
rect 5014 400 5122 430
rect 5238 400 5346 430
rect 5462 400 5570 430
rect 5686 400 5794 430
rect 5910 400 6018 430
rect 6134 400 6242 430
rect 6358 400 6466 430
rect 6582 400 6690 430
rect 6806 400 6914 430
rect 7030 400 7138 430
rect 7254 400 7362 430
rect 7478 400 7586 430
rect 7702 400 7810 430
rect 7926 400 8034 430
rect 8150 400 8258 430
rect 8374 400 8482 430
rect 8598 400 8706 430
rect 8822 400 8930 430
rect 9046 400 9154 430
rect 9270 400 9730 430
<< metal3 >>
rect 0 7616 400 7672
rect 0 7392 400 7448
rect 0 7168 400 7224
rect 0 6944 400 7000
rect 0 6720 400 6776
rect 0 6496 400 6552
rect 0 6272 400 6328
rect 0 6048 400 6104
rect 9600 5936 10000 5992
rect 0 5824 400 5880
rect 0 5600 400 5656
rect 0 5376 400 5432
rect 0 5152 400 5208
rect 0 4928 400 4984
rect 0 4704 400 4760
rect 0 4480 400 4536
rect 0 4256 400 4312
rect 0 4032 400 4088
rect 0 3808 400 3864
rect 0 3584 400 3640
rect 0 3360 400 3416
rect 0 3136 400 3192
rect 0 2912 400 2968
rect 0 2688 400 2744
rect 0 2464 400 2520
rect 0 2240 400 2296
rect 0 2016 400 2072
rect 9600 1904 10000 1960
rect 0 1792 400 1848
rect 0 1568 400 1624
rect 0 1344 400 1400
rect 0 1120 400 1176
rect 0 896 400 952
rect 0 672 400 728
rect 0 448 400 504
rect 0 224 400 280
<< obsm3 >>
rect 430 7586 9735 7658
rect 400 7478 9735 7586
rect 430 7362 9735 7478
rect 400 7254 9735 7362
rect 430 7138 9735 7254
rect 400 7030 9735 7138
rect 430 6914 9735 7030
rect 400 6806 9735 6914
rect 430 6690 9735 6806
rect 400 6582 9735 6690
rect 430 6466 9735 6582
rect 400 6358 9735 6466
rect 430 6242 9735 6358
rect 400 6134 9735 6242
rect 430 6022 9735 6134
rect 430 6018 9570 6022
rect 400 5910 9570 6018
rect 430 5906 9570 5910
rect 430 5794 9735 5906
rect 400 5686 9735 5794
rect 430 5570 9735 5686
rect 400 5462 9735 5570
rect 430 5346 9735 5462
rect 400 5238 9735 5346
rect 430 5122 9735 5238
rect 400 5014 9735 5122
rect 430 4898 9735 5014
rect 400 4790 9735 4898
rect 430 4674 9735 4790
rect 400 4566 9735 4674
rect 430 4450 9735 4566
rect 400 4342 9735 4450
rect 430 4226 9735 4342
rect 400 4118 9735 4226
rect 430 4002 9735 4118
rect 400 3894 9735 4002
rect 430 3778 9735 3894
rect 400 3670 9735 3778
rect 430 3554 9735 3670
rect 400 3446 9735 3554
rect 430 3330 9735 3446
rect 400 3222 9735 3330
rect 430 3106 9735 3222
rect 400 2998 9735 3106
rect 430 2882 9735 2998
rect 400 2774 9735 2882
rect 430 2658 9735 2774
rect 400 2550 9735 2658
rect 430 2434 9735 2550
rect 400 2326 9735 2434
rect 430 2210 9735 2326
rect 400 2102 9735 2210
rect 430 1990 9735 2102
rect 430 1986 9570 1990
rect 400 1878 9570 1986
rect 430 1874 9570 1878
rect 430 1762 9735 1874
rect 400 1654 9735 1762
rect 430 1538 9735 1654
rect 400 1430 9735 1538
rect 430 1314 9735 1430
rect 400 1206 9735 1314
rect 430 1090 9735 1206
rect 400 982 9735 1090
rect 430 866 9735 982
rect 400 758 9735 866
rect 430 642 9735 758
rect 400 534 9735 642
rect 430 418 9735 534
rect 400 310 9735 418
rect 430 238 9735 310
<< metal4 >>
rect 1670 1538 1830 6302
rect 2748 1538 2908 6302
rect 3826 1538 3986 6302
rect 4904 1538 5064 6302
rect 5982 1538 6142 6302
rect 7060 1538 7220 6302
rect 8138 1538 8298 6302
rect 9216 1538 9376 6302
<< obsm4 >>
rect 910 1508 1640 5647
rect 1860 1508 2718 5647
rect 2938 1508 3796 5647
rect 4016 1508 4874 5647
rect 5094 1508 5952 5647
rect 6172 1508 7030 5647
rect 7250 1508 8108 5647
rect 8328 1508 8834 5647
rect 910 457 8834 1508
<< labels >>
rlabel metal4 s 1670 1538 1830 6302 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 3826 1538 3986 6302 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 5982 1538 6142 6302 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 8138 1538 8298 6302 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 2748 1538 2908 6302 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 4904 1538 5064 6302 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 7060 1538 7220 6302 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 9216 1538 9376 6302 6 VSS
port 2 nsew ground bidirectional
rlabel metal3 s 9600 1904 10000 1960 6 buttons[0]
port 3 nsew signal input
rlabel metal3 s 9600 5936 10000 5992 6 buttons[1]
port 4 nsew signal input
rlabel metal2 s 8960 0 9016 400 6 clk
port 5 nsew signal input
rlabel metal2 s 1344 0 1400 400 6 i_wb_addr[0]
port 6 nsew signal input
rlabel metal2 s 4032 0 4088 400 6 i_wb_addr[10]
port 7 nsew signal input
rlabel metal2 s 4256 0 4312 400 6 i_wb_addr[11]
port 8 nsew signal input
rlabel metal2 s 4480 0 4536 400 6 i_wb_addr[12]
port 9 nsew signal input
rlabel metal2 s 4704 0 4760 400 6 i_wb_addr[13]
port 10 nsew signal input
rlabel metal2 s 4928 0 4984 400 6 i_wb_addr[14]
port 11 nsew signal input
rlabel metal2 s 5152 0 5208 400 6 i_wb_addr[15]
port 12 nsew signal input
rlabel metal2 s 5376 0 5432 400 6 i_wb_addr[16]
port 13 nsew signal input
rlabel metal2 s 5600 0 5656 400 6 i_wb_addr[17]
port 14 nsew signal input
rlabel metal2 s 5824 0 5880 400 6 i_wb_addr[18]
port 15 nsew signal input
rlabel metal2 s 6048 0 6104 400 6 i_wb_addr[19]
port 16 nsew signal input
rlabel metal2 s 1792 0 1848 400 6 i_wb_addr[1]
port 17 nsew signal input
rlabel metal2 s 6272 0 6328 400 6 i_wb_addr[20]
port 18 nsew signal input
rlabel metal2 s 6496 0 6552 400 6 i_wb_addr[21]
port 19 nsew signal input
rlabel metal2 s 6720 0 6776 400 6 i_wb_addr[22]
port 20 nsew signal input
rlabel metal2 s 6944 0 7000 400 6 i_wb_addr[23]
port 21 nsew signal input
rlabel metal2 s 7168 0 7224 400 6 i_wb_addr[24]
port 22 nsew signal input
rlabel metal2 s 7392 0 7448 400 6 i_wb_addr[25]
port 23 nsew signal input
rlabel metal2 s 7616 0 7672 400 6 i_wb_addr[26]
port 24 nsew signal input
rlabel metal2 s 7840 0 7896 400 6 i_wb_addr[27]
port 25 nsew signal input
rlabel metal2 s 8064 0 8120 400 6 i_wb_addr[28]
port 26 nsew signal input
rlabel metal2 s 8288 0 8344 400 6 i_wb_addr[29]
port 27 nsew signal input
rlabel metal2 s 2240 0 2296 400 6 i_wb_addr[2]
port 28 nsew signal input
rlabel metal2 s 8512 0 8568 400 6 i_wb_addr[30]
port 29 nsew signal input
rlabel metal2 s 8736 0 8792 400 6 i_wb_addr[31]
port 30 nsew signal input
rlabel metal2 s 2464 0 2520 400 6 i_wb_addr[3]
port 31 nsew signal input
rlabel metal2 s 2688 0 2744 400 6 i_wb_addr[4]
port 32 nsew signal input
rlabel metal2 s 2912 0 2968 400 6 i_wb_addr[5]
port 33 nsew signal input
rlabel metal2 s 3136 0 3192 400 6 i_wb_addr[6]
port 34 nsew signal input
rlabel metal2 s 3360 0 3416 400 6 i_wb_addr[7]
port 35 nsew signal input
rlabel metal2 s 3584 0 3640 400 6 i_wb_addr[8]
port 36 nsew signal input
rlabel metal2 s 3808 0 3864 400 6 i_wb_addr[9]
port 37 nsew signal input
rlabel metal2 s 672 0 728 400 6 i_wb_cyc
port 38 nsew signal input
rlabel metal2 s 1568 0 1624 400 6 i_wb_data[0]
port 39 nsew signal input
rlabel metal2 s 2016 0 2072 400 6 i_wb_data[1]
port 40 nsew signal input
rlabel metal2 s 896 0 952 400 6 i_wb_stb
port 41 nsew signal input
rlabel metal2 s 1120 0 1176 400 6 i_wb_we
port 42 nsew signal input
rlabel metal2 s 8624 7600 8680 8000 6 led_enb[0]
port 43 nsew signal output
rlabel metal2 s 3696 7600 3752 8000 6 led_enb[1]
port 44 nsew signal output
rlabel metal2 s 6160 7600 6216 8000 6 leds[0]
port 45 nsew signal output
rlabel metal2 s 1232 7600 1288 8000 6 leds[1]
port 46 nsew signal output
rlabel metal3 s 0 224 400 280 6 o_wb_ack
port 47 nsew signal output
rlabel metal3 s 0 672 400 728 6 o_wb_data[0]
port 48 nsew signal output
rlabel metal3 s 0 2912 400 2968 6 o_wb_data[10]
port 49 nsew signal output
rlabel metal3 s 0 3136 400 3192 6 o_wb_data[11]
port 50 nsew signal output
rlabel metal3 s 0 3360 400 3416 6 o_wb_data[12]
port 51 nsew signal output
rlabel metal3 s 0 3584 400 3640 6 o_wb_data[13]
port 52 nsew signal output
rlabel metal3 s 0 3808 400 3864 6 o_wb_data[14]
port 53 nsew signal output
rlabel metal3 s 0 4032 400 4088 6 o_wb_data[15]
port 54 nsew signal output
rlabel metal3 s 0 4256 400 4312 6 o_wb_data[16]
port 55 nsew signal output
rlabel metal3 s 0 4480 400 4536 6 o_wb_data[17]
port 56 nsew signal output
rlabel metal3 s 0 4704 400 4760 6 o_wb_data[18]
port 57 nsew signal output
rlabel metal3 s 0 4928 400 4984 6 o_wb_data[19]
port 58 nsew signal output
rlabel metal3 s 0 896 400 952 6 o_wb_data[1]
port 59 nsew signal output
rlabel metal3 s 0 5152 400 5208 6 o_wb_data[20]
port 60 nsew signal output
rlabel metal3 s 0 5376 400 5432 6 o_wb_data[21]
port 61 nsew signal output
rlabel metal3 s 0 5600 400 5656 6 o_wb_data[22]
port 62 nsew signal output
rlabel metal3 s 0 5824 400 5880 6 o_wb_data[23]
port 63 nsew signal output
rlabel metal3 s 0 6048 400 6104 6 o_wb_data[24]
port 64 nsew signal output
rlabel metal3 s 0 6272 400 6328 6 o_wb_data[25]
port 65 nsew signal output
rlabel metal3 s 0 6496 400 6552 6 o_wb_data[26]
port 66 nsew signal output
rlabel metal3 s 0 6720 400 6776 6 o_wb_data[27]
port 67 nsew signal output
rlabel metal3 s 0 6944 400 7000 6 o_wb_data[28]
port 68 nsew signal output
rlabel metal3 s 0 7168 400 7224 6 o_wb_data[29]
port 69 nsew signal output
rlabel metal3 s 0 1120 400 1176 6 o_wb_data[2]
port 70 nsew signal output
rlabel metal3 s 0 7392 400 7448 6 o_wb_data[30]
port 71 nsew signal output
rlabel metal3 s 0 7616 400 7672 6 o_wb_data[31]
port 72 nsew signal output
rlabel metal3 s 0 1344 400 1400 6 o_wb_data[3]
port 73 nsew signal output
rlabel metal3 s 0 1568 400 1624 6 o_wb_data[4]
port 74 nsew signal output
rlabel metal3 s 0 1792 400 1848 6 o_wb_data[5]
port 75 nsew signal output
rlabel metal3 s 0 2016 400 2072 6 o_wb_data[6]
port 76 nsew signal output
rlabel metal3 s 0 2240 400 2296 6 o_wb_data[7]
port 77 nsew signal output
rlabel metal3 s 0 2464 400 2520 6 o_wb_data[8]
port 78 nsew signal output
rlabel metal3 s 0 2688 400 2744 6 o_wb_data[9]
port 79 nsew signal output
rlabel metal3 s 0 448 400 504 6 o_wb_stall
port 80 nsew signal output
rlabel metal2 s 9184 0 9240 400 6 reset
port 81 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 10000 8000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 383116
string GDS_FILE /home/farag/carvel_riscv_soc/gf180mcu_riscv_soc/openlane/wb_buttons_leds/runs/23_11_21_18_29/results/signoff/wb_buttons_leds.magic.gds
string GDS_START 127934
<< end >>

