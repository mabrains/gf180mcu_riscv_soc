magic
tech gf180mcuD
magscale 1 10
timestamp 1700747287
<< metal1 >>
rect 1344 16490 22624 16524
rect 1344 16438 3874 16490
rect 3926 16438 3978 16490
rect 4030 16438 4082 16490
rect 4134 16438 9194 16490
rect 9246 16438 9298 16490
rect 9350 16438 9402 16490
rect 9454 16438 14514 16490
rect 14566 16438 14618 16490
rect 14670 16438 14722 16490
rect 14774 16438 19834 16490
rect 19886 16438 19938 16490
rect 19990 16438 20042 16490
rect 20094 16438 22624 16490
rect 1344 16404 22624 16438
rect 1822 16322 1874 16334
rect 1822 16258 1874 16270
rect 21758 16322 21810 16334
rect 21758 16258 21810 16270
rect 7746 16158 7758 16210
rect 7810 16158 7822 16210
rect 17042 16158 17054 16210
rect 17106 16158 17118 16210
rect 8754 16046 8766 16098
rect 8818 16046 8830 16098
rect 3838 15986 3890 15998
rect 3838 15922 3890 15934
rect 4734 15986 4786 15998
rect 4734 15922 4786 15934
rect 10558 15986 10610 15998
rect 10558 15922 10610 15934
rect 13470 15986 13522 15998
rect 13470 15922 13522 15934
rect 19294 15986 19346 15998
rect 19294 15922 19346 15934
rect 2606 15874 2658 15886
rect 2606 15810 2658 15822
rect 3390 15874 3442 15886
rect 3390 15810 3442 15822
rect 9438 15874 9490 15886
rect 9438 15810 9490 15822
rect 17726 15874 17778 15886
rect 17726 15810 17778 15822
rect 20302 15874 20354 15886
rect 20302 15810 20354 15822
rect 20974 15874 21026 15886
rect 20974 15810 21026 15822
rect 1344 15706 22784 15740
rect 1344 15654 6534 15706
rect 6586 15654 6638 15706
rect 6690 15654 6742 15706
rect 6794 15654 11854 15706
rect 11906 15654 11958 15706
rect 12010 15654 12062 15706
rect 12114 15654 17174 15706
rect 17226 15654 17278 15706
rect 17330 15654 17382 15706
rect 17434 15654 22494 15706
rect 22546 15654 22598 15706
rect 22650 15654 22702 15706
rect 22754 15654 22784 15706
rect 1344 15620 22784 15654
rect 2606 15538 2658 15550
rect 2606 15474 2658 15486
rect 3054 15538 3106 15550
rect 3054 15474 3106 15486
rect 3502 15538 3554 15550
rect 3502 15474 3554 15486
rect 1710 15426 1762 15438
rect 1710 15362 1762 15374
rect 2158 15426 2210 15438
rect 2158 15362 2210 15374
rect 22206 15090 22258 15102
rect 22206 15026 22258 15038
rect 1344 14922 22624 14956
rect 1344 14870 3874 14922
rect 3926 14870 3978 14922
rect 4030 14870 4082 14922
rect 4134 14870 9194 14922
rect 9246 14870 9298 14922
rect 9350 14870 9402 14922
rect 9454 14870 14514 14922
rect 14566 14870 14618 14922
rect 14670 14870 14722 14922
rect 14774 14870 19834 14922
rect 19886 14870 19938 14922
rect 19990 14870 20042 14922
rect 20094 14870 22624 14922
rect 1344 14836 22624 14870
rect 1710 14306 1762 14318
rect 1710 14242 1762 14254
rect 2158 14306 2210 14318
rect 2158 14242 2210 14254
rect 1344 14138 22784 14172
rect 1344 14086 6534 14138
rect 6586 14086 6638 14138
rect 6690 14086 6742 14138
rect 6794 14086 11854 14138
rect 11906 14086 11958 14138
rect 12010 14086 12062 14138
rect 12114 14086 17174 14138
rect 17226 14086 17278 14138
rect 17330 14086 17382 14138
rect 17434 14086 22494 14138
rect 22546 14086 22598 14138
rect 22650 14086 22702 14138
rect 22754 14086 22784 14138
rect 1344 14052 22784 14086
rect 1710 13858 1762 13870
rect 1710 13794 1762 13806
rect 1344 13354 22624 13388
rect 1344 13302 3874 13354
rect 3926 13302 3978 13354
rect 4030 13302 4082 13354
rect 4134 13302 9194 13354
rect 9246 13302 9298 13354
rect 9350 13302 9402 13354
rect 9454 13302 14514 13354
rect 14566 13302 14618 13354
rect 14670 13302 14722 13354
rect 14774 13302 19834 13354
rect 19886 13302 19938 13354
rect 19990 13302 20042 13354
rect 20094 13302 22624 13354
rect 1344 13268 22624 13302
rect 1710 12850 1762 12862
rect 1710 12786 1762 12798
rect 22206 12850 22258 12862
rect 22206 12786 22258 12798
rect 2158 12738 2210 12750
rect 2158 12674 2210 12686
rect 21646 12738 21698 12750
rect 21646 12674 21698 12686
rect 21870 12738 21922 12750
rect 21870 12674 21922 12686
rect 1344 12570 22784 12604
rect 1344 12518 6534 12570
rect 6586 12518 6638 12570
rect 6690 12518 6742 12570
rect 6794 12518 11854 12570
rect 11906 12518 11958 12570
rect 12010 12518 12062 12570
rect 12114 12518 17174 12570
rect 17226 12518 17278 12570
rect 17330 12518 17382 12570
rect 17434 12518 22494 12570
rect 22546 12518 22598 12570
rect 22650 12518 22702 12570
rect 22754 12518 22784 12570
rect 1344 12484 22784 12518
rect 1710 12290 1762 12302
rect 1710 12226 1762 12238
rect 2158 12290 2210 12302
rect 2158 12226 2210 12238
rect 3838 12178 3890 12190
rect 3838 12114 3890 12126
rect 2830 12066 2882 12078
rect 2830 12002 2882 12014
rect 3278 12066 3330 12078
rect 3278 12002 3330 12014
rect 4286 12066 4338 12078
rect 4286 12002 4338 12014
rect 1344 11786 22624 11820
rect 1344 11734 3874 11786
rect 3926 11734 3978 11786
rect 4030 11734 4082 11786
rect 4134 11734 9194 11786
rect 9246 11734 9298 11786
rect 9350 11734 9402 11786
rect 9454 11734 14514 11786
rect 14566 11734 14618 11786
rect 14670 11734 14722 11786
rect 14774 11734 19834 11786
rect 19886 11734 19938 11786
rect 19990 11734 20042 11786
rect 20094 11734 22624 11786
rect 1344 11700 22624 11734
rect 4958 11506 5010 11518
rect 4958 11442 5010 11454
rect 1710 11170 1762 11182
rect 1710 11106 1762 11118
rect 2158 11170 2210 11182
rect 2158 11106 2210 11118
rect 2830 11170 2882 11182
rect 2830 11106 2882 11118
rect 3390 11170 3442 11182
rect 3390 11106 3442 11118
rect 3726 11170 3778 11182
rect 3726 11106 3778 11118
rect 4510 11170 4562 11182
rect 4510 11106 4562 11118
rect 9998 11170 10050 11182
rect 9998 11106 10050 11118
rect 1344 11002 22784 11036
rect 1344 10950 6534 11002
rect 6586 10950 6638 11002
rect 6690 10950 6742 11002
rect 6794 10950 11854 11002
rect 11906 10950 11958 11002
rect 12010 10950 12062 11002
rect 12114 10950 17174 11002
rect 17226 10950 17278 11002
rect 17330 10950 17382 11002
rect 17434 10950 22494 11002
rect 22546 10950 22598 11002
rect 22650 10950 22702 11002
rect 22754 10950 22784 11002
rect 1344 10916 22784 10950
rect 1710 10722 1762 10734
rect 1710 10658 1762 10670
rect 2158 10722 2210 10734
rect 2158 10658 2210 10670
rect 2606 10722 2658 10734
rect 2606 10658 2658 10670
rect 3054 10722 3106 10734
rect 3054 10658 3106 10670
rect 10222 10722 10274 10734
rect 10222 10658 10274 10670
rect 11118 10610 11170 10622
rect 9986 10558 9998 10610
rect 10050 10558 10062 10610
rect 11118 10546 11170 10558
rect 4062 10498 4114 10510
rect 4062 10434 4114 10446
rect 4622 10498 4674 10510
rect 4622 10434 4674 10446
rect 5182 10498 5234 10510
rect 5182 10434 5234 10446
rect 5630 10498 5682 10510
rect 5630 10434 5682 10446
rect 5966 10498 6018 10510
rect 5966 10434 6018 10446
rect 6526 10498 6578 10510
rect 6526 10434 6578 10446
rect 6974 10498 7026 10510
rect 6974 10434 7026 10446
rect 8990 10498 9042 10510
rect 8990 10434 9042 10446
rect 10670 10498 10722 10510
rect 10670 10434 10722 10446
rect 11678 10498 11730 10510
rect 11678 10434 11730 10446
rect 12126 10498 12178 10510
rect 12126 10434 12178 10446
rect 5954 10334 5966 10386
rect 6018 10383 6030 10386
rect 7074 10383 7086 10386
rect 6018 10337 7086 10383
rect 6018 10334 6030 10337
rect 7074 10334 7086 10337
rect 7138 10334 7150 10386
rect 10434 10334 10446 10386
rect 10498 10383 10510 10386
rect 10994 10383 11006 10386
rect 10498 10337 11006 10383
rect 10498 10334 10510 10337
rect 10994 10334 11006 10337
rect 11058 10334 11070 10386
rect 1344 10218 22624 10252
rect 1344 10166 3874 10218
rect 3926 10166 3978 10218
rect 4030 10166 4082 10218
rect 4134 10166 9194 10218
rect 9246 10166 9298 10218
rect 9350 10166 9402 10218
rect 9454 10166 14514 10218
rect 14566 10166 14618 10218
rect 14670 10166 14722 10218
rect 14774 10166 19834 10218
rect 19886 10166 19938 10218
rect 19990 10166 20042 10218
rect 20094 10166 22624 10218
rect 1344 10132 22624 10166
rect 12238 9826 12290 9838
rect 9762 9774 9774 9826
rect 9826 9774 9838 9826
rect 10770 9774 10782 9826
rect 10834 9774 10846 9826
rect 11442 9774 11454 9826
rect 11506 9774 11518 9826
rect 12238 9762 12290 9774
rect 4958 9714 5010 9726
rect 4958 9650 5010 9662
rect 8654 9714 8706 9726
rect 8654 9650 8706 9662
rect 1710 9602 1762 9614
rect 1710 9538 1762 9550
rect 2158 9602 2210 9614
rect 2158 9538 2210 9550
rect 2606 9602 2658 9614
rect 2606 9538 2658 9550
rect 3054 9602 3106 9614
rect 3054 9538 3106 9550
rect 3726 9602 3778 9614
rect 3726 9538 3778 9550
rect 4174 9602 4226 9614
rect 4174 9538 4226 9550
rect 4622 9602 4674 9614
rect 4622 9538 4674 9550
rect 4846 9602 4898 9614
rect 4846 9538 4898 9550
rect 5854 9602 5906 9614
rect 5854 9538 5906 9550
rect 6302 9602 6354 9614
rect 6302 9538 6354 9550
rect 6974 9602 7026 9614
rect 6974 9538 7026 9550
rect 7422 9602 7474 9614
rect 7422 9538 7474 9550
rect 7870 9602 7922 9614
rect 7870 9538 7922 9550
rect 8430 9602 8482 9614
rect 8430 9538 8482 9550
rect 8990 9602 9042 9614
rect 8990 9538 9042 9550
rect 9998 9602 10050 9614
rect 9998 9538 10050 9550
rect 10558 9602 10610 9614
rect 10558 9538 10610 9550
rect 11230 9602 11282 9614
rect 11230 9538 11282 9550
rect 11902 9602 11954 9614
rect 11902 9538 11954 9550
rect 12686 9602 12738 9614
rect 12686 9538 12738 9550
rect 20862 9602 20914 9614
rect 20862 9538 20914 9550
rect 22206 9602 22258 9614
rect 22206 9538 22258 9550
rect 1344 9434 22784 9468
rect 1344 9382 6534 9434
rect 6586 9382 6638 9434
rect 6690 9382 6742 9434
rect 6794 9382 11854 9434
rect 11906 9382 11958 9434
rect 12010 9382 12062 9434
rect 12114 9382 17174 9434
rect 17226 9382 17278 9434
rect 17330 9382 17382 9434
rect 17434 9382 22494 9434
rect 22546 9382 22598 9434
rect 22650 9382 22702 9434
rect 22754 9382 22784 9434
rect 1344 9348 22784 9382
rect 15150 9266 15202 9278
rect 15150 9202 15202 9214
rect 1822 9154 1874 9166
rect 1822 9090 1874 9102
rect 2270 9154 2322 9166
rect 2270 9090 2322 9102
rect 2718 9154 2770 9166
rect 2718 9090 2770 9102
rect 3278 9154 3330 9166
rect 3278 9090 3330 9102
rect 3390 9154 3442 9166
rect 3390 9090 3442 9102
rect 7086 9154 7138 9166
rect 7086 9090 7138 9102
rect 8094 9154 8146 9166
rect 8094 9090 8146 9102
rect 10110 9154 10162 9166
rect 10110 9090 10162 9102
rect 12126 9154 12178 9166
rect 12126 9090 12178 9102
rect 6862 9042 6914 9054
rect 6514 8990 6526 9042
rect 6578 8990 6590 9042
rect 6862 8978 6914 8990
rect 7198 9042 7250 9054
rect 7198 8978 7250 8990
rect 7758 9042 7810 9054
rect 7758 8978 7810 8990
rect 8430 9042 8482 9054
rect 8430 8978 8482 8990
rect 8766 9042 8818 9054
rect 8766 8978 8818 8990
rect 8990 9042 9042 9054
rect 13694 9042 13746 9054
rect 11106 8990 11118 9042
rect 11170 8990 11182 9042
rect 11554 8990 11566 9042
rect 11618 8990 11630 9042
rect 8990 8978 9042 8990
rect 13694 8978 13746 8990
rect 14030 9042 14082 9054
rect 14030 8978 14082 8990
rect 14366 9042 14418 9054
rect 14366 8978 14418 8990
rect 8878 8930 8930 8942
rect 3714 8878 3726 8930
rect 3778 8878 3790 8930
rect 5842 8878 5854 8930
rect 5906 8878 5918 8930
rect 8878 8866 8930 8878
rect 11342 8930 11394 8942
rect 11342 8866 11394 8878
rect 14142 8930 14194 8942
rect 14142 8866 14194 8878
rect 14702 8930 14754 8942
rect 14702 8866 14754 8878
rect 20078 8930 20130 8942
rect 20078 8866 20130 8878
rect 20526 8930 20578 8942
rect 20526 8866 20578 8878
rect 21086 8930 21138 8942
rect 21086 8866 21138 8878
rect 21534 8930 21586 8942
rect 21534 8866 21586 8878
rect 22318 8930 22370 8942
rect 22318 8866 22370 8878
rect 3278 8818 3330 8830
rect 20850 8766 20862 8818
rect 20914 8815 20926 8818
rect 21410 8815 21422 8818
rect 20914 8769 21422 8815
rect 20914 8766 20926 8769
rect 21410 8766 21422 8769
rect 21474 8766 21486 8818
rect 3278 8754 3330 8766
rect 1344 8650 22624 8684
rect 1344 8598 3874 8650
rect 3926 8598 3978 8650
rect 4030 8598 4082 8650
rect 4134 8598 9194 8650
rect 9246 8598 9298 8650
rect 9350 8598 9402 8650
rect 9454 8598 14514 8650
rect 14566 8598 14618 8650
rect 14670 8598 14722 8650
rect 14774 8598 19834 8650
rect 19886 8598 19938 8650
rect 19990 8598 20042 8650
rect 20094 8598 22624 8650
rect 1344 8564 22624 8598
rect 7086 8370 7138 8382
rect 14242 8318 14254 8370
rect 14306 8318 14318 8370
rect 16370 8318 16382 8370
rect 16434 8318 16446 8370
rect 7086 8306 7138 8318
rect 3490 8206 3502 8258
rect 3554 8206 3566 8258
rect 4162 8206 4174 8258
rect 4226 8206 4238 8258
rect 4834 8206 4846 8258
rect 4898 8206 4910 8258
rect 5730 8206 5742 8258
rect 5794 8206 5806 8258
rect 7858 8206 7870 8258
rect 7922 8206 7934 8258
rect 9874 8206 9886 8258
rect 9938 8206 9950 8258
rect 12562 8206 12574 8258
rect 12626 8206 12638 8258
rect 13458 8206 13470 8258
rect 13522 8206 13534 8258
rect 5966 8146 6018 8158
rect 5966 8082 6018 8094
rect 6302 8146 6354 8158
rect 6302 8082 6354 8094
rect 6638 8146 6690 8158
rect 10446 8146 10498 8158
rect 7970 8094 7982 8146
rect 8034 8094 8046 8146
rect 6638 8082 6690 8094
rect 10446 8082 10498 8094
rect 21758 8146 21810 8158
rect 21758 8082 21810 8094
rect 1822 8034 1874 8046
rect 2718 8034 2770 8046
rect 5070 8034 5122 8046
rect 2146 7982 2158 8034
rect 2210 7982 2222 8034
rect 3042 7982 3054 8034
rect 3106 7982 3118 8034
rect 3714 7982 3726 8034
rect 3778 7982 3790 8034
rect 4386 7982 4398 8034
rect 4450 7982 4462 8034
rect 1822 7970 1874 7982
rect 2718 7970 2770 7982
rect 5070 7970 5122 7982
rect 6974 8034 7026 8046
rect 6974 7970 7026 7982
rect 7198 8034 7250 8046
rect 7198 7970 7250 7982
rect 7422 8034 7474 8046
rect 12350 8034 12402 8046
rect 9986 7982 9998 8034
rect 10050 7982 10062 8034
rect 7422 7970 7474 7982
rect 12350 7970 12402 7982
rect 16830 8034 16882 8046
rect 16830 7970 16882 7982
rect 17390 8034 17442 8046
rect 17390 7970 17442 7982
rect 18062 8034 18114 8046
rect 18062 7970 18114 7982
rect 18510 8034 18562 8046
rect 18510 7970 18562 7982
rect 19070 8034 19122 8046
rect 19070 7970 19122 7982
rect 19518 8034 19570 8046
rect 19518 7970 19570 7982
rect 19854 8034 19906 8046
rect 19854 7970 19906 7982
rect 20414 8034 20466 8046
rect 20414 7970 20466 7982
rect 20750 8034 20802 8046
rect 20750 7970 20802 7982
rect 21422 8034 21474 8046
rect 21422 7970 21474 7982
rect 22206 8034 22258 8046
rect 22206 7970 22258 7982
rect 1344 7866 22784 7900
rect 1344 7814 6534 7866
rect 6586 7814 6638 7866
rect 6690 7814 6742 7866
rect 6794 7814 11854 7866
rect 11906 7814 11958 7866
rect 12010 7814 12062 7866
rect 12114 7814 17174 7866
rect 17226 7814 17278 7866
rect 17330 7814 17382 7866
rect 17434 7814 22494 7866
rect 22546 7814 22598 7866
rect 22650 7814 22702 7866
rect 22754 7814 22784 7866
rect 1344 7780 22784 7814
rect 2046 7698 2098 7710
rect 2046 7634 2098 7646
rect 2718 7698 2770 7710
rect 2718 7634 2770 7646
rect 4062 7698 4114 7710
rect 11106 7646 11118 7698
rect 11170 7646 11182 7698
rect 4062 7634 4114 7646
rect 3390 7586 3442 7598
rect 3390 7522 3442 7534
rect 4622 7586 4674 7598
rect 4622 7522 4674 7534
rect 6302 7586 6354 7598
rect 6302 7522 6354 7534
rect 8318 7586 8370 7598
rect 12126 7586 12178 7598
rect 9538 7534 9550 7586
rect 9602 7534 9614 7586
rect 8318 7522 8370 7534
rect 12126 7522 12178 7534
rect 18622 7586 18674 7598
rect 18622 7522 18674 7534
rect 20414 7586 20466 7598
rect 20414 7522 20466 7534
rect 20862 7586 20914 7598
rect 20862 7522 20914 7534
rect 21198 7586 21250 7598
rect 21198 7522 21250 7534
rect 21534 7586 21586 7598
rect 21534 7522 21586 7534
rect 21870 7586 21922 7598
rect 21870 7522 21922 7534
rect 1710 7474 1762 7486
rect 1710 7410 1762 7422
rect 2382 7474 2434 7486
rect 8878 7474 8930 7486
rect 3042 7422 3054 7474
rect 3106 7422 3118 7474
rect 3826 7422 3838 7474
rect 3890 7422 3902 7474
rect 6738 7422 6750 7474
rect 6802 7422 6814 7474
rect 2382 7410 2434 7422
rect 8878 7410 8930 7422
rect 11230 7474 11282 7486
rect 17278 7474 17330 7486
rect 13346 7422 13358 7474
rect 13410 7422 13422 7474
rect 16482 7422 16494 7474
rect 16546 7422 16558 7474
rect 11230 7410 11282 7422
rect 17278 7410 17330 7422
rect 17614 7474 17666 7486
rect 17614 7410 17666 7422
rect 17838 7474 17890 7486
rect 20078 7474 20130 7486
rect 18386 7422 18398 7474
rect 18450 7422 18462 7474
rect 17838 7410 17890 7422
rect 20078 7410 20130 7422
rect 22206 7474 22258 7486
rect 22206 7410 22258 7422
rect 17502 7362 17554 7374
rect 7970 7310 7982 7362
rect 8034 7310 8046 7362
rect 13682 7310 13694 7362
rect 13746 7310 13758 7362
rect 15810 7310 15822 7362
rect 15874 7310 15886 7362
rect 17502 7298 17554 7310
rect 19070 7362 19122 7374
rect 19070 7298 19122 7310
rect 19518 7362 19570 7374
rect 19518 7298 19570 7310
rect 3054 7250 3106 7262
rect 20750 7250 20802 7262
rect 19394 7198 19406 7250
rect 19458 7247 19470 7250
rect 19842 7247 19854 7250
rect 19458 7201 19854 7247
rect 19458 7198 19470 7201
rect 19842 7198 19854 7201
rect 19906 7198 19918 7250
rect 3054 7186 3106 7198
rect 20750 7186 20802 7198
rect 1344 7082 22624 7116
rect 1344 7030 3874 7082
rect 3926 7030 3978 7082
rect 4030 7030 4082 7082
rect 4134 7030 9194 7082
rect 9246 7030 9298 7082
rect 9350 7030 9402 7082
rect 9454 7030 14514 7082
rect 14566 7030 14618 7082
rect 14670 7030 14722 7082
rect 14774 7030 19834 7082
rect 19886 7030 19938 7082
rect 19990 7030 20042 7082
rect 20094 7030 22624 7082
rect 1344 6996 22624 7030
rect 2146 6750 2158 6802
rect 2210 6750 2222 6802
rect 16482 6750 16494 6802
rect 16546 6750 16558 6802
rect 5966 6690 6018 6702
rect 5058 6638 5070 6690
rect 5122 6638 5134 6690
rect 5966 6626 6018 6638
rect 6414 6690 6466 6702
rect 12798 6690 12850 6702
rect 6738 6638 6750 6690
rect 6802 6638 6814 6690
rect 12338 6638 12350 6690
rect 12402 6638 12414 6690
rect 13458 6638 13470 6690
rect 13522 6638 13534 6690
rect 19282 6638 19294 6690
rect 19346 6638 19358 6690
rect 19954 6638 19966 6690
rect 20018 6638 20030 6690
rect 6414 6626 6466 6638
rect 12798 6626 12850 6638
rect 5630 6578 5682 6590
rect 4274 6526 4286 6578
rect 4338 6526 4350 6578
rect 5630 6514 5682 6526
rect 6190 6578 6242 6590
rect 12686 6578 12738 6590
rect 7298 6526 7310 6578
rect 7362 6526 7374 6578
rect 6190 6514 6242 6526
rect 12686 6514 12738 6526
rect 19742 6578 19794 6590
rect 19742 6514 19794 6526
rect 20414 6578 20466 6590
rect 20414 6514 20466 6526
rect 21310 6578 21362 6590
rect 21310 6514 21362 6526
rect 22094 6578 22146 6590
rect 22094 6514 22146 6526
rect 1710 6466 1762 6478
rect 1710 6402 1762 6414
rect 5742 6466 5794 6478
rect 5742 6402 5794 6414
rect 6302 6466 6354 6478
rect 6302 6402 6354 6414
rect 19070 6466 19122 6478
rect 19070 6402 19122 6414
rect 20750 6466 20802 6478
rect 20750 6402 20802 6414
rect 21646 6466 21698 6478
rect 21646 6402 21698 6414
rect 1344 6298 22784 6332
rect 1344 6246 6534 6298
rect 6586 6246 6638 6298
rect 6690 6246 6742 6298
rect 6794 6246 11854 6298
rect 11906 6246 11958 6298
rect 12010 6246 12062 6298
rect 12114 6246 17174 6298
rect 17226 6246 17278 6298
rect 17330 6246 17382 6298
rect 17434 6246 22494 6298
rect 22546 6246 22598 6298
rect 22650 6246 22702 6298
rect 22754 6246 22784 6298
rect 1344 6212 22784 6246
rect 2046 6130 2098 6142
rect 3502 6130 3554 6142
rect 2818 6078 2830 6130
rect 2882 6078 2894 6130
rect 2046 6066 2098 6078
rect 3502 6066 3554 6078
rect 9550 6130 9602 6142
rect 9550 6066 9602 6078
rect 16494 6130 16546 6142
rect 16494 6066 16546 6078
rect 17390 6130 17442 6142
rect 17390 6066 17442 6078
rect 17502 6130 17554 6142
rect 17502 6066 17554 6078
rect 17614 6130 17666 6142
rect 17614 6066 17666 6078
rect 1934 6018 1986 6030
rect 4734 6018 4786 6030
rect 4162 5966 4174 6018
rect 4226 5966 4238 6018
rect 1934 5954 1986 5966
rect 4734 5954 4786 5966
rect 6302 6018 6354 6030
rect 6302 5954 6354 5966
rect 7758 6018 7810 6030
rect 10334 6018 10386 6030
rect 17838 6018 17890 6030
rect 21534 6018 21586 6030
rect 10098 5966 10110 6018
rect 10162 5966 10174 6018
rect 13458 5966 13470 6018
rect 13522 5966 13534 6018
rect 20402 5966 20414 6018
rect 20466 5966 20478 6018
rect 7758 5954 7810 5966
rect 10334 5954 10386 5966
rect 17838 5954 17890 5966
rect 21534 5954 21586 5966
rect 6862 5906 6914 5918
rect 2594 5854 2606 5906
rect 2658 5854 2670 5906
rect 3266 5854 3278 5906
rect 3330 5854 3342 5906
rect 3938 5854 3950 5906
rect 4002 5854 4014 5906
rect 7186 5854 7198 5906
rect 7250 5854 7262 5906
rect 9538 5854 9550 5906
rect 9602 5854 9614 5906
rect 16146 5854 16158 5906
rect 16210 5854 16222 5906
rect 16706 5854 16718 5906
rect 16770 5854 16782 5906
rect 21186 5854 21198 5906
rect 21250 5854 21262 5906
rect 21746 5854 21758 5906
rect 21810 5854 21822 5906
rect 6862 5842 6914 5854
rect 2158 5794 2210 5806
rect 4834 5742 4846 5794
rect 4898 5742 4910 5794
rect 8306 5742 8318 5794
rect 8370 5742 8382 5794
rect 18274 5742 18286 5794
rect 18338 5742 18350 5794
rect 2158 5730 2210 5742
rect 4510 5682 4562 5694
rect 4510 5618 4562 5630
rect 9886 5682 9938 5694
rect 9886 5618 9938 5630
rect 1344 5514 22624 5548
rect 1344 5462 3874 5514
rect 3926 5462 3978 5514
rect 4030 5462 4082 5514
rect 4134 5462 9194 5514
rect 9246 5462 9298 5514
rect 9350 5462 9402 5514
rect 9454 5462 14514 5514
rect 14566 5462 14618 5514
rect 14670 5462 14722 5514
rect 14774 5462 19834 5514
rect 19886 5462 19938 5514
rect 19990 5462 20042 5514
rect 20094 5462 22624 5514
rect 1344 5428 22624 5462
rect 13582 5234 13634 5246
rect 5842 5182 5854 5234
rect 5906 5182 5918 5234
rect 7970 5182 7982 5234
rect 8034 5182 8046 5234
rect 13582 5170 13634 5182
rect 21422 5234 21474 5246
rect 21422 5170 21474 5182
rect 22094 5234 22146 5246
rect 22094 5170 22146 5182
rect 4622 5122 4674 5134
rect 2370 5070 2382 5122
rect 2434 5070 2446 5122
rect 3266 5070 3278 5122
rect 3330 5070 3342 5122
rect 3938 5070 3950 5122
rect 4002 5070 4014 5122
rect 4622 5058 4674 5070
rect 5182 5122 5234 5134
rect 12798 5122 12850 5134
rect 19070 5122 19122 5134
rect 8642 5070 8654 5122
rect 8706 5070 8718 5122
rect 10658 5070 10670 5122
rect 10722 5070 10734 5122
rect 14018 5070 14030 5122
rect 14082 5070 14094 5122
rect 16370 5070 16382 5122
rect 16434 5070 16446 5122
rect 16818 5070 16830 5122
rect 16882 5070 16894 5122
rect 5182 5058 5234 5070
rect 12798 5058 12850 5070
rect 19070 5058 19122 5070
rect 19742 5122 19794 5134
rect 19742 5058 19794 5070
rect 20078 5122 20130 5134
rect 20078 5058 20130 5070
rect 21310 5122 21362 5134
rect 21310 5058 21362 5070
rect 4734 5010 4786 5022
rect 4734 4946 4786 4958
rect 9662 5010 9714 5022
rect 15822 5010 15874 5022
rect 18734 5010 18786 5022
rect 12898 4958 12910 5010
rect 12962 4958 12974 5010
rect 18386 4958 18398 5010
rect 18450 4958 18462 5010
rect 9662 4946 9714 4958
rect 15822 4946 15874 4958
rect 18734 4946 18786 4958
rect 19406 5010 19458 5022
rect 19406 4946 19458 4958
rect 20414 5010 20466 5022
rect 20414 4946 20466 4958
rect 21534 5010 21586 5022
rect 21534 4946 21586 4958
rect 21982 5010 22034 5022
rect 21982 4946 22034 4958
rect 1710 4898 1762 4910
rect 1710 4834 1762 4846
rect 3502 4898 3554 4910
rect 3502 4834 3554 4846
rect 4174 4898 4226 4910
rect 4174 4834 4226 4846
rect 4958 4898 5010 4910
rect 13470 4898 13522 4910
rect 12786 4846 12798 4898
rect 12850 4846 12862 4898
rect 4958 4834 5010 4846
rect 13470 4834 13522 4846
rect 13694 4898 13746 4910
rect 14802 4846 14814 4898
rect 14866 4846 14878 4898
rect 13694 4834 13746 4846
rect 1344 4730 22784 4764
rect 1344 4678 6534 4730
rect 6586 4678 6638 4730
rect 6690 4678 6742 4730
rect 6794 4678 11854 4730
rect 11906 4678 11958 4730
rect 12010 4678 12062 4730
rect 12114 4678 17174 4730
rect 17226 4678 17278 4730
rect 17330 4678 17382 4730
rect 17434 4678 22494 4730
rect 22546 4678 22598 4730
rect 22650 4678 22702 4730
rect 22754 4678 22784 4730
rect 1344 4644 22784 4678
rect 9438 4562 9490 4574
rect 8866 4510 8878 4562
rect 8930 4510 8942 4562
rect 9438 4498 9490 4510
rect 9662 4562 9714 4574
rect 9662 4498 9714 4510
rect 9774 4450 9826 4462
rect 14254 4450 14306 4462
rect 18062 4450 18114 4462
rect 4050 4398 4062 4450
rect 4114 4398 4126 4450
rect 5282 4398 5294 4450
rect 5346 4398 5358 4450
rect 8978 4398 8990 4450
rect 9042 4398 9054 4450
rect 10658 4398 10670 4450
rect 10722 4398 10734 4450
rect 16706 4398 16718 4450
rect 16770 4398 16782 4450
rect 21074 4398 21086 4450
rect 21138 4398 21150 4450
rect 21858 4398 21870 4450
rect 21922 4398 21934 4450
rect 9774 4386 9826 4398
rect 14254 4386 14306 4398
rect 18062 4386 18114 4398
rect 7310 4338 7362 4350
rect 15150 4338 15202 4350
rect 4834 4286 4846 4338
rect 4898 4286 4910 4338
rect 6962 4286 6974 4338
rect 7026 4286 7038 4338
rect 11330 4286 11342 4338
rect 11394 4286 11406 4338
rect 11778 4286 11790 4338
rect 11842 4286 11854 4338
rect 13010 4286 13022 4338
rect 13074 4286 13086 4338
rect 7310 4274 7362 4286
rect 15150 4274 15202 4286
rect 17502 4338 17554 4350
rect 17502 4274 17554 4286
rect 19518 4338 19570 4350
rect 21634 4286 21646 4338
rect 21698 4286 21710 4338
rect 19518 4274 19570 4286
rect 1922 4174 1934 4226
rect 1986 4174 1998 4226
rect 10210 4174 10222 4226
rect 10274 4174 10286 4226
rect 14130 4174 14142 4226
rect 14194 4174 14206 4226
rect 19282 4174 19294 4226
rect 19346 4174 19358 4226
rect 1344 3946 22624 3980
rect 1344 3894 3874 3946
rect 3926 3894 3978 3946
rect 4030 3894 4082 3946
rect 4134 3894 9194 3946
rect 9246 3894 9298 3946
rect 9350 3894 9402 3946
rect 9454 3894 14514 3946
rect 14566 3894 14618 3946
rect 14670 3894 14722 3946
rect 14774 3894 19834 3946
rect 19886 3894 19938 3946
rect 19990 3894 20042 3946
rect 20094 3894 22624 3946
rect 1344 3860 22624 3894
rect 1934 3778 1986 3790
rect 1934 3714 1986 3726
rect 4510 3778 4562 3790
rect 4510 3714 4562 3726
rect 6974 3778 7026 3790
rect 6974 3714 7026 3726
rect 13246 3778 13298 3790
rect 16158 3778 16210 3790
rect 13794 3726 13806 3778
rect 13858 3726 13870 3778
rect 13246 3714 13298 3726
rect 16158 3714 16210 3726
rect 4846 3666 4898 3678
rect 4846 3602 4898 3614
rect 7086 3666 7138 3678
rect 16270 3666 16322 3678
rect 7746 3614 7758 3666
rect 7810 3614 7822 3666
rect 10546 3614 10558 3666
rect 10610 3614 10622 3666
rect 7086 3602 7138 3614
rect 16270 3602 16322 3614
rect 22206 3666 22258 3678
rect 22206 3602 22258 3614
rect 2718 3554 2770 3566
rect 4958 3554 5010 3566
rect 7422 3554 7474 3566
rect 13134 3554 13186 3566
rect 16830 3554 16882 3566
rect 3714 3502 3726 3554
rect 3778 3502 3790 3554
rect 4274 3502 4286 3554
rect 4338 3502 4350 3554
rect 5618 3502 5630 3554
rect 5682 3502 5694 3554
rect 7858 3502 7870 3554
rect 7922 3502 7934 3554
rect 8082 3502 8094 3554
rect 8146 3502 8158 3554
rect 9986 3502 9998 3554
rect 10050 3502 10062 3554
rect 10994 3502 11006 3554
rect 11058 3502 11070 3554
rect 14914 3502 14926 3554
rect 14978 3502 14990 3554
rect 15698 3502 15710 3554
rect 15762 3502 15774 3554
rect 16930 3502 16942 3554
rect 16994 3502 17006 3554
rect 19170 3502 19182 3554
rect 19234 3502 19246 3554
rect 20962 3502 20974 3554
rect 21026 3502 21038 3554
rect 21634 3502 21646 3554
rect 21698 3502 21710 3554
rect 2718 3490 2770 3502
rect 4958 3490 5010 3502
rect 7422 3490 7474 3502
rect 13134 3490 13186 3502
rect 16830 3490 16882 3502
rect 3054 3442 3106 3454
rect 15486 3442 15538 3454
rect 20750 3442 20802 3454
rect 4722 3390 4734 3442
rect 4786 3390 4798 3442
rect 5730 3390 5742 3442
rect 5794 3390 5806 3442
rect 6178 3390 6190 3442
rect 6242 3390 6254 3442
rect 9874 3390 9886 3442
rect 9938 3390 9950 3442
rect 10882 3390 10894 3442
rect 10946 3390 10958 3442
rect 14130 3390 14142 3442
rect 14194 3390 14206 3442
rect 18386 3390 18398 3442
rect 18450 3390 18462 3442
rect 19282 3390 19294 3442
rect 19346 3390 19358 3442
rect 3054 3378 3106 3390
rect 15486 3378 15538 3390
rect 20750 3378 20802 3390
rect 21422 3442 21474 3454
rect 21422 3378 21474 3390
rect 13246 3330 13298 3342
rect 6402 3278 6414 3330
rect 6466 3278 6478 3330
rect 13246 3266 13298 3278
rect 1344 3162 22784 3196
rect 1344 3110 6534 3162
rect 6586 3110 6638 3162
rect 6690 3110 6742 3162
rect 6794 3110 11854 3162
rect 11906 3110 11958 3162
rect 12010 3110 12062 3162
rect 12114 3110 17174 3162
rect 17226 3110 17278 3162
rect 17330 3110 17382 3162
rect 17434 3110 22494 3162
rect 22546 3110 22598 3162
rect 22650 3110 22702 3162
rect 22754 3110 22784 3162
rect 1344 3076 22784 3110
rect 3266 2942 3278 2994
rect 3330 2991 3342 2994
rect 8642 2991 8654 2994
rect 3330 2945 8654 2991
rect 3330 2942 3342 2945
rect 8642 2942 8654 2945
rect 8706 2942 8718 2994
rect 20178 2942 20190 2994
rect 20242 2991 20254 2994
rect 21746 2991 21758 2994
rect 20242 2945 21758 2991
rect 20242 2942 20254 2945
rect 21746 2942 21758 2945
rect 21810 2942 21822 2994
rect 1586 2830 1598 2882
rect 1650 2879 1662 2882
rect 4946 2879 4958 2882
rect 1650 2833 4958 2879
rect 1650 2830 1662 2833
rect 4946 2830 4958 2833
rect 5010 2830 5022 2882
<< via1 >>
rect 3874 16438 3926 16490
rect 3978 16438 4030 16490
rect 4082 16438 4134 16490
rect 9194 16438 9246 16490
rect 9298 16438 9350 16490
rect 9402 16438 9454 16490
rect 14514 16438 14566 16490
rect 14618 16438 14670 16490
rect 14722 16438 14774 16490
rect 19834 16438 19886 16490
rect 19938 16438 19990 16490
rect 20042 16438 20094 16490
rect 1822 16270 1874 16322
rect 21758 16270 21810 16322
rect 7758 16158 7810 16210
rect 17054 16158 17106 16210
rect 8766 16046 8818 16098
rect 3838 15934 3890 15986
rect 4734 15934 4786 15986
rect 10558 15934 10610 15986
rect 13470 15934 13522 15986
rect 19294 15934 19346 15986
rect 2606 15822 2658 15874
rect 3390 15822 3442 15874
rect 9438 15822 9490 15874
rect 17726 15822 17778 15874
rect 20302 15822 20354 15874
rect 20974 15822 21026 15874
rect 6534 15654 6586 15706
rect 6638 15654 6690 15706
rect 6742 15654 6794 15706
rect 11854 15654 11906 15706
rect 11958 15654 12010 15706
rect 12062 15654 12114 15706
rect 17174 15654 17226 15706
rect 17278 15654 17330 15706
rect 17382 15654 17434 15706
rect 22494 15654 22546 15706
rect 22598 15654 22650 15706
rect 22702 15654 22754 15706
rect 2606 15486 2658 15538
rect 3054 15486 3106 15538
rect 3502 15486 3554 15538
rect 1710 15374 1762 15426
rect 2158 15374 2210 15426
rect 22206 15038 22258 15090
rect 3874 14870 3926 14922
rect 3978 14870 4030 14922
rect 4082 14870 4134 14922
rect 9194 14870 9246 14922
rect 9298 14870 9350 14922
rect 9402 14870 9454 14922
rect 14514 14870 14566 14922
rect 14618 14870 14670 14922
rect 14722 14870 14774 14922
rect 19834 14870 19886 14922
rect 19938 14870 19990 14922
rect 20042 14870 20094 14922
rect 1710 14254 1762 14306
rect 2158 14254 2210 14306
rect 6534 14086 6586 14138
rect 6638 14086 6690 14138
rect 6742 14086 6794 14138
rect 11854 14086 11906 14138
rect 11958 14086 12010 14138
rect 12062 14086 12114 14138
rect 17174 14086 17226 14138
rect 17278 14086 17330 14138
rect 17382 14086 17434 14138
rect 22494 14086 22546 14138
rect 22598 14086 22650 14138
rect 22702 14086 22754 14138
rect 1710 13806 1762 13858
rect 3874 13302 3926 13354
rect 3978 13302 4030 13354
rect 4082 13302 4134 13354
rect 9194 13302 9246 13354
rect 9298 13302 9350 13354
rect 9402 13302 9454 13354
rect 14514 13302 14566 13354
rect 14618 13302 14670 13354
rect 14722 13302 14774 13354
rect 19834 13302 19886 13354
rect 19938 13302 19990 13354
rect 20042 13302 20094 13354
rect 1710 12798 1762 12850
rect 22206 12798 22258 12850
rect 2158 12686 2210 12738
rect 21646 12686 21698 12738
rect 21870 12686 21922 12738
rect 6534 12518 6586 12570
rect 6638 12518 6690 12570
rect 6742 12518 6794 12570
rect 11854 12518 11906 12570
rect 11958 12518 12010 12570
rect 12062 12518 12114 12570
rect 17174 12518 17226 12570
rect 17278 12518 17330 12570
rect 17382 12518 17434 12570
rect 22494 12518 22546 12570
rect 22598 12518 22650 12570
rect 22702 12518 22754 12570
rect 1710 12238 1762 12290
rect 2158 12238 2210 12290
rect 3838 12126 3890 12178
rect 2830 12014 2882 12066
rect 3278 12014 3330 12066
rect 4286 12014 4338 12066
rect 3874 11734 3926 11786
rect 3978 11734 4030 11786
rect 4082 11734 4134 11786
rect 9194 11734 9246 11786
rect 9298 11734 9350 11786
rect 9402 11734 9454 11786
rect 14514 11734 14566 11786
rect 14618 11734 14670 11786
rect 14722 11734 14774 11786
rect 19834 11734 19886 11786
rect 19938 11734 19990 11786
rect 20042 11734 20094 11786
rect 4958 11454 5010 11506
rect 1710 11118 1762 11170
rect 2158 11118 2210 11170
rect 2830 11118 2882 11170
rect 3390 11118 3442 11170
rect 3726 11118 3778 11170
rect 4510 11118 4562 11170
rect 9998 11118 10050 11170
rect 6534 10950 6586 11002
rect 6638 10950 6690 11002
rect 6742 10950 6794 11002
rect 11854 10950 11906 11002
rect 11958 10950 12010 11002
rect 12062 10950 12114 11002
rect 17174 10950 17226 11002
rect 17278 10950 17330 11002
rect 17382 10950 17434 11002
rect 22494 10950 22546 11002
rect 22598 10950 22650 11002
rect 22702 10950 22754 11002
rect 1710 10670 1762 10722
rect 2158 10670 2210 10722
rect 2606 10670 2658 10722
rect 3054 10670 3106 10722
rect 10222 10670 10274 10722
rect 9998 10558 10050 10610
rect 11118 10558 11170 10610
rect 4062 10446 4114 10498
rect 4622 10446 4674 10498
rect 5182 10446 5234 10498
rect 5630 10446 5682 10498
rect 5966 10446 6018 10498
rect 6526 10446 6578 10498
rect 6974 10446 7026 10498
rect 8990 10446 9042 10498
rect 10670 10446 10722 10498
rect 11678 10446 11730 10498
rect 12126 10446 12178 10498
rect 5966 10334 6018 10386
rect 7086 10334 7138 10386
rect 10446 10334 10498 10386
rect 11006 10334 11058 10386
rect 3874 10166 3926 10218
rect 3978 10166 4030 10218
rect 4082 10166 4134 10218
rect 9194 10166 9246 10218
rect 9298 10166 9350 10218
rect 9402 10166 9454 10218
rect 14514 10166 14566 10218
rect 14618 10166 14670 10218
rect 14722 10166 14774 10218
rect 19834 10166 19886 10218
rect 19938 10166 19990 10218
rect 20042 10166 20094 10218
rect 9774 9774 9826 9826
rect 10782 9774 10834 9826
rect 11454 9774 11506 9826
rect 12238 9774 12290 9826
rect 4958 9662 5010 9714
rect 8654 9662 8706 9714
rect 1710 9550 1762 9602
rect 2158 9550 2210 9602
rect 2606 9550 2658 9602
rect 3054 9550 3106 9602
rect 3726 9550 3778 9602
rect 4174 9550 4226 9602
rect 4622 9550 4674 9602
rect 4846 9550 4898 9602
rect 5854 9550 5906 9602
rect 6302 9550 6354 9602
rect 6974 9550 7026 9602
rect 7422 9550 7474 9602
rect 7870 9550 7922 9602
rect 8430 9550 8482 9602
rect 8990 9550 9042 9602
rect 9998 9550 10050 9602
rect 10558 9550 10610 9602
rect 11230 9550 11282 9602
rect 11902 9550 11954 9602
rect 12686 9550 12738 9602
rect 20862 9550 20914 9602
rect 22206 9550 22258 9602
rect 6534 9382 6586 9434
rect 6638 9382 6690 9434
rect 6742 9382 6794 9434
rect 11854 9382 11906 9434
rect 11958 9382 12010 9434
rect 12062 9382 12114 9434
rect 17174 9382 17226 9434
rect 17278 9382 17330 9434
rect 17382 9382 17434 9434
rect 22494 9382 22546 9434
rect 22598 9382 22650 9434
rect 22702 9382 22754 9434
rect 15150 9214 15202 9266
rect 1822 9102 1874 9154
rect 2270 9102 2322 9154
rect 2718 9102 2770 9154
rect 3278 9102 3330 9154
rect 3390 9102 3442 9154
rect 7086 9102 7138 9154
rect 8094 9102 8146 9154
rect 10110 9102 10162 9154
rect 12126 9102 12178 9154
rect 6526 8990 6578 9042
rect 6862 8990 6914 9042
rect 7198 8990 7250 9042
rect 7758 8990 7810 9042
rect 8430 8990 8482 9042
rect 8766 8990 8818 9042
rect 8990 8990 9042 9042
rect 11118 8990 11170 9042
rect 11566 8990 11618 9042
rect 13694 8990 13746 9042
rect 14030 8990 14082 9042
rect 14366 8990 14418 9042
rect 3726 8878 3778 8930
rect 5854 8878 5906 8930
rect 8878 8878 8930 8930
rect 11342 8878 11394 8930
rect 14142 8878 14194 8930
rect 14702 8878 14754 8930
rect 20078 8878 20130 8930
rect 20526 8878 20578 8930
rect 21086 8878 21138 8930
rect 21534 8878 21586 8930
rect 22318 8878 22370 8930
rect 3278 8766 3330 8818
rect 20862 8766 20914 8818
rect 21422 8766 21474 8818
rect 3874 8598 3926 8650
rect 3978 8598 4030 8650
rect 4082 8598 4134 8650
rect 9194 8598 9246 8650
rect 9298 8598 9350 8650
rect 9402 8598 9454 8650
rect 14514 8598 14566 8650
rect 14618 8598 14670 8650
rect 14722 8598 14774 8650
rect 19834 8598 19886 8650
rect 19938 8598 19990 8650
rect 20042 8598 20094 8650
rect 7086 8318 7138 8370
rect 14254 8318 14306 8370
rect 16382 8318 16434 8370
rect 3502 8206 3554 8258
rect 4174 8206 4226 8258
rect 4846 8206 4898 8258
rect 5742 8206 5794 8258
rect 7870 8206 7922 8258
rect 9886 8206 9938 8258
rect 12574 8206 12626 8258
rect 13470 8206 13522 8258
rect 5966 8094 6018 8146
rect 6302 8094 6354 8146
rect 6638 8094 6690 8146
rect 7982 8094 8034 8146
rect 10446 8094 10498 8146
rect 21758 8094 21810 8146
rect 1822 7982 1874 8034
rect 2158 7982 2210 8034
rect 2718 7982 2770 8034
rect 3054 7982 3106 8034
rect 3726 7982 3778 8034
rect 4398 7982 4450 8034
rect 5070 7982 5122 8034
rect 6974 7982 7026 8034
rect 7198 7982 7250 8034
rect 7422 7982 7474 8034
rect 9998 7982 10050 8034
rect 12350 7982 12402 8034
rect 16830 7982 16882 8034
rect 17390 7982 17442 8034
rect 18062 7982 18114 8034
rect 18510 7982 18562 8034
rect 19070 7982 19122 8034
rect 19518 7982 19570 8034
rect 19854 7982 19906 8034
rect 20414 7982 20466 8034
rect 20750 7982 20802 8034
rect 21422 7982 21474 8034
rect 22206 7982 22258 8034
rect 6534 7814 6586 7866
rect 6638 7814 6690 7866
rect 6742 7814 6794 7866
rect 11854 7814 11906 7866
rect 11958 7814 12010 7866
rect 12062 7814 12114 7866
rect 17174 7814 17226 7866
rect 17278 7814 17330 7866
rect 17382 7814 17434 7866
rect 22494 7814 22546 7866
rect 22598 7814 22650 7866
rect 22702 7814 22754 7866
rect 2046 7646 2098 7698
rect 2718 7646 2770 7698
rect 4062 7646 4114 7698
rect 11118 7646 11170 7698
rect 3390 7534 3442 7586
rect 4622 7534 4674 7586
rect 6302 7534 6354 7586
rect 8318 7534 8370 7586
rect 9550 7534 9602 7586
rect 12126 7534 12178 7586
rect 18622 7534 18674 7586
rect 20414 7534 20466 7586
rect 20862 7534 20914 7586
rect 21198 7534 21250 7586
rect 21534 7534 21586 7586
rect 21870 7534 21922 7586
rect 1710 7422 1762 7474
rect 2382 7422 2434 7474
rect 3054 7422 3106 7474
rect 3838 7422 3890 7474
rect 6750 7422 6802 7474
rect 8878 7422 8930 7474
rect 11230 7422 11282 7474
rect 13358 7422 13410 7474
rect 16494 7422 16546 7474
rect 17278 7422 17330 7474
rect 17614 7422 17666 7474
rect 17838 7422 17890 7474
rect 18398 7422 18450 7474
rect 20078 7422 20130 7474
rect 22206 7422 22258 7474
rect 7982 7310 8034 7362
rect 13694 7310 13746 7362
rect 15822 7310 15874 7362
rect 17502 7310 17554 7362
rect 19070 7310 19122 7362
rect 19518 7310 19570 7362
rect 3054 7198 3106 7250
rect 19406 7198 19458 7250
rect 19854 7198 19906 7250
rect 20750 7198 20802 7250
rect 3874 7030 3926 7082
rect 3978 7030 4030 7082
rect 4082 7030 4134 7082
rect 9194 7030 9246 7082
rect 9298 7030 9350 7082
rect 9402 7030 9454 7082
rect 14514 7030 14566 7082
rect 14618 7030 14670 7082
rect 14722 7030 14774 7082
rect 19834 7030 19886 7082
rect 19938 7030 19990 7082
rect 20042 7030 20094 7082
rect 2158 6750 2210 6802
rect 16494 6750 16546 6802
rect 5070 6638 5122 6690
rect 5966 6638 6018 6690
rect 6414 6638 6466 6690
rect 6750 6638 6802 6690
rect 12350 6638 12402 6690
rect 12798 6638 12850 6690
rect 13470 6638 13522 6690
rect 19294 6638 19346 6690
rect 19966 6638 20018 6690
rect 4286 6526 4338 6578
rect 5630 6526 5682 6578
rect 6190 6526 6242 6578
rect 7310 6526 7362 6578
rect 12686 6526 12738 6578
rect 19742 6526 19794 6578
rect 20414 6526 20466 6578
rect 21310 6526 21362 6578
rect 22094 6526 22146 6578
rect 1710 6414 1762 6466
rect 5742 6414 5794 6466
rect 6302 6414 6354 6466
rect 19070 6414 19122 6466
rect 20750 6414 20802 6466
rect 21646 6414 21698 6466
rect 6534 6246 6586 6298
rect 6638 6246 6690 6298
rect 6742 6246 6794 6298
rect 11854 6246 11906 6298
rect 11958 6246 12010 6298
rect 12062 6246 12114 6298
rect 17174 6246 17226 6298
rect 17278 6246 17330 6298
rect 17382 6246 17434 6298
rect 22494 6246 22546 6298
rect 22598 6246 22650 6298
rect 22702 6246 22754 6298
rect 2046 6078 2098 6130
rect 2830 6078 2882 6130
rect 3502 6078 3554 6130
rect 9550 6078 9602 6130
rect 16494 6078 16546 6130
rect 17390 6078 17442 6130
rect 17502 6078 17554 6130
rect 17614 6078 17666 6130
rect 1934 5966 1986 6018
rect 4174 5966 4226 6018
rect 4734 5966 4786 6018
rect 6302 5966 6354 6018
rect 7758 5966 7810 6018
rect 10110 5966 10162 6018
rect 10334 5966 10386 6018
rect 13470 5966 13522 6018
rect 17838 5966 17890 6018
rect 20414 5966 20466 6018
rect 21534 5966 21586 6018
rect 2606 5854 2658 5906
rect 3278 5854 3330 5906
rect 3950 5854 4002 5906
rect 6862 5854 6914 5906
rect 7198 5854 7250 5906
rect 9550 5854 9602 5906
rect 16158 5854 16210 5906
rect 16718 5854 16770 5906
rect 21198 5854 21250 5906
rect 21758 5854 21810 5906
rect 2158 5742 2210 5794
rect 4846 5742 4898 5794
rect 8318 5742 8370 5794
rect 18286 5742 18338 5794
rect 4510 5630 4562 5682
rect 9886 5630 9938 5682
rect 3874 5462 3926 5514
rect 3978 5462 4030 5514
rect 4082 5462 4134 5514
rect 9194 5462 9246 5514
rect 9298 5462 9350 5514
rect 9402 5462 9454 5514
rect 14514 5462 14566 5514
rect 14618 5462 14670 5514
rect 14722 5462 14774 5514
rect 19834 5462 19886 5514
rect 19938 5462 19990 5514
rect 20042 5462 20094 5514
rect 5854 5182 5906 5234
rect 7982 5182 8034 5234
rect 13582 5182 13634 5234
rect 21422 5182 21474 5234
rect 22094 5182 22146 5234
rect 2382 5070 2434 5122
rect 3278 5070 3330 5122
rect 3950 5070 4002 5122
rect 4622 5070 4674 5122
rect 5182 5070 5234 5122
rect 8654 5070 8706 5122
rect 10670 5070 10722 5122
rect 12798 5070 12850 5122
rect 14030 5070 14082 5122
rect 16382 5070 16434 5122
rect 16830 5070 16882 5122
rect 19070 5070 19122 5122
rect 19742 5070 19794 5122
rect 20078 5070 20130 5122
rect 21310 5070 21362 5122
rect 4734 4958 4786 5010
rect 9662 4958 9714 5010
rect 12910 4958 12962 5010
rect 15822 4958 15874 5010
rect 18398 4958 18450 5010
rect 18734 4958 18786 5010
rect 19406 4958 19458 5010
rect 20414 4958 20466 5010
rect 21534 4958 21586 5010
rect 21982 4958 22034 5010
rect 1710 4846 1762 4898
rect 3502 4846 3554 4898
rect 4174 4846 4226 4898
rect 4958 4846 5010 4898
rect 12798 4846 12850 4898
rect 13470 4846 13522 4898
rect 13694 4846 13746 4898
rect 14814 4846 14866 4898
rect 6534 4678 6586 4730
rect 6638 4678 6690 4730
rect 6742 4678 6794 4730
rect 11854 4678 11906 4730
rect 11958 4678 12010 4730
rect 12062 4678 12114 4730
rect 17174 4678 17226 4730
rect 17278 4678 17330 4730
rect 17382 4678 17434 4730
rect 22494 4678 22546 4730
rect 22598 4678 22650 4730
rect 22702 4678 22754 4730
rect 8878 4510 8930 4562
rect 9438 4510 9490 4562
rect 9662 4510 9714 4562
rect 4062 4398 4114 4450
rect 5294 4398 5346 4450
rect 8990 4398 9042 4450
rect 9774 4398 9826 4450
rect 10670 4398 10722 4450
rect 14254 4398 14306 4450
rect 16718 4398 16770 4450
rect 18062 4398 18114 4450
rect 21086 4398 21138 4450
rect 21870 4398 21922 4450
rect 4846 4286 4898 4338
rect 6974 4286 7026 4338
rect 7310 4286 7362 4338
rect 11342 4286 11394 4338
rect 11790 4286 11842 4338
rect 13022 4286 13074 4338
rect 15150 4286 15202 4338
rect 17502 4286 17554 4338
rect 19518 4286 19570 4338
rect 21646 4286 21698 4338
rect 1934 4174 1986 4226
rect 10222 4174 10274 4226
rect 14142 4174 14194 4226
rect 19294 4174 19346 4226
rect 3874 3894 3926 3946
rect 3978 3894 4030 3946
rect 4082 3894 4134 3946
rect 9194 3894 9246 3946
rect 9298 3894 9350 3946
rect 9402 3894 9454 3946
rect 14514 3894 14566 3946
rect 14618 3894 14670 3946
rect 14722 3894 14774 3946
rect 19834 3894 19886 3946
rect 19938 3894 19990 3946
rect 20042 3894 20094 3946
rect 1934 3726 1986 3778
rect 4510 3726 4562 3778
rect 6974 3726 7026 3778
rect 13246 3726 13298 3778
rect 13806 3726 13858 3778
rect 16158 3726 16210 3778
rect 4846 3614 4898 3666
rect 7086 3614 7138 3666
rect 7758 3614 7810 3666
rect 10558 3614 10610 3666
rect 16270 3614 16322 3666
rect 22206 3614 22258 3666
rect 2718 3502 2770 3554
rect 3726 3502 3778 3554
rect 4286 3502 4338 3554
rect 4958 3502 5010 3554
rect 5630 3502 5682 3554
rect 7422 3502 7474 3554
rect 7870 3502 7922 3554
rect 8094 3502 8146 3554
rect 9998 3502 10050 3554
rect 11006 3502 11058 3554
rect 13134 3502 13186 3554
rect 14926 3502 14978 3554
rect 15710 3502 15762 3554
rect 16830 3502 16882 3554
rect 16942 3502 16994 3554
rect 19182 3502 19234 3554
rect 20974 3502 21026 3554
rect 21646 3502 21698 3554
rect 3054 3390 3106 3442
rect 4734 3390 4786 3442
rect 5742 3390 5794 3442
rect 6190 3390 6242 3442
rect 9886 3390 9938 3442
rect 10894 3390 10946 3442
rect 14142 3390 14194 3442
rect 15486 3390 15538 3442
rect 18398 3390 18450 3442
rect 19294 3390 19346 3442
rect 20750 3390 20802 3442
rect 21422 3390 21474 3442
rect 6414 3278 6466 3330
rect 13246 3278 13298 3330
rect 6534 3110 6586 3162
rect 6638 3110 6690 3162
rect 6742 3110 6794 3162
rect 11854 3110 11906 3162
rect 11958 3110 12010 3162
rect 12062 3110 12114 3162
rect 17174 3110 17226 3162
rect 17278 3110 17330 3162
rect 17382 3110 17434 3162
rect 22494 3110 22546 3162
rect 22598 3110 22650 3162
rect 22702 3110 22754 3162
rect 3278 2942 3330 2994
rect 8654 2942 8706 2994
rect 20190 2942 20242 2994
rect 21758 2942 21810 2994
rect 1598 2830 1650 2882
rect 4958 2830 5010 2882
<< metal2 >>
rect 1568 19200 1680 20000
rect 4480 19200 4592 20000
rect 7392 19200 7504 20000
rect 10304 19200 10416 20000
rect 13216 19200 13328 20000
rect 16128 19200 16240 20000
rect 19040 19200 19152 20000
rect 21952 19200 22064 20000
rect 1596 16324 1652 19200
rect 3500 17332 3556 17342
rect 3052 16436 3108 16446
rect 1820 16324 1876 16334
rect 1596 16322 1876 16324
rect 1596 16270 1822 16322
rect 1874 16270 1876 16322
rect 1596 16268 1876 16270
rect 1820 16258 1876 16268
rect 2380 15988 2436 15998
rect 2436 15932 2548 15988
rect 2380 15922 2436 15932
rect 2492 15540 2548 15932
rect 2604 15876 2660 15886
rect 2604 15874 2772 15876
rect 2604 15822 2606 15874
rect 2658 15822 2772 15874
rect 2604 15820 2772 15822
rect 2604 15810 2660 15820
rect 2604 15540 2660 15550
rect 2492 15538 2660 15540
rect 2492 15486 2606 15538
rect 2658 15486 2660 15538
rect 2492 15484 2660 15486
rect 2604 15474 2660 15484
rect 1708 15426 1764 15438
rect 1708 15374 1710 15426
rect 1762 15374 1764 15426
rect 1708 14980 1764 15374
rect 2156 15426 2212 15438
rect 2156 15374 2158 15426
rect 2210 15374 2212 15426
rect 2156 15092 2212 15374
rect 2716 15148 2772 15820
rect 3052 15538 3108 16380
rect 3052 15486 3054 15538
rect 3106 15486 3108 15538
rect 3052 15474 3108 15486
rect 3388 15874 3444 15886
rect 3388 15822 3390 15874
rect 3442 15822 3444 15874
rect 3388 15540 3444 15822
rect 3388 15474 3444 15484
rect 3500 15538 3556 17276
rect 3612 16884 3668 16894
rect 3668 16828 3780 16884
rect 3612 16818 3668 16828
rect 3724 15988 3780 16828
rect 3872 16492 4136 16502
rect 3928 16436 3976 16492
rect 4032 16436 4080 16492
rect 3872 16426 4136 16436
rect 3836 15988 3892 15998
rect 3724 15986 3892 15988
rect 3724 15934 3838 15986
rect 3890 15934 3892 15986
rect 3724 15932 3892 15934
rect 4508 15988 4564 19200
rect 7420 17668 7476 19200
rect 7420 17612 7812 17668
rect 7756 16210 7812 17612
rect 9192 16492 9456 16502
rect 9248 16436 9296 16492
rect 9352 16436 9400 16492
rect 9192 16426 9456 16436
rect 7756 16158 7758 16210
rect 7810 16158 7812 16210
rect 7756 16146 7812 16158
rect 8764 16098 8820 16110
rect 8764 16046 8766 16098
rect 8818 16046 8820 16098
rect 4732 15988 4788 15998
rect 4508 15986 4788 15988
rect 4508 15934 4734 15986
rect 4786 15934 4788 15986
rect 4508 15932 4788 15934
rect 3836 15922 3892 15932
rect 4732 15922 4788 15932
rect 8764 15876 8820 16046
rect 10332 15988 10388 19200
rect 10556 15988 10612 15998
rect 10332 15986 10612 15988
rect 10332 15934 10558 15986
rect 10610 15934 10612 15986
rect 10332 15932 10612 15934
rect 13244 15988 13300 19200
rect 14512 16492 14776 16502
rect 14568 16436 14616 16492
rect 14672 16436 14720 16492
rect 14512 16426 14776 16436
rect 16156 16324 16212 19200
rect 16156 16258 16212 16268
rect 17052 16324 17108 16334
rect 17052 16210 17108 16268
rect 17052 16158 17054 16210
rect 17106 16158 17108 16210
rect 17052 16146 17108 16158
rect 13468 15988 13524 15998
rect 13244 15986 13524 15988
rect 13244 15934 13470 15986
rect 13522 15934 13524 15986
rect 13244 15932 13524 15934
rect 19068 15988 19124 19200
rect 19832 16492 20096 16502
rect 19888 16436 19936 16492
rect 19992 16436 20040 16492
rect 19832 16426 20096 16436
rect 21756 16324 21812 16334
rect 21980 16324 22036 19200
rect 21756 16322 22036 16324
rect 21756 16270 21758 16322
rect 21810 16270 22036 16322
rect 21756 16268 22036 16270
rect 22204 17332 22260 17342
rect 21756 16258 21812 16268
rect 19292 15988 19348 15998
rect 19068 15986 19348 15988
rect 19068 15934 19294 15986
rect 19346 15934 19348 15986
rect 19068 15932 19348 15934
rect 10556 15922 10612 15932
rect 13468 15922 13524 15932
rect 19292 15922 19348 15932
rect 8764 15810 8820 15820
rect 9436 15876 9492 15886
rect 9436 15782 9492 15820
rect 15932 15876 15988 15886
rect 6532 15708 6796 15718
rect 6588 15652 6636 15708
rect 6692 15652 6740 15708
rect 6532 15642 6796 15652
rect 11852 15708 12116 15718
rect 11908 15652 11956 15708
rect 12012 15652 12060 15708
rect 11852 15642 12116 15652
rect 3500 15486 3502 15538
rect 3554 15486 3556 15538
rect 3500 15474 3556 15486
rect 2156 15026 2212 15036
rect 2380 15092 2772 15148
rect 1708 14914 1764 14924
rect 1708 14306 1764 14318
rect 1708 14254 1710 14306
rect 1762 14254 1764 14306
rect 1708 14084 1764 14254
rect 2156 14308 2212 14318
rect 2156 14214 2212 14252
rect 1708 14018 1764 14028
rect 1708 13858 1764 13870
rect 1708 13806 1710 13858
rect 1762 13806 1764 13858
rect 1708 13300 1764 13806
rect 1708 13234 1764 13244
rect 1708 12852 1764 12862
rect 1708 12758 1764 12796
rect 2156 12740 2212 12750
rect 2156 12646 2212 12684
rect 1708 12290 1764 12302
rect 1708 12238 1710 12290
rect 1762 12238 1764 12290
rect 1708 11956 1764 12238
rect 1708 11890 1764 11900
rect 2156 12290 2212 12302
rect 2156 12238 2158 12290
rect 2210 12238 2212 12290
rect 2156 11508 2212 12238
rect 2380 11788 2436 15092
rect 3872 14924 4136 14934
rect 3928 14868 3976 14924
rect 4032 14868 4080 14924
rect 3872 14858 4136 14868
rect 9192 14924 9456 14934
rect 9248 14868 9296 14924
rect 9352 14868 9400 14924
rect 9192 14858 9456 14868
rect 14512 14924 14776 14934
rect 14568 14868 14616 14924
rect 14672 14868 14720 14924
rect 14512 14858 14776 14868
rect 6532 14140 6796 14150
rect 6588 14084 6636 14140
rect 6692 14084 6740 14140
rect 6532 14074 6796 14084
rect 11852 14140 12116 14150
rect 11908 14084 11956 14140
rect 12012 14084 12060 14140
rect 11852 14074 12116 14084
rect 3872 13356 4136 13366
rect 3928 13300 3976 13356
rect 4032 13300 4080 13356
rect 3872 13290 4136 13300
rect 9192 13356 9456 13366
rect 9248 13300 9296 13356
rect 9352 13300 9400 13356
rect 9192 13290 9456 13300
rect 14512 13356 14776 13366
rect 14568 13300 14616 13356
rect 14672 13300 14720 13356
rect 14512 13290 14776 13300
rect 6532 12572 6796 12582
rect 6588 12516 6636 12572
rect 6692 12516 6740 12572
rect 6532 12506 6796 12516
rect 11852 12572 12116 12582
rect 11908 12516 11956 12572
rect 12012 12516 12060 12572
rect 11852 12506 12116 12516
rect 3836 12178 3892 12190
rect 3836 12126 3838 12178
rect 3890 12126 3892 12178
rect 2828 12068 2884 12078
rect 3276 12068 3332 12078
rect 2604 12066 2884 12068
rect 2604 12014 2830 12066
rect 2882 12014 2884 12066
rect 2604 12012 2884 12014
rect 2604 11788 2660 12012
rect 2828 12002 2884 12012
rect 2940 12066 3332 12068
rect 2940 12014 3278 12066
rect 3330 12014 3332 12066
rect 2940 12012 3332 12014
rect 2156 11442 2212 11452
rect 2268 11732 2436 11788
rect 2492 11732 2660 11788
rect 1708 11172 1764 11182
rect 2156 11172 2212 11182
rect 1708 11078 1764 11116
rect 2044 11170 2212 11172
rect 2044 11118 2158 11170
rect 2210 11118 2212 11170
rect 2044 11116 2212 11118
rect 1708 10722 1764 10734
rect 1708 10670 1710 10722
rect 1762 10670 1764 10722
rect 1708 10164 1764 10670
rect 2044 10612 2100 11116
rect 2156 11106 2212 11116
rect 2044 10546 2100 10556
rect 2156 10722 2212 10734
rect 2156 10670 2158 10722
rect 2210 10670 2212 10722
rect 1708 10098 1764 10108
rect 2156 9828 2212 10670
rect 1820 9772 2212 9828
rect 1708 9604 1764 9614
rect 1708 9510 1764 9548
rect 1820 9380 1876 9772
rect 1708 9324 1876 9380
rect 2156 9602 2212 9614
rect 2156 9550 2158 9602
rect 2210 9550 2212 9602
rect 1708 7924 1764 9324
rect 2156 9268 2212 9550
rect 2268 9380 2324 11732
rect 2492 11172 2548 11732
rect 2828 11172 2884 11182
rect 2492 11106 2548 11116
rect 2716 11170 2884 11172
rect 2716 11118 2830 11170
rect 2882 11118 2884 11170
rect 2716 11116 2884 11118
rect 2604 10724 2660 10734
rect 2492 10722 2660 10724
rect 2492 10670 2606 10722
rect 2658 10670 2660 10722
rect 2492 10668 2660 10670
rect 2268 9324 2436 9380
rect 2156 9202 2212 9212
rect 1820 9154 1876 9166
rect 1820 9102 1822 9154
rect 1874 9102 1876 9154
rect 1820 8484 1876 9102
rect 2044 9156 2100 9166
rect 1820 8418 1876 8428
rect 1932 8596 1988 8606
rect 1484 7868 1764 7924
rect 1820 8034 1876 8046
rect 1820 7982 1822 8034
rect 1874 7982 1876 8034
rect 1820 7924 1876 7982
rect 1484 4564 1540 7868
rect 1820 7858 1876 7868
rect 1820 7700 1876 7710
rect 1708 7588 1764 7598
rect 1708 7476 1764 7532
rect 1484 4498 1540 4508
rect 1596 7474 1764 7476
rect 1596 7422 1710 7474
rect 1762 7422 1764 7474
rect 1596 7420 1764 7422
rect 1596 2882 1652 7420
rect 1708 7410 1764 7420
rect 1708 6466 1764 6478
rect 1708 6414 1710 6466
rect 1762 6414 1764 6466
rect 1708 6132 1764 6414
rect 1708 6066 1764 6076
rect 1596 2830 1598 2882
rect 1650 2830 1652 2882
rect 1596 2818 1652 2830
rect 1708 4898 1764 4910
rect 1708 4846 1710 4898
rect 1762 4846 1764 4898
rect 1708 2548 1764 4846
rect 1820 4788 1876 7644
rect 1932 6468 1988 8540
rect 2044 7698 2100 9100
rect 2268 9154 2324 9166
rect 2268 9102 2270 9154
rect 2322 9102 2324 9154
rect 2268 8596 2324 9102
rect 2268 8530 2324 8540
rect 2044 7646 2046 7698
rect 2098 7646 2100 7698
rect 2044 7634 2100 7646
rect 2156 8034 2212 8046
rect 2380 8036 2436 9324
rect 2492 8820 2548 10668
rect 2604 10658 2660 10668
rect 2492 8754 2548 8764
rect 2604 9602 2660 9614
rect 2604 9550 2606 9602
rect 2658 9550 2660 9602
rect 2604 8484 2660 9550
rect 2716 9380 2772 11116
rect 2828 11106 2884 11116
rect 2940 10836 2996 12012
rect 3276 12002 3332 12012
rect 3724 12068 3780 12078
rect 3836 12068 3892 12126
rect 3780 12012 3892 12068
rect 4284 12066 4340 12078
rect 4284 12014 4286 12066
rect 4338 12014 4340 12066
rect 3724 12002 3780 12012
rect 3872 11788 4136 11798
rect 3928 11732 3976 11788
rect 4032 11732 4080 11788
rect 4284 11788 4340 12014
rect 9192 11788 9456 11798
rect 4284 11732 4452 11788
rect 3872 11722 4136 11732
rect 3388 11172 3444 11182
rect 3388 11078 3444 11116
rect 3724 11170 3780 11182
rect 3724 11118 3726 11170
rect 3778 11118 3780 11170
rect 2716 9314 2772 9324
rect 2828 10780 2996 10836
rect 2716 9156 2772 9166
rect 2716 9062 2772 9100
rect 2604 8418 2660 8428
rect 2828 8260 2884 10780
rect 3052 10724 3108 10734
rect 2940 10722 3108 10724
rect 2940 10670 3054 10722
rect 3106 10670 3108 10722
rect 2940 10668 3108 10670
rect 2940 8484 2996 10668
rect 3052 10658 3108 10668
rect 3724 10612 3780 11118
rect 3724 10546 3780 10556
rect 4060 10498 4116 10510
rect 4060 10446 4062 10498
rect 4114 10446 4116 10498
rect 4060 10388 4116 10446
rect 3500 10332 4116 10388
rect 2940 8418 2996 8428
rect 3052 9602 3108 9614
rect 3052 9550 3054 9602
rect 3106 9550 3108 9602
rect 2156 7982 2158 8034
rect 2210 7982 2212 8034
rect 2156 7364 2212 7982
rect 2156 7298 2212 7308
rect 2268 7980 2436 8036
rect 2492 8204 2884 8260
rect 3052 8260 3108 9550
rect 3388 9380 3444 9390
rect 3276 9156 3332 9166
rect 3276 9062 3332 9100
rect 3388 9154 3444 9324
rect 3388 9102 3390 9154
rect 3442 9102 3444 9154
rect 3388 9090 3444 9102
rect 3276 8818 3332 8830
rect 3276 8766 3278 8818
rect 3330 8766 3332 8818
rect 3052 8204 3220 8260
rect 2156 6804 2212 6814
rect 2268 6804 2324 7980
rect 2380 7812 2436 7822
rect 2380 7476 2436 7756
rect 2492 7588 2548 8204
rect 2716 8036 2772 8046
rect 2716 7942 2772 7980
rect 3052 8034 3108 8046
rect 3052 7982 3054 8034
rect 3106 7982 3108 8034
rect 2940 7924 2996 7934
rect 2828 7868 2940 7924
rect 2716 7700 2772 7710
rect 2828 7700 2884 7868
rect 2940 7858 2996 7868
rect 2716 7698 2884 7700
rect 2716 7646 2718 7698
rect 2770 7646 2884 7698
rect 2716 7644 2884 7646
rect 3052 7700 3108 7982
rect 2716 7634 2772 7644
rect 3052 7634 3108 7644
rect 2492 7532 2660 7588
rect 2380 7474 2548 7476
rect 2380 7422 2382 7474
rect 2434 7422 2548 7474
rect 2380 7420 2548 7422
rect 2380 7410 2436 7420
rect 2156 6802 2324 6804
rect 2156 6750 2158 6802
rect 2210 6750 2324 6802
rect 2156 6748 2324 6750
rect 2156 6738 2212 6748
rect 1932 6402 1988 6412
rect 2044 6132 2100 6142
rect 2268 6132 2324 6142
rect 2044 6130 2268 6132
rect 2044 6078 2046 6130
rect 2098 6078 2268 6130
rect 2044 6076 2268 6078
rect 2044 6066 2100 6076
rect 2268 6066 2324 6076
rect 1932 6018 1988 6030
rect 1932 5966 1934 6018
rect 1986 5966 1988 6018
rect 1932 5348 1988 5966
rect 2156 5796 2212 5806
rect 2156 5702 2212 5740
rect 1932 5282 1988 5292
rect 2380 5124 2436 5134
rect 1820 4722 1876 4732
rect 1932 5122 2436 5124
rect 1932 5070 2382 5122
rect 2434 5070 2436 5122
rect 1932 5068 2436 5070
rect 1932 4226 1988 5068
rect 2380 5058 2436 5068
rect 2492 4340 2548 7420
rect 2604 5906 2660 7532
rect 3052 7476 3108 7486
rect 2940 7474 3108 7476
rect 2940 7422 3054 7474
rect 3106 7422 3108 7474
rect 2940 7420 3108 7422
rect 2828 6356 2884 6366
rect 2828 6130 2884 6300
rect 2828 6078 2830 6130
rect 2882 6078 2884 6130
rect 2828 6066 2884 6078
rect 2940 6132 2996 7420
rect 3052 7410 3108 7420
rect 2940 6066 2996 6076
rect 3052 7250 3108 7262
rect 3052 7198 3054 7250
rect 3106 7198 3108 7250
rect 2604 5854 2606 5906
rect 2658 5854 2660 5906
rect 2604 4676 2660 5854
rect 3052 5796 3108 7198
rect 2828 5740 3108 5796
rect 2604 4610 2660 4620
rect 2716 5124 2772 5134
rect 2492 4274 2548 4284
rect 1932 4174 1934 4226
rect 1986 4174 1988 4226
rect 1932 4162 1988 4174
rect 1932 3780 1988 3790
rect 1932 3686 1988 3724
rect 2716 3554 2772 5068
rect 2828 4452 2884 5740
rect 3164 4564 3220 8204
rect 3276 7588 3332 8766
rect 3500 8258 3556 10332
rect 3872 10220 4136 10230
rect 3928 10164 3976 10220
rect 4032 10164 4080 10220
rect 3872 10154 4136 10164
rect 3724 9604 3780 9614
rect 3500 8206 3502 8258
rect 3554 8206 3556 8258
rect 3388 7588 3444 7598
rect 3276 7586 3444 7588
rect 3276 7534 3390 7586
rect 3442 7534 3444 7586
rect 3276 7532 3444 7534
rect 3388 7522 3444 7532
rect 3388 7140 3444 7150
rect 3276 5908 3332 5918
rect 3276 5814 3332 5852
rect 2828 4386 2884 4396
rect 3052 4508 3220 4564
rect 3276 5572 3332 5582
rect 3276 5122 3332 5516
rect 3276 5070 3278 5122
rect 3330 5070 3332 5122
rect 3052 3668 3108 4508
rect 2716 3502 2718 3554
rect 2770 3502 2772 3554
rect 2716 3490 2772 3502
rect 2828 3612 3108 3668
rect 3164 4340 3220 4350
rect 2828 3388 2884 3612
rect 2492 3332 2884 3388
rect 3052 3444 3108 3482
rect 3052 3378 3108 3388
rect 2492 2996 2548 3332
rect 2492 2930 2548 2940
rect 1708 2482 1764 2492
rect 3164 800 3220 4284
rect 3276 2994 3332 5070
rect 3388 3388 3444 7084
rect 3500 6916 3556 8206
rect 3612 9602 3780 9604
rect 3612 9550 3726 9602
rect 3778 9550 3780 9602
rect 3612 9548 3780 9550
rect 3612 8148 3668 9548
rect 3724 9538 3780 9548
rect 4172 9604 4228 9614
rect 4172 9510 4228 9548
rect 4396 9380 4452 11732
rect 9248 11732 9296 11788
rect 9352 11732 9400 11788
rect 9192 11722 9456 11732
rect 14512 11788 14776 11798
rect 14568 11732 14616 11788
rect 14672 11732 14720 11788
rect 14512 11722 14776 11732
rect 4956 11508 5012 11518
rect 4956 11414 5012 11452
rect 4508 11170 4564 11182
rect 4508 11118 4510 11170
rect 4562 11118 4564 11170
rect 4508 10948 4564 11118
rect 9996 11172 10052 11182
rect 9996 11078 10052 11116
rect 15148 11172 15204 11182
rect 6532 11004 6796 11014
rect 6588 10948 6636 11004
rect 6692 10948 6740 11004
rect 6532 10938 6796 10948
rect 11852 11004 12116 11014
rect 11908 10948 11956 11004
rect 12012 10948 12060 11004
rect 11852 10938 12116 10948
rect 4508 10882 4564 10892
rect 10220 10722 10276 10734
rect 10220 10670 10222 10722
rect 10274 10670 10276 10722
rect 9996 10612 10052 10622
rect 9996 10610 10164 10612
rect 9996 10558 9998 10610
rect 10050 10558 10164 10610
rect 9996 10556 10164 10558
rect 9996 10546 10052 10556
rect 4620 10500 4676 10510
rect 4396 9314 4452 9324
rect 4508 10498 4676 10500
rect 4508 10446 4622 10498
rect 4674 10446 4676 10498
rect 4508 10444 4676 10446
rect 3724 8930 3780 8942
rect 3724 8878 3726 8930
rect 3778 8878 3780 8930
rect 3724 8260 3780 8878
rect 3872 8652 4136 8662
rect 3928 8596 3976 8652
rect 4032 8596 4080 8652
rect 3872 8586 4136 8596
rect 4172 8260 4228 8270
rect 4508 8260 4564 10444
rect 4620 10434 4676 10444
rect 5180 10498 5236 10510
rect 5628 10500 5684 10510
rect 5180 10446 5182 10498
rect 5234 10446 5236 10498
rect 4956 9714 5012 9726
rect 4956 9662 4958 9714
rect 5010 9662 5012 9714
rect 3724 8204 3892 8260
rect 3612 8082 3668 8092
rect 3724 8036 3780 8046
rect 3724 7942 3780 7980
rect 3836 7812 3892 8204
rect 4172 8258 4564 8260
rect 4172 8206 4174 8258
rect 4226 8206 4564 8258
rect 4172 8204 4564 8206
rect 4172 8194 4228 8204
rect 3724 7756 3892 7812
rect 4060 8036 4116 8046
rect 4396 8036 4452 8046
rect 3724 7588 3780 7756
rect 4060 7698 4116 7980
rect 4060 7646 4062 7698
rect 4114 7646 4116 7698
rect 4060 7634 4116 7646
rect 4284 8034 4452 8036
rect 4284 7982 4398 8034
rect 4450 7982 4452 8034
rect 4284 7980 4452 7982
rect 3724 7252 3780 7532
rect 3836 7476 3892 7486
rect 3836 7382 3892 7420
rect 3724 7186 3780 7196
rect 3872 7084 4136 7094
rect 3928 7028 3976 7084
rect 4032 7028 4080 7084
rect 3872 7018 4136 7028
rect 4284 7028 4340 7980
rect 4396 7970 4452 7980
rect 4508 7812 4564 8204
rect 4284 6962 4340 6972
rect 4396 7756 4564 7812
rect 4620 9602 4676 9614
rect 4620 9550 4622 9602
rect 4674 9550 4676 9602
rect 4620 7812 4676 9550
rect 4844 9604 4900 9614
rect 4844 9510 4900 9548
rect 4844 9156 4900 9166
rect 4956 9156 5012 9662
rect 4900 9100 5012 9156
rect 4844 8484 4900 9100
rect 4844 8418 4900 8428
rect 4956 8932 5012 8942
rect 4844 8258 4900 8270
rect 4844 8206 4846 8258
rect 4898 8206 4900 8258
rect 4844 8148 4900 8206
rect 4844 8082 4900 8092
rect 4620 7756 4788 7812
rect 3500 6860 3780 6916
rect 3500 6692 3556 6702
rect 3500 6130 3556 6636
rect 3500 6078 3502 6130
rect 3554 6078 3556 6130
rect 3500 6066 3556 6078
rect 3500 4898 3556 4910
rect 3500 4846 3502 4898
rect 3554 4846 3556 4898
rect 3500 4340 3556 4846
rect 3500 4274 3556 4284
rect 3724 3780 3780 6860
rect 4284 6578 4340 6590
rect 4284 6526 4286 6578
rect 4338 6526 4340 6578
rect 4284 6468 4340 6526
rect 4284 6402 4340 6412
rect 4172 6018 4228 6030
rect 4172 5966 4174 6018
rect 4226 5966 4228 6018
rect 3948 5906 4004 5918
rect 3948 5854 3950 5906
rect 4002 5854 4004 5906
rect 3948 5796 4004 5854
rect 4172 5908 4228 5966
rect 4172 5842 4228 5852
rect 3948 5730 4004 5740
rect 4284 5684 4340 5694
rect 3872 5516 4136 5526
rect 3928 5460 3976 5516
rect 4032 5460 4080 5516
rect 3872 5450 4136 5460
rect 3948 5236 4004 5246
rect 3948 5122 4004 5180
rect 3948 5070 3950 5122
rect 4002 5070 4004 5122
rect 3948 4228 4004 5070
rect 4172 4900 4228 4910
rect 4172 4806 4228 4844
rect 4060 4452 4116 4462
rect 4060 4358 4116 4396
rect 3948 4162 4004 4172
rect 4284 4116 4340 5628
rect 4284 4050 4340 4060
rect 3872 3948 4136 3958
rect 3928 3892 3976 3948
rect 4032 3892 4080 3948
rect 3872 3882 4136 3892
rect 3724 3724 4116 3780
rect 3724 3556 3780 3566
rect 3724 3462 3780 3500
rect 3388 3332 3668 3388
rect 3276 2942 3278 2994
rect 3330 2942 3332 2994
rect 3276 2930 3332 2942
rect 3612 800 3668 3332
rect 4060 800 4116 3724
rect 4284 3556 4340 3566
rect 4284 3462 4340 3500
rect 4396 3332 4452 7756
rect 4620 7586 4676 7598
rect 4620 7534 4622 7586
rect 4674 7534 4676 7586
rect 4620 6580 4676 7534
rect 4732 7140 4788 7756
rect 4732 7074 4788 7084
rect 4620 6514 4676 6524
rect 4844 6692 4900 6702
rect 4732 6020 4788 6030
rect 4732 5926 4788 5964
rect 4844 5794 4900 6636
rect 4844 5742 4846 5794
rect 4898 5742 4900 5794
rect 4844 5730 4900 5742
rect 4508 5682 4564 5694
rect 4508 5630 4510 5682
rect 4562 5630 4564 5682
rect 4508 5572 4564 5630
rect 4508 3778 4564 5516
rect 4620 5180 4900 5236
rect 4620 5122 4676 5180
rect 4620 5070 4622 5122
rect 4674 5070 4676 5122
rect 4620 5058 4676 5070
rect 4508 3726 4510 3778
rect 4562 3726 4564 3778
rect 4508 3714 4564 3726
rect 4732 5010 4788 5022
rect 4732 4958 4734 5010
rect 4786 4958 4788 5010
rect 4732 3668 4788 4958
rect 4844 5012 4900 5180
rect 4844 4946 4900 4956
rect 4956 4898 5012 8876
rect 5068 8034 5124 8046
rect 5068 7982 5070 8034
rect 5122 7982 5124 8034
rect 5068 7252 5124 7982
rect 5180 7476 5236 10446
rect 5404 10498 5684 10500
rect 5404 10446 5630 10498
rect 5682 10446 5684 10498
rect 5404 10444 5684 10446
rect 5180 7410 5236 7420
rect 5292 9268 5348 9278
rect 5068 7186 5124 7196
rect 5180 7140 5236 7150
rect 4956 4846 4958 4898
rect 5010 4846 5012 4898
rect 4956 4834 5012 4846
rect 5068 6916 5124 6926
rect 5068 6690 5124 6860
rect 5068 6638 5070 6690
rect 5122 6638 5124 6690
rect 4844 4340 4900 4350
rect 5068 4340 5124 6638
rect 5180 6692 5236 7084
rect 5180 6626 5236 6636
rect 5180 5236 5236 5246
rect 5180 5122 5236 5180
rect 5180 5070 5182 5122
rect 5234 5070 5236 5122
rect 5180 5058 5236 5070
rect 5292 4450 5348 9212
rect 5404 8820 5460 10444
rect 5628 10434 5684 10444
rect 5964 10498 6020 10510
rect 6524 10500 6580 10510
rect 5964 10446 5966 10498
rect 6018 10446 6020 10498
rect 5964 10386 6020 10446
rect 5964 10334 5966 10386
rect 6018 10334 6020 10386
rect 5852 9602 5908 9614
rect 5852 9550 5854 9602
rect 5906 9550 5908 9602
rect 5852 9156 5908 9550
rect 5964 9380 6020 10334
rect 6412 10498 6580 10500
rect 6412 10446 6526 10498
rect 6578 10446 6580 10498
rect 6412 10444 6580 10446
rect 5964 9314 6020 9324
rect 6300 9602 6356 9614
rect 6300 9550 6302 9602
rect 6354 9550 6356 9602
rect 5404 8754 5460 8764
rect 5516 9100 5908 9156
rect 5404 8372 5460 8382
rect 5404 7700 5460 8316
rect 5404 5796 5460 7644
rect 5404 5730 5460 5740
rect 5516 8148 5572 9100
rect 6300 9044 6356 9550
rect 6412 9268 6468 10444
rect 6524 10434 6580 10444
rect 6972 10500 7028 10510
rect 8988 10500 9044 10510
rect 6972 10498 7140 10500
rect 6972 10446 6974 10498
rect 7026 10446 7140 10498
rect 6972 10444 7140 10446
rect 6972 10434 7028 10444
rect 7084 10386 7140 10444
rect 7084 10334 7086 10386
rect 7138 10334 7140 10386
rect 6972 9602 7028 9614
rect 6972 9550 6974 9602
rect 7026 9550 7028 9602
rect 6532 9436 6796 9446
rect 6588 9380 6636 9436
rect 6692 9380 6740 9436
rect 6532 9370 6796 9380
rect 6412 9212 6692 9268
rect 6524 9044 6580 9054
rect 6076 8988 6356 9044
rect 6412 9042 6580 9044
rect 6412 8990 6526 9042
rect 6578 8990 6580 9042
rect 6412 8988 6580 8990
rect 5852 8932 5908 8942
rect 5852 8838 5908 8876
rect 6076 8708 6132 8988
rect 5852 8652 6132 8708
rect 6188 8820 6244 8830
rect 5292 4398 5294 4450
rect 5346 4398 5348 4450
rect 5292 4386 5348 4398
rect 5404 4676 5460 4686
rect 4844 4338 5124 4340
rect 4844 4286 4846 4338
rect 4898 4286 5124 4338
rect 4844 4284 5124 4286
rect 4844 4274 4900 4284
rect 4844 4116 4900 4126
rect 4900 4060 5012 4116
rect 4844 4050 4900 4060
rect 4844 3668 4900 3678
rect 4732 3666 4900 3668
rect 4732 3614 4846 3666
rect 4898 3614 4900 3666
rect 4732 3612 4900 3614
rect 4844 3602 4900 3612
rect 4956 3554 5012 4060
rect 4956 3502 4958 3554
rect 5010 3502 5012 3554
rect 4956 3490 5012 3502
rect 4732 3444 4788 3482
rect 4732 3378 4788 3388
rect 4396 3276 4564 3332
rect 4508 800 4564 3276
rect 4956 2882 5012 2894
rect 4956 2830 4958 2882
rect 5010 2830 5012 2882
rect 4956 800 5012 2830
rect 5404 800 5460 4620
rect 5516 3220 5572 8092
rect 5740 8260 5796 8270
rect 5852 8260 5908 8652
rect 5740 8258 5908 8260
rect 5740 8206 5742 8258
rect 5794 8206 5908 8258
rect 5740 8204 5908 8206
rect 5964 8260 6020 8270
rect 5740 8148 5796 8204
rect 5740 8082 5796 8092
rect 5964 8146 6020 8204
rect 5964 8094 5966 8146
rect 6018 8094 6020 8146
rect 5964 8082 6020 8094
rect 6076 7588 6132 7598
rect 6188 7588 6244 8764
rect 6300 8372 6356 8382
rect 6300 8146 6356 8316
rect 6300 8094 6302 8146
rect 6354 8094 6356 8146
rect 6300 7812 6356 8094
rect 6300 7746 6356 7756
rect 6412 7700 6468 8988
rect 6524 8978 6580 8988
rect 6636 8596 6692 9212
rect 6860 9042 6916 9054
rect 6860 8990 6862 9042
rect 6914 8990 6916 9042
rect 6860 8820 6916 8990
rect 6860 8754 6916 8764
rect 6636 8530 6692 8540
rect 6972 8372 7028 9550
rect 7084 9604 7140 10334
rect 8876 10498 9044 10500
rect 8876 10446 8990 10498
rect 9042 10446 9044 10498
rect 8876 10444 9044 10446
rect 8652 9716 8708 9726
rect 8876 9716 8932 10444
rect 8988 10434 9044 10444
rect 9192 10220 9456 10230
rect 9248 10164 9296 10220
rect 9352 10164 9400 10220
rect 9192 10154 9456 10164
rect 8540 9714 8932 9716
rect 8540 9662 8654 9714
rect 8706 9662 8932 9714
rect 8540 9660 8932 9662
rect 9772 9826 9828 9838
rect 9772 9774 9774 9826
rect 9826 9774 9828 9826
rect 7420 9604 7476 9614
rect 7084 9548 7420 9604
rect 7420 9510 7476 9548
rect 7868 9602 7924 9614
rect 7868 9550 7870 9602
rect 7922 9550 7924 9602
rect 7084 9156 7140 9166
rect 7084 9062 7140 9100
rect 7196 9044 7252 9054
rect 7756 9044 7812 9054
rect 7868 9044 7924 9550
rect 8428 9604 8484 9614
rect 8428 9510 8484 9548
rect 8092 9156 8148 9166
rect 8092 9154 8372 9156
rect 8092 9102 8094 9154
rect 8146 9102 8372 9154
rect 8092 9100 8372 9102
rect 8092 9090 8148 9100
rect 7196 9042 7364 9044
rect 7196 8990 7198 9042
rect 7250 8990 7364 9042
rect 7196 8988 7364 8990
rect 7196 8978 7252 8988
rect 6972 8306 7028 8316
rect 7084 8932 7140 8942
rect 7084 8370 7140 8876
rect 7084 8318 7086 8370
rect 7138 8318 7140 8370
rect 7084 8306 7140 8318
rect 6636 8148 6692 8158
rect 6636 8054 6692 8092
rect 6972 8034 7028 8046
rect 7196 8036 7252 8046
rect 6972 7982 6974 8034
rect 7026 7982 7028 8034
rect 6532 7868 6796 7878
rect 6588 7812 6636 7868
rect 6692 7812 6740 7868
rect 6532 7802 6796 7812
rect 6412 7644 6580 7700
rect 6300 7588 6356 7598
rect 6188 7586 6356 7588
rect 6188 7534 6302 7586
rect 6354 7534 6356 7586
rect 6188 7532 6356 7534
rect 6076 7140 6132 7532
rect 6300 7522 6356 7532
rect 6076 7084 6468 7140
rect 6076 6916 6132 6926
rect 5964 6692 6020 6702
rect 6076 6692 6132 6860
rect 5964 6690 6132 6692
rect 5964 6638 5966 6690
rect 6018 6638 6132 6690
rect 5964 6636 6132 6638
rect 6188 6804 6244 6814
rect 5964 6626 6020 6636
rect 5628 6578 5684 6590
rect 5628 6526 5630 6578
rect 5682 6526 5684 6578
rect 5628 6468 5684 6526
rect 6188 6578 6244 6748
rect 6412 6690 6468 7084
rect 6412 6638 6414 6690
rect 6466 6638 6468 6690
rect 6412 6626 6468 6638
rect 6188 6526 6190 6578
rect 6242 6526 6244 6578
rect 6188 6514 6244 6526
rect 6524 6580 6580 7644
rect 6860 7588 6916 7598
rect 6748 7476 6804 7486
rect 6636 7474 6804 7476
rect 6636 7422 6750 7474
rect 6802 7422 6804 7474
rect 6636 7420 6804 7422
rect 6636 6804 6692 7420
rect 6748 7410 6804 7420
rect 6860 6916 6916 7532
rect 6972 7140 7028 7982
rect 6972 7074 7028 7084
rect 7084 8034 7252 8036
rect 7084 7982 7198 8034
rect 7250 7982 7252 8034
rect 7084 7980 7252 7982
rect 6860 6850 6916 6860
rect 6636 6738 6692 6748
rect 6748 6692 6804 6702
rect 6748 6598 6804 6636
rect 6524 6514 6580 6524
rect 5628 6402 5684 6412
rect 5740 6466 5796 6478
rect 5740 6414 5742 6466
rect 5794 6414 5796 6466
rect 5740 6356 5796 6414
rect 6300 6468 6356 6478
rect 6300 6466 6468 6468
rect 6300 6414 6302 6466
rect 6354 6414 6468 6466
rect 6300 6412 6468 6414
rect 6300 6402 6356 6412
rect 6076 6356 6132 6366
rect 5740 6300 6020 6356
rect 5852 6132 5908 6142
rect 5628 6020 5684 6030
rect 5628 3556 5684 5964
rect 5628 3462 5684 3500
rect 5740 5796 5796 5806
rect 5740 3442 5796 5740
rect 5852 5234 5908 6076
rect 5852 5182 5854 5234
rect 5906 5182 5908 5234
rect 5852 5124 5908 5182
rect 5852 5058 5908 5068
rect 5964 3780 6020 6300
rect 6132 6300 6244 6356
rect 6076 6290 6132 6300
rect 6188 6020 6244 6300
rect 6300 6020 6356 6030
rect 6188 6018 6356 6020
rect 6188 5966 6302 6018
rect 6354 5966 6356 6018
rect 6188 5964 6356 5966
rect 6412 6020 6468 6412
rect 6532 6300 6796 6310
rect 6588 6244 6636 6300
rect 6692 6244 6740 6300
rect 6532 6234 6796 6244
rect 7084 6132 7140 7980
rect 7196 7970 7252 7980
rect 7308 7700 7364 8988
rect 7644 9042 7924 9044
rect 7644 8990 7758 9042
rect 7810 8990 7924 9042
rect 7644 8988 7924 8990
rect 7420 8034 7476 8046
rect 7420 7982 7422 8034
rect 7474 7982 7476 8034
rect 7420 7924 7476 7982
rect 7420 7858 7476 7868
rect 7308 7644 7476 7700
rect 7084 6066 7140 6076
rect 7196 7028 7252 7038
rect 6412 5964 6580 6020
rect 6188 5572 6244 5582
rect 5964 3714 6020 3724
rect 6076 4452 6132 4462
rect 5740 3390 5742 3442
rect 5794 3390 5796 3442
rect 5740 3378 5796 3390
rect 6076 3220 6132 4396
rect 6188 3442 6244 5516
rect 6300 3668 6356 5964
rect 6300 3602 6356 3612
rect 6412 5796 6468 5806
rect 6412 3556 6468 5740
rect 6524 5124 6580 5964
rect 6524 5058 6580 5068
rect 6860 5908 6916 5918
rect 7196 5908 7252 6972
rect 7308 6580 7364 6590
rect 7308 6486 7364 6524
rect 7420 6468 7476 7644
rect 6860 5124 6916 5852
rect 6860 5058 6916 5068
rect 7084 5906 7252 5908
rect 7084 5854 7198 5906
rect 7250 5854 7252 5906
rect 7084 5852 7252 5854
rect 6860 4900 6916 4910
rect 6532 4732 6796 4742
rect 6588 4676 6636 4732
rect 6692 4676 6740 4732
rect 6532 4666 6796 4676
rect 6412 3490 6468 3500
rect 6188 3390 6190 3442
rect 6242 3390 6244 3442
rect 6188 3378 6244 3390
rect 6412 3332 6468 3342
rect 6412 3238 6468 3276
rect 5516 3164 5908 3220
rect 6076 3164 6356 3220
rect 5852 800 5908 3164
rect 6300 800 6356 3164
rect 6532 3164 6796 3174
rect 6588 3108 6636 3164
rect 6692 3108 6740 3164
rect 6532 3098 6796 3108
rect 6860 2996 6916 4844
rect 6972 4788 7028 4798
rect 6972 4338 7028 4732
rect 7084 4564 7140 5852
rect 7196 5842 7252 5852
rect 7308 6132 7364 6142
rect 7084 4498 7140 4508
rect 6972 4286 6974 4338
rect 7026 4286 7028 4338
rect 6972 4274 7028 4286
rect 7308 4338 7364 6076
rect 7308 4286 7310 4338
rect 7362 4286 7364 4338
rect 7308 4274 7364 4286
rect 7196 4228 7252 4238
rect 6972 3780 7028 3790
rect 6972 3686 7028 3724
rect 7084 3668 7140 3678
rect 7084 3574 7140 3612
rect 6748 2940 6916 2996
rect 6748 800 6804 2940
rect 7196 800 7252 4172
rect 7420 3554 7476 6412
rect 7420 3502 7422 3554
rect 7474 3502 7476 3554
rect 7420 3490 7476 3502
rect 7644 800 7700 8988
rect 7756 8978 7812 8988
rect 8204 8708 8260 8718
rect 8092 8652 8204 8708
rect 7868 8258 7924 8270
rect 7868 8206 7870 8258
rect 7922 8206 7924 8258
rect 7868 8036 7924 8206
rect 7980 8148 8036 8158
rect 7980 8054 8036 8092
rect 7868 7970 7924 7980
rect 7756 7364 7812 7374
rect 7756 6020 7812 7308
rect 7980 7362 8036 7374
rect 7980 7310 7982 7362
rect 8034 7310 8036 7362
rect 7980 6244 8036 7310
rect 7756 6018 7924 6020
rect 7756 5966 7758 6018
rect 7810 5966 7924 6018
rect 7756 5964 7924 5966
rect 7756 5954 7812 5964
rect 7756 5124 7812 5134
rect 7756 3666 7812 5068
rect 7868 5012 7924 5964
rect 7980 5796 8036 6188
rect 7980 5730 8036 5740
rect 7980 5236 8036 5246
rect 8092 5236 8148 8652
rect 8204 8642 8260 8652
rect 8316 8148 8372 9100
rect 8428 9042 8484 9054
rect 8428 8990 8430 9042
rect 8482 8990 8484 9042
rect 8428 8932 8484 8990
rect 8428 8866 8484 8876
rect 8316 8082 8372 8092
rect 7980 5234 8148 5236
rect 7980 5182 7982 5234
rect 8034 5182 8148 5234
rect 7980 5180 8148 5182
rect 8204 7700 8260 7710
rect 7980 5170 8036 5180
rect 7868 4956 8148 5012
rect 7980 4676 8036 4686
rect 7756 3614 7758 3666
rect 7810 3614 7812 3666
rect 7756 3602 7812 3614
rect 7868 4564 7924 4574
rect 7868 3554 7924 4508
rect 7868 3502 7870 3554
rect 7922 3502 7924 3554
rect 7868 3490 7924 3502
rect 7980 3444 8036 4620
rect 8092 3554 8148 4956
rect 8092 3502 8094 3554
rect 8146 3502 8148 3554
rect 8092 3490 8148 3502
rect 8204 3388 8260 7644
rect 8316 7586 8372 7598
rect 8316 7534 8318 7586
rect 8370 7534 8372 7586
rect 8316 7476 8372 7534
rect 8316 7410 8372 7420
rect 8428 7364 8484 7374
rect 7980 3378 8036 3388
rect 8092 3332 8260 3388
rect 8316 5794 8372 5806
rect 8316 5742 8318 5794
rect 8370 5742 8372 5794
rect 8316 3444 8372 5742
rect 8428 4788 8484 7308
rect 8540 4900 8596 9660
rect 8652 9650 8708 9660
rect 8988 9604 9044 9614
rect 9772 9604 9828 9774
rect 10108 9828 10164 10556
rect 10220 10388 10276 10670
rect 11116 10612 11172 10622
rect 10892 10610 11172 10612
rect 10892 10558 11118 10610
rect 11170 10558 11172 10610
rect 10892 10556 11172 10558
rect 10668 10498 10724 10510
rect 10668 10446 10670 10498
rect 10722 10446 10724 10498
rect 10444 10388 10500 10398
rect 10220 10386 10500 10388
rect 10220 10334 10446 10386
rect 10498 10334 10500 10386
rect 10220 10332 10500 10334
rect 10444 10322 10500 10332
rect 10668 9828 10724 10446
rect 10108 9772 10724 9828
rect 10780 9828 10836 9838
rect 10892 9828 10948 10556
rect 11116 10546 11172 10556
rect 11676 10498 11732 10510
rect 11676 10446 11678 10498
rect 11730 10446 11732 10498
rect 10780 9826 10948 9828
rect 10780 9774 10782 9826
rect 10834 9774 10948 9826
rect 10780 9772 10948 9774
rect 11004 10386 11060 10398
rect 11004 10334 11006 10386
rect 11058 10334 11060 10386
rect 8988 9602 9156 9604
rect 8988 9550 8990 9602
rect 9042 9550 9156 9602
rect 8988 9548 9156 9550
rect 8988 9538 9044 9548
rect 8764 9042 8820 9054
rect 8764 8990 8766 9042
rect 8818 8990 8820 9042
rect 8652 6916 8708 6926
rect 8652 5122 8708 6860
rect 8764 6132 8820 8990
rect 8988 9042 9044 9054
rect 8988 8990 8990 9042
rect 9042 8990 9044 9042
rect 8876 8930 8932 8942
rect 8876 8878 8878 8930
rect 8930 8878 8932 8930
rect 8876 8708 8932 8878
rect 8876 8642 8932 8652
rect 8876 7474 8932 7486
rect 8876 7422 8878 7474
rect 8930 7422 8932 7474
rect 8876 7364 8932 7422
rect 8876 7298 8932 7308
rect 8988 6580 9044 8990
rect 9100 9044 9156 9548
rect 9212 9044 9268 9054
rect 9100 8988 9212 9044
rect 9212 8978 9268 8988
rect 9192 8652 9456 8662
rect 9248 8596 9296 8652
rect 9352 8596 9400 8652
rect 9192 8586 9456 8596
rect 9548 7588 9604 7598
rect 9548 7494 9604 7532
rect 9192 7084 9456 7094
rect 9248 7028 9296 7084
rect 9352 7028 9400 7084
rect 9192 7018 9456 7028
rect 8988 6524 9716 6580
rect 9548 6132 9604 6142
rect 8764 6130 9604 6132
rect 8764 6078 9550 6130
rect 9602 6078 9604 6130
rect 8764 6076 9604 6078
rect 9548 6066 9604 6076
rect 9548 5908 9604 5918
rect 9548 5814 9604 5852
rect 9660 5684 9716 6524
rect 9548 5628 9716 5684
rect 9192 5516 9456 5526
rect 9248 5460 9296 5516
rect 9352 5460 9400 5516
rect 9192 5450 9456 5460
rect 9548 5348 9604 5628
rect 9772 5460 9828 9548
rect 9996 9602 10052 9614
rect 9996 9550 9998 9602
rect 10050 9550 10052 9602
rect 9996 9156 10052 9550
rect 9996 9090 10052 9100
rect 10108 9154 10164 9166
rect 10108 9102 10110 9154
rect 10162 9102 10164 9154
rect 10108 8820 10164 9102
rect 10108 8754 10164 8764
rect 9884 8260 9940 8270
rect 9884 8166 9940 8204
rect 9996 8034 10052 8046
rect 9996 7982 9998 8034
rect 10050 7982 10052 8034
rect 9884 5684 9940 5694
rect 9884 5590 9940 5628
rect 9772 5404 9940 5460
rect 8652 5070 8654 5122
rect 8706 5070 8708 5122
rect 8652 5058 8708 5070
rect 9436 5292 9604 5348
rect 9660 5348 9716 5358
rect 9716 5292 9828 5348
rect 8988 5012 9044 5022
rect 8540 4844 8820 4900
rect 8428 4732 8596 4788
rect 8316 3378 8372 3388
rect 8092 800 8148 3332
rect 8540 800 8596 4732
rect 8652 3668 8708 3678
rect 8652 2994 8708 3612
rect 8764 3388 8820 4844
rect 8876 4562 8932 4574
rect 8876 4510 8878 4562
rect 8930 4510 8932 4562
rect 8876 4452 8932 4510
rect 8876 4386 8932 4396
rect 8988 4450 9044 4956
rect 9436 4562 9492 5292
rect 9660 5282 9716 5292
rect 9660 5012 9716 5022
rect 9436 4510 9438 4562
rect 9490 4510 9492 4562
rect 9436 4498 9492 4510
rect 9548 5010 9716 5012
rect 9548 4958 9662 5010
rect 9714 4958 9716 5010
rect 9548 4956 9716 4958
rect 8988 4398 8990 4450
rect 9042 4398 9044 4450
rect 8988 4386 9044 4398
rect 9192 3948 9456 3958
rect 9248 3892 9296 3948
rect 9352 3892 9400 3948
rect 9192 3882 9456 3892
rect 9548 3780 9604 4956
rect 9660 4946 9716 4956
rect 9660 4564 9716 4574
rect 9660 4470 9716 4508
rect 9772 4450 9828 5292
rect 9772 4398 9774 4450
rect 9826 4398 9828 4450
rect 9772 4386 9828 4398
rect 9884 4116 9940 5404
rect 9212 3724 9604 3780
rect 9772 4060 9940 4116
rect 9996 4228 10052 7982
rect 10332 7924 10388 9772
rect 10556 9602 10612 9614
rect 10556 9550 10558 9602
rect 10610 9550 10612 9602
rect 10444 8148 10500 8158
rect 10444 8054 10500 8092
rect 10332 7868 10500 7924
rect 10220 7588 10276 7598
rect 10108 6468 10164 6478
rect 10108 6018 10164 6412
rect 10108 5966 10110 6018
rect 10162 5966 10164 6018
rect 10108 5954 10164 5966
rect 9212 3388 9268 3724
rect 9772 3388 9828 4060
rect 9996 3554 10052 4172
rect 10220 4226 10276 7532
rect 10332 6244 10388 6254
rect 10332 6018 10388 6188
rect 10332 5966 10334 6018
rect 10386 5966 10388 6018
rect 10332 5954 10388 5966
rect 10220 4174 10222 4226
rect 10274 4174 10276 4226
rect 10220 4162 10276 4174
rect 9996 3502 9998 3554
rect 10050 3502 10052 3554
rect 9996 3490 10052 3502
rect 8764 3332 9044 3388
rect 9212 3332 9380 3388
rect 8652 2942 8654 2994
rect 8706 2942 8708 2994
rect 8652 2930 8708 2942
rect 8988 800 9044 3332
rect 9324 3266 9380 3276
rect 9436 3332 9828 3388
rect 9884 3444 9940 3482
rect 10108 3444 10164 3454
rect 9884 3378 9940 3388
rect 9996 3332 10164 3388
rect 10444 3388 10500 7868
rect 10556 4900 10612 9550
rect 10668 6692 10724 6702
rect 10668 5684 10724 6636
rect 10668 5618 10724 5628
rect 10556 4834 10612 4844
rect 10668 5122 10724 5134
rect 10668 5070 10670 5122
rect 10722 5070 10724 5122
rect 10668 4676 10724 5070
rect 10556 4620 10724 4676
rect 10556 3666 10612 4620
rect 10668 4450 10724 4462
rect 10668 4398 10670 4450
rect 10722 4398 10724 4450
rect 10668 4228 10724 4398
rect 10668 4162 10724 4172
rect 10556 3614 10558 3666
rect 10610 3614 10612 3666
rect 10556 3602 10612 3614
rect 10444 3332 10612 3388
rect 9436 800 9492 3332
rect 9996 2212 10052 3332
rect 9884 2156 10052 2212
rect 10332 3276 10612 3332
rect 9884 800 9940 2156
rect 10332 800 10388 3276
rect 10780 800 10836 9772
rect 11004 9044 11060 10334
rect 11452 9826 11508 9838
rect 11452 9774 11454 9826
rect 11506 9774 11508 9826
rect 11228 9602 11284 9614
rect 11228 9550 11230 9602
rect 11282 9550 11284 9602
rect 11228 9268 11284 9550
rect 11228 9202 11284 9212
rect 11452 9604 11508 9774
rect 11116 9044 11172 9054
rect 11004 9042 11172 9044
rect 11004 8990 11118 9042
rect 11170 8990 11172 9042
rect 11004 8988 11172 8990
rect 11116 8978 11172 8988
rect 11340 8930 11396 8942
rect 11340 8878 11342 8930
rect 11394 8878 11396 8930
rect 11116 7698 11172 7710
rect 11116 7646 11118 7698
rect 11170 7646 11172 7698
rect 11116 5348 11172 7646
rect 11228 7476 11284 7486
rect 11228 6804 11284 7420
rect 11228 6738 11284 6748
rect 11116 4900 11172 5292
rect 11116 4834 11172 4844
rect 10892 4452 10948 4462
rect 10892 3442 10948 4396
rect 11340 4340 11396 8878
rect 11004 4338 11396 4340
rect 11004 4286 11342 4338
rect 11394 4286 11396 4338
rect 11004 4284 11396 4286
rect 11004 3554 11060 4284
rect 11340 4274 11396 4284
rect 11004 3502 11006 3554
rect 11058 3502 11060 3554
rect 11004 3490 11060 3502
rect 10892 3390 10894 3442
rect 10946 3390 10948 3442
rect 10892 3378 10948 3390
rect 11452 3388 11508 9548
rect 11676 9828 11732 10446
rect 12124 10500 12180 10510
rect 12124 10406 12180 10444
rect 14512 10220 14776 10230
rect 14568 10164 14616 10220
rect 14672 10164 14720 10220
rect 14512 10154 14776 10164
rect 12236 9828 12292 9838
rect 11676 9826 12292 9828
rect 11676 9774 12238 9826
rect 12290 9774 12292 9826
rect 11676 9772 12292 9774
rect 11564 9044 11620 9054
rect 11564 8950 11620 8988
rect 11228 3332 11508 3388
rect 11228 800 11284 3332
rect 11676 800 11732 9772
rect 12236 9762 12292 9772
rect 11900 9604 11956 9614
rect 12684 9604 12740 9614
rect 11900 9602 12292 9604
rect 11900 9550 11902 9602
rect 11954 9550 12292 9602
rect 11900 9548 12292 9550
rect 11900 9538 11956 9548
rect 11852 9436 12116 9446
rect 11908 9380 11956 9436
rect 12012 9380 12060 9436
rect 11852 9370 12116 9380
rect 12124 9156 12180 9166
rect 12124 9062 12180 9100
rect 12236 8260 12292 9548
rect 12684 9510 12740 9548
rect 15148 9266 15204 11116
rect 15148 9214 15150 9266
rect 15202 9214 15204 9266
rect 13692 9044 13748 9054
rect 13580 9042 13748 9044
rect 13580 8990 13694 9042
rect 13746 8990 13748 9042
rect 13580 8988 13748 8990
rect 12908 8932 12964 8942
rect 12236 8194 12292 8204
rect 12460 8260 12516 8270
rect 12572 8260 12628 8270
rect 12516 8258 12628 8260
rect 12516 8206 12574 8258
rect 12626 8206 12628 8258
rect 12516 8204 12628 8206
rect 12348 8036 12404 8046
rect 12236 8034 12404 8036
rect 12236 7982 12350 8034
rect 12402 7982 12404 8034
rect 12236 7980 12404 7982
rect 11852 7868 12116 7878
rect 11908 7812 11956 7868
rect 12012 7812 12060 7868
rect 11852 7802 12116 7812
rect 12124 7588 12180 7598
rect 12124 7494 12180 7532
rect 11852 6300 12116 6310
rect 11908 6244 11956 6300
rect 12012 6244 12060 6300
rect 11852 6234 12116 6244
rect 12236 6132 12292 7980
rect 12348 7970 12404 7980
rect 12348 6692 12404 6702
rect 12348 6598 12404 6636
rect 12236 6066 12292 6076
rect 11852 4732 12116 4742
rect 11908 4676 11956 4732
rect 12012 4676 12060 4732
rect 11852 4666 12116 4676
rect 11788 4452 11844 4462
rect 11788 4338 11844 4396
rect 11788 4286 11790 4338
rect 11842 4286 11844 4338
rect 11788 4274 11844 4286
rect 11852 3164 12116 3174
rect 11908 3108 11956 3164
rect 12012 3108 12060 3164
rect 11852 3098 12116 3108
rect 12460 2996 12516 8204
rect 12572 8194 12628 8204
rect 12796 6690 12852 6702
rect 12796 6638 12798 6690
rect 12850 6638 12852 6690
rect 12684 6578 12740 6590
rect 12684 6526 12686 6578
rect 12738 6526 12740 6578
rect 12684 6356 12740 6526
rect 12796 6580 12852 6638
rect 12796 6514 12852 6524
rect 12908 6356 12964 8876
rect 13468 8258 13524 8270
rect 13468 8206 13470 8258
rect 13522 8206 13524 8258
rect 12684 6300 12964 6356
rect 13020 7476 13076 7486
rect 13020 6020 13076 7420
rect 12796 5964 13076 6020
rect 13356 7474 13412 7486
rect 13356 7422 13358 7474
rect 13410 7422 13412 7474
rect 13356 7364 13412 7422
rect 12796 5124 12852 5964
rect 12684 5122 12852 5124
rect 12684 5070 12798 5122
rect 12850 5070 12852 5122
rect 12684 5068 12852 5070
rect 12124 2940 12516 2996
rect 12572 3668 12628 3678
rect 12124 800 12180 2940
rect 12572 800 12628 3612
rect 12684 3556 12740 5068
rect 12796 5058 12852 5068
rect 13244 5236 13300 5246
rect 12908 5012 12964 5022
rect 12908 4918 12964 4956
rect 12796 4900 12852 4910
rect 12796 4806 12852 4844
rect 13132 4788 13188 4798
rect 13020 4340 13076 4350
rect 13020 4246 13076 4284
rect 12684 3490 12740 3500
rect 13132 3554 13188 4732
rect 13244 3778 13300 5180
rect 13356 5012 13412 7308
rect 13468 6916 13524 8206
rect 13468 6850 13524 6860
rect 13468 6692 13524 6702
rect 13468 6018 13524 6636
rect 13468 5966 13470 6018
rect 13522 5966 13524 6018
rect 13468 5954 13524 5966
rect 13356 4946 13412 4956
rect 13468 5796 13524 5806
rect 13468 4900 13524 5740
rect 13580 5234 13636 8988
rect 13692 8978 13748 8988
rect 14028 9042 14084 9054
rect 14028 8990 14030 9042
rect 14082 8990 14084 9042
rect 13692 7476 13748 7486
rect 13692 7362 13748 7420
rect 13692 7310 13694 7362
rect 13746 7310 13748 7362
rect 13692 7298 13748 7310
rect 14028 6804 14084 8990
rect 14364 9042 14420 9054
rect 14364 8990 14366 9042
rect 14418 8990 14420 9042
rect 14140 8930 14196 8942
rect 14140 8878 14142 8930
rect 14194 8878 14196 8930
rect 14140 8372 14196 8878
rect 14252 8372 14308 8382
rect 14140 8370 14308 8372
rect 14140 8318 14254 8370
rect 14306 8318 14308 8370
rect 14140 8316 14308 8318
rect 14252 8306 14308 8316
rect 14028 6738 14084 6748
rect 14140 7252 14196 7262
rect 13580 5182 13582 5234
rect 13634 5182 13636 5234
rect 13580 5170 13636 5182
rect 14028 6020 14084 6030
rect 14028 5684 14084 5964
rect 14028 5122 14084 5628
rect 14028 5070 14030 5122
rect 14082 5070 14084 5122
rect 14028 5058 14084 5070
rect 13804 5012 13860 5022
rect 13468 4806 13524 4844
rect 13692 4900 13748 4910
rect 13692 4564 13748 4844
rect 13692 4498 13748 4508
rect 13244 3726 13246 3778
rect 13298 3726 13300 3778
rect 13244 3714 13300 3726
rect 13804 3778 13860 4956
rect 14140 5012 14196 7196
rect 14252 6132 14308 6142
rect 14364 6132 14420 8990
rect 14700 8932 14756 8942
rect 14700 8930 14980 8932
rect 14700 8878 14702 8930
rect 14754 8878 14980 8930
rect 14700 8876 14980 8878
rect 14700 8866 14756 8876
rect 14512 8652 14776 8662
rect 14568 8596 14616 8652
rect 14672 8596 14720 8652
rect 14512 8586 14776 8596
rect 14512 7084 14776 7094
rect 14568 7028 14616 7084
rect 14672 7028 14720 7084
rect 14512 7018 14776 7028
rect 14308 6076 14420 6132
rect 14252 6066 14308 6076
rect 14924 6020 14980 8876
rect 14924 5954 14980 5964
rect 14512 5516 14776 5526
rect 14568 5460 14616 5516
rect 14672 5460 14720 5516
rect 14512 5450 14776 5460
rect 14140 4946 14196 4956
rect 15036 5348 15092 5358
rect 14812 4900 14868 4910
rect 14812 4898 14980 4900
rect 14812 4846 14814 4898
rect 14866 4846 14980 4898
rect 14812 4844 14980 4846
rect 14812 4834 14868 4844
rect 14252 4452 14308 4462
rect 14252 4358 14308 4396
rect 14364 4340 14420 4350
rect 14140 4226 14196 4238
rect 14140 4174 14142 4226
rect 14194 4174 14196 4226
rect 13804 3726 13806 3778
rect 13858 3726 13860 3778
rect 13804 3714 13860 3726
rect 13916 4116 13972 4126
rect 13132 3502 13134 3554
rect 13186 3502 13188 3554
rect 13132 3490 13188 3502
rect 13580 3668 13636 3678
rect 13020 3444 13076 3454
rect 13020 800 13076 3388
rect 13244 3332 13300 3342
rect 13244 3238 13300 3276
rect 13580 1876 13636 3612
rect 13468 1820 13636 1876
rect 13468 800 13524 1820
rect 13916 800 13972 4060
rect 14140 3442 14196 4174
rect 14140 3390 14142 3442
rect 14194 3390 14196 3442
rect 14140 3378 14196 3390
rect 14364 800 14420 4284
rect 14512 3948 14776 3958
rect 14568 3892 14616 3948
rect 14672 3892 14720 3948
rect 14512 3882 14776 3892
rect 14924 3554 14980 4844
rect 14924 3502 14926 3554
rect 14978 3502 14980 3554
rect 14924 3490 14980 3502
rect 15036 3332 15092 5292
rect 15148 4900 15204 9214
rect 15484 9604 15540 9614
rect 15148 4834 15204 4844
rect 15260 5908 15316 5918
rect 15148 4338 15204 4350
rect 15148 4286 15150 4338
rect 15202 4286 15204 4338
rect 15148 3780 15204 4286
rect 15148 3714 15204 3724
rect 14812 3276 15092 3332
rect 14812 800 14868 3276
rect 15260 800 15316 5852
rect 15484 4676 15540 9548
rect 15820 7364 15876 7374
rect 15820 7270 15876 7308
rect 15596 6804 15652 6814
rect 15652 6748 15764 6804
rect 15596 6738 15652 6748
rect 15708 4788 15764 6748
rect 15932 6580 15988 15820
rect 17724 15874 17780 15886
rect 17724 15822 17726 15874
rect 17778 15822 17780 15874
rect 17172 15708 17436 15718
rect 17228 15652 17276 15708
rect 17332 15652 17380 15708
rect 17172 15642 17436 15652
rect 17172 14140 17436 14150
rect 17228 14084 17276 14140
rect 17332 14084 17380 14140
rect 17172 14074 17436 14084
rect 17172 12572 17436 12582
rect 17228 12516 17276 12572
rect 17332 12516 17380 12572
rect 17172 12506 17436 12516
rect 17724 11788 17780 15822
rect 20300 15876 20356 15886
rect 20972 15876 21028 15886
rect 20300 15874 21028 15876
rect 20300 15822 20302 15874
rect 20354 15822 20974 15874
rect 21026 15822 21028 15874
rect 20300 15820 21028 15822
rect 19832 14924 20096 14934
rect 19888 14868 19936 14924
rect 19992 14868 20040 14924
rect 19832 14858 20096 14868
rect 19832 13356 20096 13366
rect 19888 13300 19936 13356
rect 19992 13300 20040 13356
rect 19832 13290 20096 13300
rect 19832 11788 20096 11798
rect 17724 11732 18004 11788
rect 16380 11172 16436 11182
rect 16380 8370 16436 11116
rect 17172 11004 17436 11014
rect 17228 10948 17276 11004
rect 17332 10948 17380 11004
rect 17172 10938 17436 10948
rect 17172 9436 17436 9446
rect 17228 9380 17276 9436
rect 17332 9380 17380 9436
rect 17172 9370 17436 9380
rect 16380 8318 16382 8370
rect 16434 8318 16436 8370
rect 16380 8306 16436 8318
rect 16828 8034 16884 8046
rect 17388 8036 17444 8046
rect 16828 7982 16830 8034
rect 16882 7982 16884 8034
rect 16492 7474 16548 7486
rect 16492 7422 16494 7474
rect 16546 7422 16548 7474
rect 16492 6916 16548 7422
rect 16492 6802 16548 6860
rect 16492 6750 16494 6802
rect 16546 6750 16548 6802
rect 16492 6738 16548 6750
rect 16716 7252 16772 7262
rect 15932 6514 15988 6524
rect 16716 6468 16772 7196
rect 16716 6402 16772 6412
rect 16828 6244 16884 7982
rect 17052 8034 17444 8036
rect 17052 7982 17390 8034
rect 17442 7982 17444 8034
rect 17052 7980 17444 7982
rect 16716 6188 16884 6244
rect 16940 6804 16996 6814
rect 16492 6132 16548 6142
rect 15820 6130 16548 6132
rect 15820 6078 16494 6130
rect 16546 6078 16548 6130
rect 15820 6076 16548 6078
rect 15820 5010 15876 6076
rect 16492 6066 16548 6076
rect 16156 5906 16212 5918
rect 16156 5854 16158 5906
rect 16210 5854 16212 5906
rect 16156 5124 16212 5854
rect 16716 5906 16772 6188
rect 16716 5854 16718 5906
rect 16770 5854 16772 5906
rect 16492 5572 16548 5582
rect 16156 5058 16212 5068
rect 16380 5236 16436 5246
rect 16380 5122 16436 5180
rect 16380 5070 16382 5122
rect 16434 5070 16436 5122
rect 16380 5058 16436 5070
rect 15820 4958 15822 5010
rect 15874 4958 15876 5010
rect 15820 4946 15876 4958
rect 16268 5012 16324 5022
rect 15708 4732 16212 4788
rect 15484 4620 15764 4676
rect 15484 4452 15540 4462
rect 15484 3442 15540 4396
rect 15484 3390 15486 3442
rect 15538 3390 15540 3442
rect 15484 3378 15540 3390
rect 15708 3554 15764 4620
rect 15708 3502 15710 3554
rect 15762 3502 15764 3554
rect 15708 3444 15764 3502
rect 15932 3780 15988 3790
rect 15932 3388 15988 3724
rect 16156 3778 16212 4732
rect 16156 3726 16158 3778
rect 16210 3726 16212 3778
rect 16156 3714 16212 3726
rect 16268 3666 16324 4956
rect 16268 3614 16270 3666
rect 16322 3614 16324 3666
rect 16268 3602 16324 3614
rect 15708 3378 15764 3388
rect 15820 3332 15988 3388
rect 15820 3220 15876 3332
rect 16492 3220 16548 5516
rect 15708 3164 15876 3220
rect 16156 3164 16548 3220
rect 16604 5460 16660 5470
rect 15708 800 15764 3164
rect 16156 800 16212 3164
rect 16604 800 16660 5404
rect 16716 5348 16772 5854
rect 16716 5282 16772 5292
rect 16828 5122 16884 5134
rect 16828 5070 16830 5122
rect 16882 5070 16884 5122
rect 16716 4450 16772 4462
rect 16716 4398 16718 4450
rect 16770 4398 16772 4450
rect 16716 3444 16772 4398
rect 16828 4340 16884 5070
rect 16828 4274 16884 4284
rect 16828 3556 16884 3566
rect 16828 3462 16884 3500
rect 16940 3554 16996 6748
rect 17052 5012 17108 7980
rect 17388 7970 17444 7980
rect 17172 7868 17436 7878
rect 17228 7812 17276 7868
rect 17332 7812 17380 7868
rect 17172 7802 17436 7812
rect 17276 7474 17332 7486
rect 17276 7422 17278 7474
rect 17330 7422 17332 7474
rect 17276 6468 17332 7422
rect 17612 7474 17668 7486
rect 17612 7422 17614 7474
rect 17666 7422 17668 7474
rect 17500 7364 17556 7374
rect 17500 7270 17556 7308
rect 17612 6916 17668 7422
rect 17388 6860 17668 6916
rect 17836 7474 17892 7486
rect 17836 7422 17838 7474
rect 17890 7422 17892 7474
rect 17388 6692 17444 6860
rect 17388 6626 17444 6636
rect 17836 6468 17892 7422
rect 17276 6402 17332 6412
rect 17500 6412 17892 6468
rect 17948 7476 18004 11732
rect 19888 11732 19936 11788
rect 19992 11732 20040 11788
rect 19832 11722 20096 11732
rect 20300 11172 20356 15820
rect 20972 15810 21028 15820
rect 22204 15090 22260 17276
rect 22492 15708 22756 15718
rect 22548 15652 22596 15708
rect 22652 15652 22700 15708
rect 22492 15642 22756 15652
rect 22204 15038 22206 15090
rect 22258 15038 22260 15090
rect 22204 15026 22260 15038
rect 22492 14140 22756 14150
rect 22548 14084 22596 14140
rect 22652 14084 22700 14140
rect 22492 14074 22756 14084
rect 22204 12850 22260 12862
rect 22204 12798 22206 12850
rect 22258 12798 22260 12850
rect 21084 12740 21140 12750
rect 20300 11106 20356 11116
rect 20972 12684 21084 12740
rect 19832 10220 20096 10230
rect 19888 10164 19936 10220
rect 19992 10164 20040 10220
rect 19832 10154 20096 10164
rect 20860 9602 20916 9614
rect 20860 9550 20862 9602
rect 20914 9550 20916 9602
rect 20076 8930 20132 8942
rect 20076 8878 20078 8930
rect 20130 8878 20132 8930
rect 20076 8820 20132 8878
rect 20524 8932 20580 8942
rect 20524 8930 20692 8932
rect 20524 8878 20526 8930
rect 20578 8878 20692 8930
rect 20524 8876 20692 8878
rect 20524 8866 20580 8876
rect 19292 8764 20132 8820
rect 18060 8034 18116 8046
rect 18060 7982 18062 8034
rect 18114 7982 18116 8034
rect 18060 7476 18116 7982
rect 18508 8034 18564 8046
rect 18508 7982 18510 8034
rect 18562 7982 18564 8034
rect 18396 7476 18452 7486
rect 18060 7474 18452 7476
rect 18060 7422 18398 7474
rect 18450 7422 18452 7474
rect 18060 7420 18452 7422
rect 17172 6300 17436 6310
rect 17228 6244 17276 6300
rect 17332 6244 17380 6300
rect 17172 6234 17436 6244
rect 17388 6132 17444 6142
rect 17388 6038 17444 6076
rect 17500 6130 17556 6412
rect 17500 6078 17502 6130
rect 17554 6078 17556 6130
rect 17500 6066 17556 6078
rect 17612 6244 17668 6254
rect 17612 6130 17668 6188
rect 17948 6244 18004 7420
rect 17948 6178 18004 6188
rect 18172 6692 18228 6702
rect 17612 6078 17614 6130
rect 17666 6078 17668 6130
rect 17612 6066 17668 6078
rect 17836 6020 17892 6030
rect 17836 5926 17892 5964
rect 18060 6020 18116 6030
rect 17836 5796 17892 5806
rect 17500 5124 17556 5134
rect 17164 5012 17220 5022
rect 17052 4956 17164 5012
rect 17164 4946 17220 4956
rect 17172 4732 17436 4742
rect 17228 4676 17276 4732
rect 17332 4676 17380 4732
rect 17172 4666 17436 4676
rect 17500 4564 17556 5068
rect 16940 3502 16942 3554
rect 16994 3502 16996 3554
rect 16940 3490 16996 3502
rect 17164 4508 17556 4564
rect 16716 3378 16772 3388
rect 17164 3332 17220 4508
rect 17500 4338 17556 4350
rect 17500 4286 17502 4338
rect 17554 4286 17556 4338
rect 17500 4228 17556 4286
rect 17500 4162 17556 4172
rect 17836 3388 17892 5740
rect 18060 5684 18116 5964
rect 17052 3276 17220 3332
rect 17500 3332 17892 3388
rect 17948 5628 18116 5684
rect 17052 800 17108 3276
rect 17172 3164 17436 3174
rect 17228 3108 17276 3164
rect 17332 3108 17380 3164
rect 17172 3098 17436 3108
rect 17500 800 17556 3332
rect 17948 800 18004 5628
rect 18060 5348 18116 5358
rect 18060 4450 18116 5292
rect 18172 5124 18228 6636
rect 18284 6580 18340 6590
rect 18284 5794 18340 6524
rect 18284 5742 18286 5794
rect 18338 5742 18340 5794
rect 18284 5730 18340 5742
rect 18284 5572 18340 5582
rect 18396 5572 18452 7420
rect 18340 5516 18452 5572
rect 18284 5506 18340 5516
rect 18172 5058 18228 5068
rect 18396 5124 18452 5134
rect 18396 5010 18452 5068
rect 18396 4958 18398 5010
rect 18450 4958 18452 5010
rect 18396 4946 18452 4958
rect 18060 4398 18062 4450
rect 18114 4398 18116 4450
rect 18060 4386 18116 4398
rect 18284 4900 18340 4910
rect 18284 2436 18340 4844
rect 18396 4788 18452 4798
rect 18396 3442 18452 4732
rect 18508 4452 18564 7982
rect 19068 8034 19124 8046
rect 19068 7982 19070 8034
rect 19122 7982 19124 8034
rect 19068 7700 19124 7982
rect 18732 7644 19124 7700
rect 18620 7586 18676 7598
rect 18620 7534 18622 7586
rect 18674 7534 18676 7586
rect 18620 7140 18676 7534
rect 18620 7074 18676 7084
rect 18508 4386 18564 4396
rect 18620 6916 18676 6926
rect 18620 3780 18676 6860
rect 18732 5460 18788 7644
rect 18956 7476 19012 7486
rect 18732 5394 18788 5404
rect 18844 6580 18900 6590
rect 18732 5236 18788 5246
rect 18732 5010 18788 5180
rect 18732 4958 18734 5010
rect 18786 4958 18788 5010
rect 18732 4946 18788 4958
rect 18732 3780 18788 3790
rect 18620 3724 18732 3780
rect 18732 3714 18788 3724
rect 18396 3390 18398 3442
rect 18450 3390 18452 3442
rect 18396 3378 18452 3390
rect 18284 2380 18452 2436
rect 18396 800 18452 2380
rect 18844 800 18900 6524
rect 18956 3220 19012 7420
rect 19068 7362 19124 7374
rect 19068 7310 19070 7362
rect 19122 7310 19124 7362
rect 19068 6692 19124 7310
rect 19180 6916 19236 6926
rect 19292 6916 19348 8764
rect 19832 8652 20096 8662
rect 19888 8596 19936 8652
rect 19992 8596 20040 8652
rect 19832 8586 20096 8596
rect 19516 8036 19572 8046
rect 19516 8034 19684 8036
rect 19516 7982 19518 8034
rect 19570 7982 19684 8034
rect 19516 7980 19684 7982
rect 19516 7970 19572 7980
rect 19516 7362 19572 7374
rect 19516 7310 19518 7362
rect 19570 7310 19572 7362
rect 19236 6860 19348 6916
rect 19404 7250 19460 7262
rect 19404 7198 19406 7250
rect 19458 7198 19460 7250
rect 19180 6850 19236 6860
rect 19292 6692 19348 6702
rect 19068 6690 19348 6692
rect 19068 6638 19294 6690
rect 19346 6638 19348 6690
rect 19068 6636 19348 6638
rect 19068 6466 19124 6478
rect 19068 6414 19070 6466
rect 19122 6414 19124 6466
rect 19068 5460 19124 6414
rect 19292 5796 19348 6636
rect 19404 5908 19460 7198
rect 19516 6132 19572 7310
rect 19628 6356 19684 7980
rect 19852 8034 19908 8046
rect 20412 8036 20468 8046
rect 19852 7982 19854 8034
rect 19906 7982 19908 8034
rect 19852 7250 19908 7982
rect 20188 8034 20468 8036
rect 20188 7982 20414 8034
rect 20466 7982 20468 8034
rect 20188 7980 20468 7982
rect 20188 7588 20244 7980
rect 20412 7970 20468 7980
rect 20076 7476 20132 7486
rect 20076 7382 20132 7420
rect 19852 7198 19854 7250
rect 19906 7198 19908 7250
rect 19852 7186 19908 7198
rect 19832 7084 20096 7094
rect 19888 7028 19936 7084
rect 19992 7028 20040 7084
rect 19832 7018 20096 7028
rect 19740 6804 19796 6814
rect 19740 6578 19796 6748
rect 19740 6526 19742 6578
rect 19794 6526 19796 6578
rect 19740 6514 19796 6526
rect 19964 6690 20020 6702
rect 19964 6638 19966 6690
rect 20018 6638 20020 6690
rect 19964 6356 20020 6638
rect 19628 6300 20020 6356
rect 19516 6066 19572 6076
rect 19964 6020 20020 6300
rect 19964 5954 20020 5964
rect 19404 5842 19460 5852
rect 19292 5730 19348 5740
rect 19832 5516 20096 5526
rect 19628 5460 19684 5470
rect 19068 5404 19572 5460
rect 19292 5236 19348 5246
rect 19180 5180 19292 5236
rect 19068 5122 19124 5134
rect 19068 5070 19070 5122
rect 19122 5070 19124 5122
rect 19068 4452 19124 5070
rect 19068 4386 19124 4396
rect 19180 3554 19236 5180
rect 19292 5170 19348 5180
rect 19404 5124 19460 5134
rect 19404 5010 19460 5068
rect 19404 4958 19406 5010
rect 19458 4958 19460 5010
rect 19404 4946 19460 4958
rect 19516 4338 19572 5404
rect 19888 5460 19936 5516
rect 19992 5460 20040 5516
rect 19832 5450 20096 5460
rect 19628 5348 19684 5404
rect 19628 5292 20132 5348
rect 19740 5124 19796 5134
rect 19740 5030 19796 5068
rect 20076 5122 20132 5292
rect 20076 5070 20078 5122
rect 20130 5070 20132 5122
rect 20076 5058 20132 5070
rect 19516 4286 19518 4338
rect 19570 4286 19572 4338
rect 19516 4274 19572 4286
rect 19628 5012 19684 5022
rect 19180 3502 19182 3554
rect 19234 3502 19236 3554
rect 19180 3490 19236 3502
rect 19292 4226 19348 4238
rect 19292 4174 19294 4226
rect 19346 4174 19348 4226
rect 19292 3442 19348 4174
rect 19292 3390 19294 3442
rect 19346 3390 19348 3442
rect 19292 3378 19348 3390
rect 19628 3388 19684 4956
rect 20188 4900 20244 7532
rect 20412 7588 20468 7598
rect 20412 7586 20580 7588
rect 20412 7534 20414 7586
rect 20466 7534 20580 7586
rect 20412 7532 20580 7534
rect 20412 7522 20468 7532
rect 20412 6916 20468 6926
rect 20188 4834 20244 4844
rect 20300 6860 20412 6916
rect 20300 4788 20356 6860
rect 20412 6850 20468 6860
rect 20412 6580 20468 6590
rect 20412 6486 20468 6524
rect 20412 6132 20468 6142
rect 20412 6018 20468 6076
rect 20412 5966 20414 6018
rect 20466 5966 20468 6018
rect 20412 5572 20468 5966
rect 20524 5796 20580 7532
rect 20636 7028 20692 8876
rect 20860 8818 20916 9550
rect 20860 8766 20862 8818
rect 20914 8766 20916 8818
rect 20860 8754 20916 8766
rect 20748 8034 20804 8046
rect 20748 7982 20750 8034
rect 20802 7982 20804 8034
rect 20748 7476 20804 7982
rect 20860 7588 20916 7598
rect 20972 7588 21028 12684
rect 21084 12674 21140 12684
rect 21644 12738 21700 12750
rect 21644 12686 21646 12738
rect 21698 12686 21700 12738
rect 21644 12404 21700 12686
rect 21868 12740 21924 12750
rect 21868 12646 21924 12684
rect 21644 12338 21700 12348
rect 22204 12404 22260 12798
rect 22492 12572 22756 12582
rect 22548 12516 22596 12572
rect 22652 12516 22700 12572
rect 22492 12506 22756 12516
rect 22204 12338 22260 12348
rect 22492 11004 22756 11014
rect 22548 10948 22596 11004
rect 22652 10948 22700 11004
rect 22492 10938 22756 10948
rect 22204 9604 22260 9614
rect 22204 9510 22260 9548
rect 22492 9436 22756 9446
rect 22548 9380 22596 9436
rect 22652 9380 22700 9436
rect 22492 9370 22756 9380
rect 21420 9100 21812 9156
rect 20860 7586 21028 7588
rect 20860 7534 20862 7586
rect 20914 7534 21028 7586
rect 20860 7532 21028 7534
rect 21084 8930 21140 8942
rect 21084 8878 21086 8930
rect 21138 8878 21140 8930
rect 20860 7522 20916 7532
rect 20748 7410 20804 7420
rect 20748 7252 20804 7262
rect 20748 7158 20804 7196
rect 20636 6972 20916 7028
rect 20524 5730 20580 5740
rect 20636 6468 20692 6478
rect 20412 5516 20580 5572
rect 20412 5348 20468 5358
rect 20412 5010 20468 5292
rect 20412 4958 20414 5010
rect 20466 4958 20468 5010
rect 20412 4946 20468 4958
rect 20300 4722 20356 4732
rect 20524 4564 20580 5516
rect 20524 4498 20580 4508
rect 19832 3948 20096 3958
rect 19888 3892 19936 3948
rect 19992 3892 20040 3948
rect 19832 3882 20096 3892
rect 19628 3332 19796 3388
rect 18956 3164 19348 3220
rect 19292 800 19348 3164
rect 19740 800 19796 3332
rect 20188 2994 20244 3006
rect 20188 2942 20190 2994
rect 20242 2942 20244 2994
rect 20188 800 20244 2942
rect 20636 800 20692 6412
rect 20748 6466 20804 6478
rect 20748 6414 20750 6466
rect 20802 6414 20804 6466
rect 20748 5124 20804 6414
rect 20748 5058 20804 5068
rect 20860 3668 20916 6972
rect 20972 6468 21028 6478
rect 21084 6468 21140 8878
rect 21420 8818 21476 9100
rect 21532 8932 21588 8942
rect 21532 8930 21700 8932
rect 21532 8878 21534 8930
rect 21586 8878 21700 8930
rect 21532 8876 21700 8878
rect 21532 8866 21588 8876
rect 21420 8766 21422 8818
rect 21474 8766 21476 8818
rect 21420 8754 21476 8766
rect 21420 8034 21476 8046
rect 21420 7982 21422 8034
rect 21474 7982 21476 8034
rect 21196 7586 21252 7598
rect 21196 7534 21198 7586
rect 21250 7534 21252 7586
rect 21196 6916 21252 7534
rect 21196 6850 21252 6860
rect 21308 6578 21364 6590
rect 21308 6526 21310 6578
rect 21362 6526 21364 6578
rect 21308 6468 21364 6526
rect 21028 6412 21364 6468
rect 20972 6402 21028 6412
rect 21420 6244 21476 7982
rect 21532 7588 21588 7598
rect 21532 7494 21588 7532
rect 21644 6692 21700 8876
rect 21756 8146 21812 9100
rect 22316 8932 22372 8942
rect 21756 8094 21758 8146
rect 21810 8094 21812 8146
rect 21756 6916 21812 8094
rect 22092 8930 22372 8932
rect 22092 8878 22318 8930
rect 22370 8878 22372 8930
rect 22092 8876 22372 8878
rect 21868 7588 21924 7598
rect 21868 7586 22036 7588
rect 21868 7534 21870 7586
rect 21922 7534 22036 7586
rect 21868 7532 22036 7534
rect 21868 7522 21924 7532
rect 21756 6850 21812 6860
rect 21644 6636 21812 6692
rect 20972 6188 21476 6244
rect 21644 6466 21700 6478
rect 21644 6414 21646 6466
rect 21698 6414 21700 6466
rect 20972 4452 21028 6188
rect 21532 6020 21588 6030
rect 21196 6018 21588 6020
rect 21196 5966 21534 6018
rect 21586 5966 21588 6018
rect 21196 5964 21588 5966
rect 21196 5906 21252 5964
rect 21532 5954 21588 5964
rect 21196 5854 21198 5906
rect 21250 5854 21252 5906
rect 21196 5842 21252 5854
rect 21420 5796 21476 5806
rect 21476 5740 21588 5796
rect 21420 5730 21476 5740
rect 21420 5236 21476 5246
rect 21420 5142 21476 5180
rect 21308 5124 21364 5134
rect 21308 5030 21364 5068
rect 21532 5010 21588 5740
rect 21532 4958 21534 5010
rect 21586 4958 21588 5010
rect 21532 4946 21588 4958
rect 21084 4452 21140 4462
rect 20972 4450 21140 4452
rect 20972 4398 21086 4450
rect 21138 4398 21140 4450
rect 20972 4396 21140 4398
rect 21084 4386 21140 4396
rect 21420 4340 21476 4350
rect 20972 3668 21028 3678
rect 20860 3612 20972 3668
rect 20972 3554 21028 3612
rect 20972 3502 20974 3554
rect 21026 3502 21028 3554
rect 20972 3490 21028 3502
rect 20748 3444 20804 3482
rect 20748 3378 20804 3388
rect 21420 3442 21476 4284
rect 21644 4338 21700 6414
rect 21644 4286 21646 4338
rect 21698 4286 21700 4338
rect 21644 4274 21700 4286
rect 21756 5906 21812 6636
rect 21756 5854 21758 5906
rect 21810 5854 21812 5906
rect 21532 3780 21588 3790
rect 21532 3556 21588 3724
rect 21644 3556 21700 3566
rect 21532 3554 21700 3556
rect 21532 3502 21646 3554
rect 21698 3502 21700 3554
rect 21532 3500 21700 3502
rect 21644 3490 21700 3500
rect 21420 3390 21422 3442
rect 21474 3390 21476 3442
rect 21420 3378 21476 3390
rect 21756 2994 21812 5854
rect 21868 5684 21924 5694
rect 21868 5124 21924 5628
rect 21980 5236 22036 7532
rect 22092 7476 22148 8876
rect 22316 8866 22372 8876
rect 22204 8036 22260 8046
rect 22204 8034 22372 8036
rect 22204 7982 22206 8034
rect 22258 7982 22372 8034
rect 22204 7980 22372 7982
rect 22204 7970 22260 7980
rect 22204 7476 22260 7486
rect 22092 7474 22260 7476
rect 22092 7422 22206 7474
rect 22258 7422 22260 7474
rect 22092 7420 22260 7422
rect 22316 7476 22372 7980
rect 22492 7868 22756 7878
rect 22548 7812 22596 7868
rect 22652 7812 22700 7868
rect 22492 7802 22756 7812
rect 22428 7476 22484 7486
rect 22316 7420 22428 7476
rect 22204 6804 22260 7420
rect 22428 7410 22484 7420
rect 22204 6748 22372 6804
rect 22092 6580 22148 6590
rect 22092 6486 22148 6524
rect 22092 5236 22148 5246
rect 21980 5234 22148 5236
rect 21980 5182 22094 5234
rect 22146 5182 22148 5234
rect 21980 5180 22148 5182
rect 22092 5170 22148 5180
rect 21868 5068 22036 5124
rect 21980 5010 22036 5068
rect 21980 4958 21982 5010
rect 22034 4958 22036 5010
rect 21980 4946 22036 4958
rect 21868 4564 21924 4574
rect 21868 4452 21924 4508
rect 21868 4450 22260 4452
rect 21868 4398 21870 4450
rect 21922 4398 22260 4450
rect 21868 4396 22260 4398
rect 21868 4386 21924 4396
rect 22204 3666 22260 4396
rect 22204 3614 22206 3666
rect 22258 3614 22260 3666
rect 22204 3602 22260 3614
rect 21756 2942 21758 2994
rect 21810 2942 21812 2994
rect 21756 2930 21812 2942
rect 22316 2548 22372 6748
rect 22492 6300 22756 6310
rect 22548 6244 22596 6300
rect 22652 6244 22700 6300
rect 22492 6234 22756 6244
rect 22492 4732 22756 4742
rect 22548 4676 22596 4732
rect 22652 4676 22700 4732
rect 22492 4666 22756 4676
rect 22492 3164 22756 3174
rect 22548 3108 22596 3164
rect 22652 3108 22700 3164
rect 22492 3098 22756 3108
rect 22316 2482 22372 2492
rect 3136 0 3248 800
rect 3584 0 3696 800
rect 4032 0 4144 800
rect 4480 0 4592 800
rect 4928 0 5040 800
rect 5376 0 5488 800
rect 5824 0 5936 800
rect 6272 0 6384 800
rect 6720 0 6832 800
rect 7168 0 7280 800
rect 7616 0 7728 800
rect 8064 0 8176 800
rect 8512 0 8624 800
rect 8960 0 9072 800
rect 9408 0 9520 800
rect 9856 0 9968 800
rect 10304 0 10416 800
rect 10752 0 10864 800
rect 11200 0 11312 800
rect 11648 0 11760 800
rect 12096 0 12208 800
rect 12544 0 12656 800
rect 12992 0 13104 800
rect 13440 0 13552 800
rect 13888 0 14000 800
rect 14336 0 14448 800
rect 14784 0 14896 800
rect 15232 0 15344 800
rect 15680 0 15792 800
rect 16128 0 16240 800
rect 16576 0 16688 800
rect 17024 0 17136 800
rect 17472 0 17584 800
rect 17920 0 18032 800
rect 18368 0 18480 800
rect 18816 0 18928 800
rect 19264 0 19376 800
rect 19712 0 19824 800
rect 20160 0 20272 800
rect 20608 0 20720 800
<< via2 >>
rect 3500 17276 3556 17332
rect 3052 16380 3108 16436
rect 2380 15932 2436 15988
rect 3388 15484 3444 15540
rect 3612 16828 3668 16884
rect 3872 16490 3928 16492
rect 3872 16438 3874 16490
rect 3874 16438 3926 16490
rect 3926 16438 3928 16490
rect 3872 16436 3928 16438
rect 3976 16490 4032 16492
rect 3976 16438 3978 16490
rect 3978 16438 4030 16490
rect 4030 16438 4032 16490
rect 3976 16436 4032 16438
rect 4080 16490 4136 16492
rect 4080 16438 4082 16490
rect 4082 16438 4134 16490
rect 4134 16438 4136 16490
rect 4080 16436 4136 16438
rect 9192 16490 9248 16492
rect 9192 16438 9194 16490
rect 9194 16438 9246 16490
rect 9246 16438 9248 16490
rect 9192 16436 9248 16438
rect 9296 16490 9352 16492
rect 9296 16438 9298 16490
rect 9298 16438 9350 16490
rect 9350 16438 9352 16490
rect 9296 16436 9352 16438
rect 9400 16490 9456 16492
rect 9400 16438 9402 16490
rect 9402 16438 9454 16490
rect 9454 16438 9456 16490
rect 9400 16436 9456 16438
rect 14512 16490 14568 16492
rect 14512 16438 14514 16490
rect 14514 16438 14566 16490
rect 14566 16438 14568 16490
rect 14512 16436 14568 16438
rect 14616 16490 14672 16492
rect 14616 16438 14618 16490
rect 14618 16438 14670 16490
rect 14670 16438 14672 16490
rect 14616 16436 14672 16438
rect 14720 16490 14776 16492
rect 14720 16438 14722 16490
rect 14722 16438 14774 16490
rect 14774 16438 14776 16490
rect 14720 16436 14776 16438
rect 16156 16268 16212 16324
rect 17052 16268 17108 16324
rect 19832 16490 19888 16492
rect 19832 16438 19834 16490
rect 19834 16438 19886 16490
rect 19886 16438 19888 16490
rect 19832 16436 19888 16438
rect 19936 16490 19992 16492
rect 19936 16438 19938 16490
rect 19938 16438 19990 16490
rect 19990 16438 19992 16490
rect 19936 16436 19992 16438
rect 20040 16490 20096 16492
rect 20040 16438 20042 16490
rect 20042 16438 20094 16490
rect 20094 16438 20096 16490
rect 20040 16436 20096 16438
rect 22204 17276 22260 17332
rect 8764 15820 8820 15876
rect 9436 15874 9492 15876
rect 9436 15822 9438 15874
rect 9438 15822 9490 15874
rect 9490 15822 9492 15874
rect 9436 15820 9492 15822
rect 15932 15820 15988 15876
rect 6532 15706 6588 15708
rect 6532 15654 6534 15706
rect 6534 15654 6586 15706
rect 6586 15654 6588 15706
rect 6532 15652 6588 15654
rect 6636 15706 6692 15708
rect 6636 15654 6638 15706
rect 6638 15654 6690 15706
rect 6690 15654 6692 15706
rect 6636 15652 6692 15654
rect 6740 15706 6796 15708
rect 6740 15654 6742 15706
rect 6742 15654 6794 15706
rect 6794 15654 6796 15706
rect 6740 15652 6796 15654
rect 11852 15706 11908 15708
rect 11852 15654 11854 15706
rect 11854 15654 11906 15706
rect 11906 15654 11908 15706
rect 11852 15652 11908 15654
rect 11956 15706 12012 15708
rect 11956 15654 11958 15706
rect 11958 15654 12010 15706
rect 12010 15654 12012 15706
rect 11956 15652 12012 15654
rect 12060 15706 12116 15708
rect 12060 15654 12062 15706
rect 12062 15654 12114 15706
rect 12114 15654 12116 15706
rect 12060 15652 12116 15654
rect 2156 15036 2212 15092
rect 1708 14924 1764 14980
rect 2156 14306 2212 14308
rect 2156 14254 2158 14306
rect 2158 14254 2210 14306
rect 2210 14254 2212 14306
rect 2156 14252 2212 14254
rect 1708 14028 1764 14084
rect 1708 13244 1764 13300
rect 1708 12850 1764 12852
rect 1708 12798 1710 12850
rect 1710 12798 1762 12850
rect 1762 12798 1764 12850
rect 1708 12796 1764 12798
rect 2156 12738 2212 12740
rect 2156 12686 2158 12738
rect 2158 12686 2210 12738
rect 2210 12686 2212 12738
rect 2156 12684 2212 12686
rect 1708 11900 1764 11956
rect 3872 14922 3928 14924
rect 3872 14870 3874 14922
rect 3874 14870 3926 14922
rect 3926 14870 3928 14922
rect 3872 14868 3928 14870
rect 3976 14922 4032 14924
rect 3976 14870 3978 14922
rect 3978 14870 4030 14922
rect 4030 14870 4032 14922
rect 3976 14868 4032 14870
rect 4080 14922 4136 14924
rect 4080 14870 4082 14922
rect 4082 14870 4134 14922
rect 4134 14870 4136 14922
rect 4080 14868 4136 14870
rect 9192 14922 9248 14924
rect 9192 14870 9194 14922
rect 9194 14870 9246 14922
rect 9246 14870 9248 14922
rect 9192 14868 9248 14870
rect 9296 14922 9352 14924
rect 9296 14870 9298 14922
rect 9298 14870 9350 14922
rect 9350 14870 9352 14922
rect 9296 14868 9352 14870
rect 9400 14922 9456 14924
rect 9400 14870 9402 14922
rect 9402 14870 9454 14922
rect 9454 14870 9456 14922
rect 9400 14868 9456 14870
rect 14512 14922 14568 14924
rect 14512 14870 14514 14922
rect 14514 14870 14566 14922
rect 14566 14870 14568 14922
rect 14512 14868 14568 14870
rect 14616 14922 14672 14924
rect 14616 14870 14618 14922
rect 14618 14870 14670 14922
rect 14670 14870 14672 14922
rect 14616 14868 14672 14870
rect 14720 14922 14776 14924
rect 14720 14870 14722 14922
rect 14722 14870 14774 14922
rect 14774 14870 14776 14922
rect 14720 14868 14776 14870
rect 6532 14138 6588 14140
rect 6532 14086 6534 14138
rect 6534 14086 6586 14138
rect 6586 14086 6588 14138
rect 6532 14084 6588 14086
rect 6636 14138 6692 14140
rect 6636 14086 6638 14138
rect 6638 14086 6690 14138
rect 6690 14086 6692 14138
rect 6636 14084 6692 14086
rect 6740 14138 6796 14140
rect 6740 14086 6742 14138
rect 6742 14086 6794 14138
rect 6794 14086 6796 14138
rect 6740 14084 6796 14086
rect 11852 14138 11908 14140
rect 11852 14086 11854 14138
rect 11854 14086 11906 14138
rect 11906 14086 11908 14138
rect 11852 14084 11908 14086
rect 11956 14138 12012 14140
rect 11956 14086 11958 14138
rect 11958 14086 12010 14138
rect 12010 14086 12012 14138
rect 11956 14084 12012 14086
rect 12060 14138 12116 14140
rect 12060 14086 12062 14138
rect 12062 14086 12114 14138
rect 12114 14086 12116 14138
rect 12060 14084 12116 14086
rect 3872 13354 3928 13356
rect 3872 13302 3874 13354
rect 3874 13302 3926 13354
rect 3926 13302 3928 13354
rect 3872 13300 3928 13302
rect 3976 13354 4032 13356
rect 3976 13302 3978 13354
rect 3978 13302 4030 13354
rect 4030 13302 4032 13354
rect 3976 13300 4032 13302
rect 4080 13354 4136 13356
rect 4080 13302 4082 13354
rect 4082 13302 4134 13354
rect 4134 13302 4136 13354
rect 4080 13300 4136 13302
rect 9192 13354 9248 13356
rect 9192 13302 9194 13354
rect 9194 13302 9246 13354
rect 9246 13302 9248 13354
rect 9192 13300 9248 13302
rect 9296 13354 9352 13356
rect 9296 13302 9298 13354
rect 9298 13302 9350 13354
rect 9350 13302 9352 13354
rect 9296 13300 9352 13302
rect 9400 13354 9456 13356
rect 9400 13302 9402 13354
rect 9402 13302 9454 13354
rect 9454 13302 9456 13354
rect 9400 13300 9456 13302
rect 14512 13354 14568 13356
rect 14512 13302 14514 13354
rect 14514 13302 14566 13354
rect 14566 13302 14568 13354
rect 14512 13300 14568 13302
rect 14616 13354 14672 13356
rect 14616 13302 14618 13354
rect 14618 13302 14670 13354
rect 14670 13302 14672 13354
rect 14616 13300 14672 13302
rect 14720 13354 14776 13356
rect 14720 13302 14722 13354
rect 14722 13302 14774 13354
rect 14774 13302 14776 13354
rect 14720 13300 14776 13302
rect 6532 12570 6588 12572
rect 6532 12518 6534 12570
rect 6534 12518 6586 12570
rect 6586 12518 6588 12570
rect 6532 12516 6588 12518
rect 6636 12570 6692 12572
rect 6636 12518 6638 12570
rect 6638 12518 6690 12570
rect 6690 12518 6692 12570
rect 6636 12516 6692 12518
rect 6740 12570 6796 12572
rect 6740 12518 6742 12570
rect 6742 12518 6794 12570
rect 6794 12518 6796 12570
rect 6740 12516 6796 12518
rect 11852 12570 11908 12572
rect 11852 12518 11854 12570
rect 11854 12518 11906 12570
rect 11906 12518 11908 12570
rect 11852 12516 11908 12518
rect 11956 12570 12012 12572
rect 11956 12518 11958 12570
rect 11958 12518 12010 12570
rect 12010 12518 12012 12570
rect 11956 12516 12012 12518
rect 12060 12570 12116 12572
rect 12060 12518 12062 12570
rect 12062 12518 12114 12570
rect 12114 12518 12116 12570
rect 12060 12516 12116 12518
rect 2156 11452 2212 11508
rect 1708 11170 1764 11172
rect 1708 11118 1710 11170
rect 1710 11118 1762 11170
rect 1762 11118 1764 11170
rect 1708 11116 1764 11118
rect 2044 10556 2100 10612
rect 1708 10108 1764 10164
rect 1708 9602 1764 9604
rect 1708 9550 1710 9602
rect 1710 9550 1762 9602
rect 1762 9550 1764 9602
rect 1708 9548 1764 9550
rect 2492 11116 2548 11172
rect 2156 9212 2212 9268
rect 2044 9100 2100 9156
rect 1820 8428 1876 8484
rect 1932 8540 1988 8596
rect 1820 7868 1876 7924
rect 1820 7644 1876 7700
rect 1708 7532 1764 7588
rect 1484 4508 1540 4564
rect 1708 6076 1764 6132
rect 2268 8540 2324 8596
rect 2492 8764 2548 8820
rect 3724 12012 3780 12068
rect 3872 11786 3928 11788
rect 3872 11734 3874 11786
rect 3874 11734 3926 11786
rect 3926 11734 3928 11786
rect 3872 11732 3928 11734
rect 3976 11786 4032 11788
rect 3976 11734 3978 11786
rect 3978 11734 4030 11786
rect 4030 11734 4032 11786
rect 3976 11732 4032 11734
rect 4080 11786 4136 11788
rect 4080 11734 4082 11786
rect 4082 11734 4134 11786
rect 4134 11734 4136 11786
rect 4080 11732 4136 11734
rect 3388 11170 3444 11172
rect 3388 11118 3390 11170
rect 3390 11118 3442 11170
rect 3442 11118 3444 11170
rect 3388 11116 3444 11118
rect 2716 9324 2772 9380
rect 2716 9154 2772 9156
rect 2716 9102 2718 9154
rect 2718 9102 2770 9154
rect 2770 9102 2772 9154
rect 2716 9100 2772 9102
rect 2604 8428 2660 8484
rect 3724 10556 3780 10612
rect 2940 8428 2996 8484
rect 2156 7308 2212 7364
rect 3388 9324 3444 9380
rect 3276 9154 3332 9156
rect 3276 9102 3278 9154
rect 3278 9102 3330 9154
rect 3330 9102 3332 9154
rect 3276 9100 3332 9102
rect 2380 7756 2436 7812
rect 2716 8034 2772 8036
rect 2716 7982 2718 8034
rect 2718 7982 2770 8034
rect 2770 7982 2772 8034
rect 2716 7980 2772 7982
rect 2940 7868 2996 7924
rect 3052 7644 3108 7700
rect 1932 6412 1988 6468
rect 2268 6076 2324 6132
rect 2156 5794 2212 5796
rect 2156 5742 2158 5794
rect 2158 5742 2210 5794
rect 2210 5742 2212 5794
rect 2156 5740 2212 5742
rect 1932 5292 1988 5348
rect 1820 4732 1876 4788
rect 2828 6300 2884 6356
rect 2940 6076 2996 6132
rect 2604 4620 2660 4676
rect 2716 5068 2772 5124
rect 2492 4284 2548 4340
rect 1932 3778 1988 3780
rect 1932 3726 1934 3778
rect 1934 3726 1986 3778
rect 1986 3726 1988 3778
rect 1932 3724 1988 3726
rect 3872 10218 3928 10220
rect 3872 10166 3874 10218
rect 3874 10166 3926 10218
rect 3926 10166 3928 10218
rect 3872 10164 3928 10166
rect 3976 10218 4032 10220
rect 3976 10166 3978 10218
rect 3978 10166 4030 10218
rect 4030 10166 4032 10218
rect 3976 10164 4032 10166
rect 4080 10218 4136 10220
rect 4080 10166 4082 10218
rect 4082 10166 4134 10218
rect 4134 10166 4136 10218
rect 4080 10164 4136 10166
rect 3388 7084 3444 7140
rect 3276 5906 3332 5908
rect 3276 5854 3278 5906
rect 3278 5854 3330 5906
rect 3330 5854 3332 5906
rect 3276 5852 3332 5854
rect 2828 4396 2884 4452
rect 3276 5516 3332 5572
rect 3164 4284 3220 4340
rect 3052 3442 3108 3444
rect 3052 3390 3054 3442
rect 3054 3390 3106 3442
rect 3106 3390 3108 3442
rect 3052 3388 3108 3390
rect 2492 2940 2548 2996
rect 1708 2492 1764 2548
rect 4172 9602 4228 9604
rect 4172 9550 4174 9602
rect 4174 9550 4226 9602
rect 4226 9550 4228 9602
rect 4172 9548 4228 9550
rect 9192 11786 9248 11788
rect 9192 11734 9194 11786
rect 9194 11734 9246 11786
rect 9246 11734 9248 11786
rect 9192 11732 9248 11734
rect 9296 11786 9352 11788
rect 9296 11734 9298 11786
rect 9298 11734 9350 11786
rect 9350 11734 9352 11786
rect 9296 11732 9352 11734
rect 9400 11786 9456 11788
rect 9400 11734 9402 11786
rect 9402 11734 9454 11786
rect 9454 11734 9456 11786
rect 9400 11732 9456 11734
rect 14512 11786 14568 11788
rect 14512 11734 14514 11786
rect 14514 11734 14566 11786
rect 14566 11734 14568 11786
rect 14512 11732 14568 11734
rect 14616 11786 14672 11788
rect 14616 11734 14618 11786
rect 14618 11734 14670 11786
rect 14670 11734 14672 11786
rect 14616 11732 14672 11734
rect 14720 11786 14776 11788
rect 14720 11734 14722 11786
rect 14722 11734 14774 11786
rect 14774 11734 14776 11786
rect 14720 11732 14776 11734
rect 4956 11506 5012 11508
rect 4956 11454 4958 11506
rect 4958 11454 5010 11506
rect 5010 11454 5012 11506
rect 4956 11452 5012 11454
rect 9996 11170 10052 11172
rect 9996 11118 9998 11170
rect 9998 11118 10050 11170
rect 10050 11118 10052 11170
rect 9996 11116 10052 11118
rect 15148 11116 15204 11172
rect 4508 10892 4564 10948
rect 6532 11002 6588 11004
rect 6532 10950 6534 11002
rect 6534 10950 6586 11002
rect 6586 10950 6588 11002
rect 6532 10948 6588 10950
rect 6636 11002 6692 11004
rect 6636 10950 6638 11002
rect 6638 10950 6690 11002
rect 6690 10950 6692 11002
rect 6636 10948 6692 10950
rect 6740 11002 6796 11004
rect 6740 10950 6742 11002
rect 6742 10950 6794 11002
rect 6794 10950 6796 11002
rect 6740 10948 6796 10950
rect 11852 11002 11908 11004
rect 11852 10950 11854 11002
rect 11854 10950 11906 11002
rect 11906 10950 11908 11002
rect 11852 10948 11908 10950
rect 11956 11002 12012 11004
rect 11956 10950 11958 11002
rect 11958 10950 12010 11002
rect 12010 10950 12012 11002
rect 11956 10948 12012 10950
rect 12060 11002 12116 11004
rect 12060 10950 12062 11002
rect 12062 10950 12114 11002
rect 12114 10950 12116 11002
rect 12060 10948 12116 10950
rect 4396 9324 4452 9380
rect 3872 8650 3928 8652
rect 3872 8598 3874 8650
rect 3874 8598 3926 8650
rect 3926 8598 3928 8650
rect 3872 8596 3928 8598
rect 3976 8650 4032 8652
rect 3976 8598 3978 8650
rect 3978 8598 4030 8650
rect 4030 8598 4032 8650
rect 3976 8596 4032 8598
rect 4080 8650 4136 8652
rect 4080 8598 4082 8650
rect 4082 8598 4134 8650
rect 4134 8598 4136 8650
rect 4080 8596 4136 8598
rect 3612 8092 3668 8148
rect 3724 8034 3780 8036
rect 3724 7982 3726 8034
rect 3726 7982 3778 8034
rect 3778 7982 3780 8034
rect 3724 7980 3780 7982
rect 4060 7980 4116 8036
rect 3724 7532 3780 7588
rect 3836 7474 3892 7476
rect 3836 7422 3838 7474
rect 3838 7422 3890 7474
rect 3890 7422 3892 7474
rect 3836 7420 3892 7422
rect 3724 7196 3780 7252
rect 3872 7082 3928 7084
rect 3872 7030 3874 7082
rect 3874 7030 3926 7082
rect 3926 7030 3928 7082
rect 3872 7028 3928 7030
rect 3976 7082 4032 7084
rect 3976 7030 3978 7082
rect 3978 7030 4030 7082
rect 4030 7030 4032 7082
rect 3976 7028 4032 7030
rect 4080 7082 4136 7084
rect 4080 7030 4082 7082
rect 4082 7030 4134 7082
rect 4134 7030 4136 7082
rect 4080 7028 4136 7030
rect 4284 6972 4340 7028
rect 4844 9602 4900 9604
rect 4844 9550 4846 9602
rect 4846 9550 4898 9602
rect 4898 9550 4900 9602
rect 4844 9548 4900 9550
rect 4844 9100 4900 9156
rect 4844 8428 4900 8484
rect 4956 8876 5012 8932
rect 4844 8092 4900 8148
rect 3500 6636 3556 6692
rect 3500 4284 3556 4340
rect 4284 6412 4340 6468
rect 4172 5852 4228 5908
rect 3948 5740 4004 5796
rect 4284 5628 4340 5684
rect 3872 5514 3928 5516
rect 3872 5462 3874 5514
rect 3874 5462 3926 5514
rect 3926 5462 3928 5514
rect 3872 5460 3928 5462
rect 3976 5514 4032 5516
rect 3976 5462 3978 5514
rect 3978 5462 4030 5514
rect 4030 5462 4032 5514
rect 3976 5460 4032 5462
rect 4080 5514 4136 5516
rect 4080 5462 4082 5514
rect 4082 5462 4134 5514
rect 4134 5462 4136 5514
rect 4080 5460 4136 5462
rect 3948 5180 4004 5236
rect 4172 4898 4228 4900
rect 4172 4846 4174 4898
rect 4174 4846 4226 4898
rect 4226 4846 4228 4898
rect 4172 4844 4228 4846
rect 4060 4450 4116 4452
rect 4060 4398 4062 4450
rect 4062 4398 4114 4450
rect 4114 4398 4116 4450
rect 4060 4396 4116 4398
rect 3948 4172 4004 4228
rect 4284 4060 4340 4116
rect 3872 3946 3928 3948
rect 3872 3894 3874 3946
rect 3874 3894 3926 3946
rect 3926 3894 3928 3946
rect 3872 3892 3928 3894
rect 3976 3946 4032 3948
rect 3976 3894 3978 3946
rect 3978 3894 4030 3946
rect 4030 3894 4032 3946
rect 3976 3892 4032 3894
rect 4080 3946 4136 3948
rect 4080 3894 4082 3946
rect 4082 3894 4134 3946
rect 4134 3894 4136 3946
rect 4080 3892 4136 3894
rect 3724 3554 3780 3556
rect 3724 3502 3726 3554
rect 3726 3502 3778 3554
rect 3778 3502 3780 3554
rect 3724 3500 3780 3502
rect 4284 3554 4340 3556
rect 4284 3502 4286 3554
rect 4286 3502 4338 3554
rect 4338 3502 4340 3554
rect 4284 3500 4340 3502
rect 4732 7084 4788 7140
rect 4620 6524 4676 6580
rect 4844 6636 4900 6692
rect 4732 6018 4788 6020
rect 4732 5966 4734 6018
rect 4734 5966 4786 6018
rect 4786 5966 4788 6018
rect 4732 5964 4788 5966
rect 4508 5516 4564 5572
rect 4844 4956 4900 5012
rect 5180 7420 5236 7476
rect 5292 9212 5348 9268
rect 5068 7196 5124 7252
rect 5180 7084 5236 7140
rect 5068 6860 5124 6916
rect 5180 6636 5236 6692
rect 5180 5180 5236 5236
rect 5964 9324 6020 9380
rect 5404 8764 5460 8820
rect 5404 8316 5460 8372
rect 5404 7644 5460 7700
rect 5404 5740 5460 5796
rect 6532 9434 6588 9436
rect 6532 9382 6534 9434
rect 6534 9382 6586 9434
rect 6586 9382 6588 9434
rect 6532 9380 6588 9382
rect 6636 9434 6692 9436
rect 6636 9382 6638 9434
rect 6638 9382 6690 9434
rect 6690 9382 6692 9434
rect 6636 9380 6692 9382
rect 6740 9434 6796 9436
rect 6740 9382 6742 9434
rect 6742 9382 6794 9434
rect 6794 9382 6796 9434
rect 6740 9380 6796 9382
rect 5852 8930 5908 8932
rect 5852 8878 5854 8930
rect 5854 8878 5906 8930
rect 5906 8878 5908 8930
rect 5852 8876 5908 8878
rect 6188 8764 6244 8820
rect 5516 8092 5572 8148
rect 5404 4620 5460 4676
rect 4844 4060 4900 4116
rect 4732 3442 4788 3444
rect 4732 3390 4734 3442
rect 4734 3390 4786 3442
rect 4786 3390 4788 3442
rect 4732 3388 4788 3390
rect 5964 8204 6020 8260
rect 5740 8092 5796 8148
rect 6076 7532 6132 7588
rect 6300 8316 6356 8372
rect 6300 7756 6356 7812
rect 6860 8764 6916 8820
rect 6636 8540 6692 8596
rect 9192 10218 9248 10220
rect 9192 10166 9194 10218
rect 9194 10166 9246 10218
rect 9246 10166 9248 10218
rect 9192 10164 9248 10166
rect 9296 10218 9352 10220
rect 9296 10166 9298 10218
rect 9298 10166 9350 10218
rect 9350 10166 9352 10218
rect 9296 10164 9352 10166
rect 9400 10218 9456 10220
rect 9400 10166 9402 10218
rect 9402 10166 9454 10218
rect 9454 10166 9456 10218
rect 9400 10164 9456 10166
rect 7420 9602 7476 9604
rect 7420 9550 7422 9602
rect 7422 9550 7474 9602
rect 7474 9550 7476 9602
rect 7420 9548 7476 9550
rect 7084 9154 7140 9156
rect 7084 9102 7086 9154
rect 7086 9102 7138 9154
rect 7138 9102 7140 9154
rect 7084 9100 7140 9102
rect 8428 9602 8484 9604
rect 8428 9550 8430 9602
rect 8430 9550 8482 9602
rect 8482 9550 8484 9602
rect 8428 9548 8484 9550
rect 6972 8316 7028 8372
rect 7084 8876 7140 8932
rect 6636 8146 6692 8148
rect 6636 8094 6638 8146
rect 6638 8094 6690 8146
rect 6690 8094 6692 8146
rect 6636 8092 6692 8094
rect 6532 7866 6588 7868
rect 6532 7814 6534 7866
rect 6534 7814 6586 7866
rect 6586 7814 6588 7866
rect 6532 7812 6588 7814
rect 6636 7866 6692 7868
rect 6636 7814 6638 7866
rect 6638 7814 6690 7866
rect 6690 7814 6692 7866
rect 6636 7812 6692 7814
rect 6740 7866 6796 7868
rect 6740 7814 6742 7866
rect 6742 7814 6794 7866
rect 6794 7814 6796 7866
rect 6740 7812 6796 7814
rect 6076 6860 6132 6916
rect 6188 6748 6244 6804
rect 6860 7532 6916 7588
rect 6972 7084 7028 7140
rect 6860 6860 6916 6916
rect 6636 6748 6692 6804
rect 6748 6690 6804 6692
rect 6748 6638 6750 6690
rect 6750 6638 6802 6690
rect 6802 6638 6804 6690
rect 6748 6636 6804 6638
rect 6524 6524 6580 6580
rect 5628 6412 5684 6468
rect 5852 6076 5908 6132
rect 5628 5964 5684 6020
rect 5628 3554 5684 3556
rect 5628 3502 5630 3554
rect 5630 3502 5682 3554
rect 5682 3502 5684 3554
rect 5628 3500 5684 3502
rect 5740 5740 5796 5796
rect 5852 5068 5908 5124
rect 6076 6300 6132 6356
rect 6532 6298 6588 6300
rect 6532 6246 6534 6298
rect 6534 6246 6586 6298
rect 6586 6246 6588 6298
rect 6532 6244 6588 6246
rect 6636 6298 6692 6300
rect 6636 6246 6638 6298
rect 6638 6246 6690 6298
rect 6690 6246 6692 6298
rect 6636 6244 6692 6246
rect 6740 6298 6796 6300
rect 6740 6246 6742 6298
rect 6742 6246 6794 6298
rect 6794 6246 6796 6298
rect 6740 6244 6796 6246
rect 7420 7868 7476 7924
rect 7084 6076 7140 6132
rect 7196 6972 7252 7028
rect 6188 5516 6244 5572
rect 5964 3724 6020 3780
rect 6076 4396 6132 4452
rect 6300 3612 6356 3668
rect 6412 5740 6468 5796
rect 6524 5068 6580 5124
rect 7308 6578 7364 6580
rect 7308 6526 7310 6578
rect 7310 6526 7362 6578
rect 7362 6526 7364 6578
rect 7308 6524 7364 6526
rect 7420 6412 7476 6468
rect 6860 5906 6916 5908
rect 6860 5854 6862 5906
rect 6862 5854 6914 5906
rect 6914 5854 6916 5906
rect 6860 5852 6916 5854
rect 6860 5068 6916 5124
rect 6860 4844 6916 4900
rect 6532 4730 6588 4732
rect 6532 4678 6534 4730
rect 6534 4678 6586 4730
rect 6586 4678 6588 4730
rect 6532 4676 6588 4678
rect 6636 4730 6692 4732
rect 6636 4678 6638 4730
rect 6638 4678 6690 4730
rect 6690 4678 6692 4730
rect 6636 4676 6692 4678
rect 6740 4730 6796 4732
rect 6740 4678 6742 4730
rect 6742 4678 6794 4730
rect 6794 4678 6796 4730
rect 6740 4676 6796 4678
rect 6412 3500 6468 3556
rect 6412 3330 6468 3332
rect 6412 3278 6414 3330
rect 6414 3278 6466 3330
rect 6466 3278 6468 3330
rect 6412 3276 6468 3278
rect 6532 3162 6588 3164
rect 6532 3110 6534 3162
rect 6534 3110 6586 3162
rect 6586 3110 6588 3162
rect 6532 3108 6588 3110
rect 6636 3162 6692 3164
rect 6636 3110 6638 3162
rect 6638 3110 6690 3162
rect 6690 3110 6692 3162
rect 6636 3108 6692 3110
rect 6740 3162 6796 3164
rect 6740 3110 6742 3162
rect 6742 3110 6794 3162
rect 6794 3110 6796 3162
rect 6740 3108 6796 3110
rect 6972 4732 7028 4788
rect 7308 6076 7364 6132
rect 7084 4508 7140 4564
rect 7196 4172 7252 4228
rect 6972 3778 7028 3780
rect 6972 3726 6974 3778
rect 6974 3726 7026 3778
rect 7026 3726 7028 3778
rect 6972 3724 7028 3726
rect 7084 3666 7140 3668
rect 7084 3614 7086 3666
rect 7086 3614 7138 3666
rect 7138 3614 7140 3666
rect 7084 3612 7140 3614
rect 8204 8652 8260 8708
rect 7980 8146 8036 8148
rect 7980 8094 7982 8146
rect 7982 8094 8034 8146
rect 8034 8094 8036 8146
rect 7980 8092 8036 8094
rect 7868 7980 7924 8036
rect 7756 7308 7812 7364
rect 7980 6188 8036 6244
rect 7756 5068 7812 5124
rect 7980 5740 8036 5796
rect 8428 8876 8484 8932
rect 8316 8092 8372 8148
rect 8204 7644 8260 7700
rect 7980 4620 8036 4676
rect 7868 4508 7924 4564
rect 7980 3388 8036 3444
rect 8316 7420 8372 7476
rect 8428 7308 8484 7364
rect 8652 6860 8708 6916
rect 8876 8652 8932 8708
rect 8876 7308 8932 7364
rect 9772 9548 9828 9604
rect 9212 8988 9268 9044
rect 9192 8650 9248 8652
rect 9192 8598 9194 8650
rect 9194 8598 9246 8650
rect 9246 8598 9248 8650
rect 9192 8596 9248 8598
rect 9296 8650 9352 8652
rect 9296 8598 9298 8650
rect 9298 8598 9350 8650
rect 9350 8598 9352 8650
rect 9296 8596 9352 8598
rect 9400 8650 9456 8652
rect 9400 8598 9402 8650
rect 9402 8598 9454 8650
rect 9454 8598 9456 8650
rect 9400 8596 9456 8598
rect 9548 7586 9604 7588
rect 9548 7534 9550 7586
rect 9550 7534 9602 7586
rect 9602 7534 9604 7586
rect 9548 7532 9604 7534
rect 9192 7082 9248 7084
rect 9192 7030 9194 7082
rect 9194 7030 9246 7082
rect 9246 7030 9248 7082
rect 9192 7028 9248 7030
rect 9296 7082 9352 7084
rect 9296 7030 9298 7082
rect 9298 7030 9350 7082
rect 9350 7030 9352 7082
rect 9296 7028 9352 7030
rect 9400 7082 9456 7084
rect 9400 7030 9402 7082
rect 9402 7030 9454 7082
rect 9454 7030 9456 7082
rect 9400 7028 9456 7030
rect 9548 5906 9604 5908
rect 9548 5854 9550 5906
rect 9550 5854 9602 5906
rect 9602 5854 9604 5906
rect 9548 5852 9604 5854
rect 9192 5514 9248 5516
rect 9192 5462 9194 5514
rect 9194 5462 9246 5514
rect 9246 5462 9248 5514
rect 9192 5460 9248 5462
rect 9296 5514 9352 5516
rect 9296 5462 9298 5514
rect 9298 5462 9350 5514
rect 9350 5462 9352 5514
rect 9296 5460 9352 5462
rect 9400 5514 9456 5516
rect 9400 5462 9402 5514
rect 9402 5462 9454 5514
rect 9454 5462 9456 5514
rect 9400 5460 9456 5462
rect 9996 9100 10052 9156
rect 10108 8764 10164 8820
rect 9884 8258 9940 8260
rect 9884 8206 9886 8258
rect 9886 8206 9938 8258
rect 9938 8206 9940 8258
rect 9884 8204 9940 8206
rect 9884 5682 9940 5684
rect 9884 5630 9886 5682
rect 9886 5630 9938 5682
rect 9938 5630 9940 5682
rect 9884 5628 9940 5630
rect 9660 5292 9716 5348
rect 8988 4956 9044 5012
rect 8316 3388 8372 3444
rect 8652 3612 8708 3668
rect 8876 4396 8932 4452
rect 9192 3946 9248 3948
rect 9192 3894 9194 3946
rect 9194 3894 9246 3946
rect 9246 3894 9248 3946
rect 9192 3892 9248 3894
rect 9296 3946 9352 3948
rect 9296 3894 9298 3946
rect 9298 3894 9350 3946
rect 9350 3894 9352 3946
rect 9296 3892 9352 3894
rect 9400 3946 9456 3948
rect 9400 3894 9402 3946
rect 9402 3894 9454 3946
rect 9454 3894 9456 3946
rect 9400 3892 9456 3894
rect 9660 4562 9716 4564
rect 9660 4510 9662 4562
rect 9662 4510 9714 4562
rect 9714 4510 9716 4562
rect 9660 4508 9716 4510
rect 10444 8146 10500 8148
rect 10444 8094 10446 8146
rect 10446 8094 10498 8146
rect 10498 8094 10500 8146
rect 10444 8092 10500 8094
rect 10220 7532 10276 7588
rect 10108 6412 10164 6468
rect 9996 4172 10052 4228
rect 10332 6188 10388 6244
rect 9324 3276 9380 3332
rect 9884 3442 9940 3444
rect 9884 3390 9886 3442
rect 9886 3390 9938 3442
rect 9938 3390 9940 3442
rect 9884 3388 9940 3390
rect 10108 3388 10164 3444
rect 10668 6636 10724 6692
rect 10668 5628 10724 5684
rect 10556 4844 10612 4900
rect 10668 4172 10724 4228
rect 11228 9212 11284 9268
rect 11452 9548 11508 9604
rect 11228 7474 11284 7476
rect 11228 7422 11230 7474
rect 11230 7422 11282 7474
rect 11282 7422 11284 7474
rect 11228 7420 11284 7422
rect 11228 6748 11284 6804
rect 11116 5292 11172 5348
rect 11116 4844 11172 4900
rect 10892 4396 10948 4452
rect 12124 10498 12180 10500
rect 12124 10446 12126 10498
rect 12126 10446 12178 10498
rect 12178 10446 12180 10498
rect 12124 10444 12180 10446
rect 14512 10218 14568 10220
rect 14512 10166 14514 10218
rect 14514 10166 14566 10218
rect 14566 10166 14568 10218
rect 14512 10164 14568 10166
rect 14616 10218 14672 10220
rect 14616 10166 14618 10218
rect 14618 10166 14670 10218
rect 14670 10166 14672 10218
rect 14616 10164 14672 10166
rect 14720 10218 14776 10220
rect 14720 10166 14722 10218
rect 14722 10166 14774 10218
rect 14774 10166 14776 10218
rect 14720 10164 14776 10166
rect 11564 9042 11620 9044
rect 11564 8990 11566 9042
rect 11566 8990 11618 9042
rect 11618 8990 11620 9042
rect 11564 8988 11620 8990
rect 11852 9434 11908 9436
rect 11852 9382 11854 9434
rect 11854 9382 11906 9434
rect 11906 9382 11908 9434
rect 11852 9380 11908 9382
rect 11956 9434 12012 9436
rect 11956 9382 11958 9434
rect 11958 9382 12010 9434
rect 12010 9382 12012 9434
rect 11956 9380 12012 9382
rect 12060 9434 12116 9436
rect 12060 9382 12062 9434
rect 12062 9382 12114 9434
rect 12114 9382 12116 9434
rect 12060 9380 12116 9382
rect 12124 9154 12180 9156
rect 12124 9102 12126 9154
rect 12126 9102 12178 9154
rect 12178 9102 12180 9154
rect 12124 9100 12180 9102
rect 12684 9602 12740 9604
rect 12684 9550 12686 9602
rect 12686 9550 12738 9602
rect 12738 9550 12740 9602
rect 12684 9548 12740 9550
rect 12908 8876 12964 8932
rect 12236 8204 12292 8260
rect 12460 8204 12516 8260
rect 11852 7866 11908 7868
rect 11852 7814 11854 7866
rect 11854 7814 11906 7866
rect 11906 7814 11908 7866
rect 11852 7812 11908 7814
rect 11956 7866 12012 7868
rect 11956 7814 11958 7866
rect 11958 7814 12010 7866
rect 12010 7814 12012 7866
rect 11956 7812 12012 7814
rect 12060 7866 12116 7868
rect 12060 7814 12062 7866
rect 12062 7814 12114 7866
rect 12114 7814 12116 7866
rect 12060 7812 12116 7814
rect 12124 7586 12180 7588
rect 12124 7534 12126 7586
rect 12126 7534 12178 7586
rect 12178 7534 12180 7586
rect 12124 7532 12180 7534
rect 11852 6298 11908 6300
rect 11852 6246 11854 6298
rect 11854 6246 11906 6298
rect 11906 6246 11908 6298
rect 11852 6244 11908 6246
rect 11956 6298 12012 6300
rect 11956 6246 11958 6298
rect 11958 6246 12010 6298
rect 12010 6246 12012 6298
rect 11956 6244 12012 6246
rect 12060 6298 12116 6300
rect 12060 6246 12062 6298
rect 12062 6246 12114 6298
rect 12114 6246 12116 6298
rect 12060 6244 12116 6246
rect 12348 6690 12404 6692
rect 12348 6638 12350 6690
rect 12350 6638 12402 6690
rect 12402 6638 12404 6690
rect 12348 6636 12404 6638
rect 12236 6076 12292 6132
rect 11852 4730 11908 4732
rect 11852 4678 11854 4730
rect 11854 4678 11906 4730
rect 11906 4678 11908 4730
rect 11852 4676 11908 4678
rect 11956 4730 12012 4732
rect 11956 4678 11958 4730
rect 11958 4678 12010 4730
rect 12010 4678 12012 4730
rect 11956 4676 12012 4678
rect 12060 4730 12116 4732
rect 12060 4678 12062 4730
rect 12062 4678 12114 4730
rect 12114 4678 12116 4730
rect 12060 4676 12116 4678
rect 11788 4396 11844 4452
rect 11852 3162 11908 3164
rect 11852 3110 11854 3162
rect 11854 3110 11906 3162
rect 11906 3110 11908 3162
rect 11852 3108 11908 3110
rect 11956 3162 12012 3164
rect 11956 3110 11958 3162
rect 11958 3110 12010 3162
rect 12010 3110 12012 3162
rect 11956 3108 12012 3110
rect 12060 3162 12116 3164
rect 12060 3110 12062 3162
rect 12062 3110 12114 3162
rect 12114 3110 12116 3162
rect 12060 3108 12116 3110
rect 12796 6524 12852 6580
rect 13020 7420 13076 7476
rect 13356 7308 13412 7364
rect 12572 3612 12628 3668
rect 13244 5180 13300 5236
rect 12908 5010 12964 5012
rect 12908 4958 12910 5010
rect 12910 4958 12962 5010
rect 12962 4958 12964 5010
rect 12908 4956 12964 4958
rect 12796 4898 12852 4900
rect 12796 4846 12798 4898
rect 12798 4846 12850 4898
rect 12850 4846 12852 4898
rect 12796 4844 12852 4846
rect 13132 4732 13188 4788
rect 13020 4338 13076 4340
rect 13020 4286 13022 4338
rect 13022 4286 13074 4338
rect 13074 4286 13076 4338
rect 13020 4284 13076 4286
rect 12684 3500 12740 3556
rect 13468 6860 13524 6916
rect 13468 6690 13524 6692
rect 13468 6638 13470 6690
rect 13470 6638 13522 6690
rect 13522 6638 13524 6690
rect 13468 6636 13524 6638
rect 13356 4956 13412 5012
rect 13468 5740 13524 5796
rect 13692 7420 13748 7476
rect 14028 6748 14084 6804
rect 14140 7196 14196 7252
rect 14028 5964 14084 6020
rect 14028 5628 14084 5684
rect 13804 4956 13860 5012
rect 13468 4898 13524 4900
rect 13468 4846 13470 4898
rect 13470 4846 13522 4898
rect 13522 4846 13524 4898
rect 13468 4844 13524 4846
rect 13692 4898 13748 4900
rect 13692 4846 13694 4898
rect 13694 4846 13746 4898
rect 13746 4846 13748 4898
rect 13692 4844 13748 4846
rect 13692 4508 13748 4564
rect 14512 8650 14568 8652
rect 14512 8598 14514 8650
rect 14514 8598 14566 8650
rect 14566 8598 14568 8650
rect 14512 8596 14568 8598
rect 14616 8650 14672 8652
rect 14616 8598 14618 8650
rect 14618 8598 14670 8650
rect 14670 8598 14672 8650
rect 14616 8596 14672 8598
rect 14720 8650 14776 8652
rect 14720 8598 14722 8650
rect 14722 8598 14774 8650
rect 14774 8598 14776 8650
rect 14720 8596 14776 8598
rect 14512 7082 14568 7084
rect 14512 7030 14514 7082
rect 14514 7030 14566 7082
rect 14566 7030 14568 7082
rect 14512 7028 14568 7030
rect 14616 7082 14672 7084
rect 14616 7030 14618 7082
rect 14618 7030 14670 7082
rect 14670 7030 14672 7082
rect 14616 7028 14672 7030
rect 14720 7082 14776 7084
rect 14720 7030 14722 7082
rect 14722 7030 14774 7082
rect 14774 7030 14776 7082
rect 14720 7028 14776 7030
rect 14252 6076 14308 6132
rect 14924 5964 14980 6020
rect 14512 5514 14568 5516
rect 14512 5462 14514 5514
rect 14514 5462 14566 5514
rect 14566 5462 14568 5514
rect 14512 5460 14568 5462
rect 14616 5514 14672 5516
rect 14616 5462 14618 5514
rect 14618 5462 14670 5514
rect 14670 5462 14672 5514
rect 14616 5460 14672 5462
rect 14720 5514 14776 5516
rect 14720 5462 14722 5514
rect 14722 5462 14774 5514
rect 14774 5462 14776 5514
rect 14720 5460 14776 5462
rect 14140 4956 14196 5012
rect 15036 5292 15092 5348
rect 14252 4450 14308 4452
rect 14252 4398 14254 4450
rect 14254 4398 14306 4450
rect 14306 4398 14308 4450
rect 14252 4396 14308 4398
rect 14364 4284 14420 4340
rect 13916 4060 13972 4116
rect 13580 3612 13636 3668
rect 13020 3388 13076 3444
rect 13244 3330 13300 3332
rect 13244 3278 13246 3330
rect 13246 3278 13298 3330
rect 13298 3278 13300 3330
rect 13244 3276 13300 3278
rect 14512 3946 14568 3948
rect 14512 3894 14514 3946
rect 14514 3894 14566 3946
rect 14566 3894 14568 3946
rect 14512 3892 14568 3894
rect 14616 3946 14672 3948
rect 14616 3894 14618 3946
rect 14618 3894 14670 3946
rect 14670 3894 14672 3946
rect 14616 3892 14672 3894
rect 14720 3946 14776 3948
rect 14720 3894 14722 3946
rect 14722 3894 14774 3946
rect 14774 3894 14776 3946
rect 14720 3892 14776 3894
rect 15484 9548 15540 9604
rect 15148 4844 15204 4900
rect 15260 5852 15316 5908
rect 15148 3724 15204 3780
rect 15820 7362 15876 7364
rect 15820 7310 15822 7362
rect 15822 7310 15874 7362
rect 15874 7310 15876 7362
rect 15820 7308 15876 7310
rect 15596 6748 15652 6804
rect 17172 15706 17228 15708
rect 17172 15654 17174 15706
rect 17174 15654 17226 15706
rect 17226 15654 17228 15706
rect 17172 15652 17228 15654
rect 17276 15706 17332 15708
rect 17276 15654 17278 15706
rect 17278 15654 17330 15706
rect 17330 15654 17332 15706
rect 17276 15652 17332 15654
rect 17380 15706 17436 15708
rect 17380 15654 17382 15706
rect 17382 15654 17434 15706
rect 17434 15654 17436 15706
rect 17380 15652 17436 15654
rect 17172 14138 17228 14140
rect 17172 14086 17174 14138
rect 17174 14086 17226 14138
rect 17226 14086 17228 14138
rect 17172 14084 17228 14086
rect 17276 14138 17332 14140
rect 17276 14086 17278 14138
rect 17278 14086 17330 14138
rect 17330 14086 17332 14138
rect 17276 14084 17332 14086
rect 17380 14138 17436 14140
rect 17380 14086 17382 14138
rect 17382 14086 17434 14138
rect 17434 14086 17436 14138
rect 17380 14084 17436 14086
rect 17172 12570 17228 12572
rect 17172 12518 17174 12570
rect 17174 12518 17226 12570
rect 17226 12518 17228 12570
rect 17172 12516 17228 12518
rect 17276 12570 17332 12572
rect 17276 12518 17278 12570
rect 17278 12518 17330 12570
rect 17330 12518 17332 12570
rect 17276 12516 17332 12518
rect 17380 12570 17436 12572
rect 17380 12518 17382 12570
rect 17382 12518 17434 12570
rect 17434 12518 17436 12570
rect 17380 12516 17436 12518
rect 19832 14922 19888 14924
rect 19832 14870 19834 14922
rect 19834 14870 19886 14922
rect 19886 14870 19888 14922
rect 19832 14868 19888 14870
rect 19936 14922 19992 14924
rect 19936 14870 19938 14922
rect 19938 14870 19990 14922
rect 19990 14870 19992 14922
rect 19936 14868 19992 14870
rect 20040 14922 20096 14924
rect 20040 14870 20042 14922
rect 20042 14870 20094 14922
rect 20094 14870 20096 14922
rect 20040 14868 20096 14870
rect 19832 13354 19888 13356
rect 19832 13302 19834 13354
rect 19834 13302 19886 13354
rect 19886 13302 19888 13354
rect 19832 13300 19888 13302
rect 19936 13354 19992 13356
rect 19936 13302 19938 13354
rect 19938 13302 19990 13354
rect 19990 13302 19992 13354
rect 19936 13300 19992 13302
rect 20040 13354 20096 13356
rect 20040 13302 20042 13354
rect 20042 13302 20094 13354
rect 20094 13302 20096 13354
rect 20040 13300 20096 13302
rect 16380 11116 16436 11172
rect 17172 11002 17228 11004
rect 17172 10950 17174 11002
rect 17174 10950 17226 11002
rect 17226 10950 17228 11002
rect 17172 10948 17228 10950
rect 17276 11002 17332 11004
rect 17276 10950 17278 11002
rect 17278 10950 17330 11002
rect 17330 10950 17332 11002
rect 17276 10948 17332 10950
rect 17380 11002 17436 11004
rect 17380 10950 17382 11002
rect 17382 10950 17434 11002
rect 17434 10950 17436 11002
rect 17380 10948 17436 10950
rect 17172 9434 17228 9436
rect 17172 9382 17174 9434
rect 17174 9382 17226 9434
rect 17226 9382 17228 9434
rect 17172 9380 17228 9382
rect 17276 9434 17332 9436
rect 17276 9382 17278 9434
rect 17278 9382 17330 9434
rect 17330 9382 17332 9434
rect 17276 9380 17332 9382
rect 17380 9434 17436 9436
rect 17380 9382 17382 9434
rect 17382 9382 17434 9434
rect 17434 9382 17436 9434
rect 17380 9380 17436 9382
rect 16492 6860 16548 6916
rect 16716 7196 16772 7252
rect 15932 6524 15988 6580
rect 16716 6412 16772 6468
rect 16940 6748 16996 6804
rect 16492 5516 16548 5572
rect 16156 5068 16212 5124
rect 16380 5180 16436 5236
rect 16268 4956 16324 5012
rect 15484 4396 15540 4452
rect 15708 3388 15764 3444
rect 15932 3724 15988 3780
rect 16604 5404 16660 5460
rect 16716 5292 16772 5348
rect 16828 4284 16884 4340
rect 16828 3554 16884 3556
rect 16828 3502 16830 3554
rect 16830 3502 16882 3554
rect 16882 3502 16884 3554
rect 16828 3500 16884 3502
rect 17172 7866 17228 7868
rect 17172 7814 17174 7866
rect 17174 7814 17226 7866
rect 17226 7814 17228 7866
rect 17172 7812 17228 7814
rect 17276 7866 17332 7868
rect 17276 7814 17278 7866
rect 17278 7814 17330 7866
rect 17330 7814 17332 7866
rect 17276 7812 17332 7814
rect 17380 7866 17436 7868
rect 17380 7814 17382 7866
rect 17382 7814 17434 7866
rect 17434 7814 17436 7866
rect 17380 7812 17436 7814
rect 17500 7362 17556 7364
rect 17500 7310 17502 7362
rect 17502 7310 17554 7362
rect 17554 7310 17556 7362
rect 17500 7308 17556 7310
rect 17388 6636 17444 6692
rect 17276 6412 17332 6468
rect 19832 11786 19888 11788
rect 19832 11734 19834 11786
rect 19834 11734 19886 11786
rect 19886 11734 19888 11786
rect 19832 11732 19888 11734
rect 19936 11786 19992 11788
rect 19936 11734 19938 11786
rect 19938 11734 19990 11786
rect 19990 11734 19992 11786
rect 19936 11732 19992 11734
rect 20040 11786 20096 11788
rect 20040 11734 20042 11786
rect 20042 11734 20094 11786
rect 20094 11734 20096 11786
rect 20040 11732 20096 11734
rect 22492 15706 22548 15708
rect 22492 15654 22494 15706
rect 22494 15654 22546 15706
rect 22546 15654 22548 15706
rect 22492 15652 22548 15654
rect 22596 15706 22652 15708
rect 22596 15654 22598 15706
rect 22598 15654 22650 15706
rect 22650 15654 22652 15706
rect 22596 15652 22652 15654
rect 22700 15706 22756 15708
rect 22700 15654 22702 15706
rect 22702 15654 22754 15706
rect 22754 15654 22756 15706
rect 22700 15652 22756 15654
rect 22492 14138 22548 14140
rect 22492 14086 22494 14138
rect 22494 14086 22546 14138
rect 22546 14086 22548 14138
rect 22492 14084 22548 14086
rect 22596 14138 22652 14140
rect 22596 14086 22598 14138
rect 22598 14086 22650 14138
rect 22650 14086 22652 14138
rect 22596 14084 22652 14086
rect 22700 14138 22756 14140
rect 22700 14086 22702 14138
rect 22702 14086 22754 14138
rect 22754 14086 22756 14138
rect 22700 14084 22756 14086
rect 20300 11116 20356 11172
rect 21084 12684 21140 12740
rect 19832 10218 19888 10220
rect 19832 10166 19834 10218
rect 19834 10166 19886 10218
rect 19886 10166 19888 10218
rect 19832 10164 19888 10166
rect 19936 10218 19992 10220
rect 19936 10166 19938 10218
rect 19938 10166 19990 10218
rect 19990 10166 19992 10218
rect 19936 10164 19992 10166
rect 20040 10218 20096 10220
rect 20040 10166 20042 10218
rect 20042 10166 20094 10218
rect 20094 10166 20096 10218
rect 20040 10164 20096 10166
rect 17948 7420 18004 7476
rect 17172 6298 17228 6300
rect 17172 6246 17174 6298
rect 17174 6246 17226 6298
rect 17226 6246 17228 6298
rect 17172 6244 17228 6246
rect 17276 6298 17332 6300
rect 17276 6246 17278 6298
rect 17278 6246 17330 6298
rect 17330 6246 17332 6298
rect 17276 6244 17332 6246
rect 17380 6298 17436 6300
rect 17380 6246 17382 6298
rect 17382 6246 17434 6298
rect 17434 6246 17436 6298
rect 17380 6244 17436 6246
rect 17388 6130 17444 6132
rect 17388 6078 17390 6130
rect 17390 6078 17442 6130
rect 17442 6078 17444 6130
rect 17388 6076 17444 6078
rect 17612 6188 17668 6244
rect 17948 6188 18004 6244
rect 18172 6636 18228 6692
rect 17836 6018 17892 6020
rect 17836 5966 17838 6018
rect 17838 5966 17890 6018
rect 17890 5966 17892 6018
rect 17836 5964 17892 5966
rect 18060 5964 18116 6020
rect 17836 5740 17892 5796
rect 17500 5068 17556 5124
rect 17164 4956 17220 5012
rect 17172 4730 17228 4732
rect 17172 4678 17174 4730
rect 17174 4678 17226 4730
rect 17226 4678 17228 4730
rect 17172 4676 17228 4678
rect 17276 4730 17332 4732
rect 17276 4678 17278 4730
rect 17278 4678 17330 4730
rect 17330 4678 17332 4730
rect 17276 4676 17332 4678
rect 17380 4730 17436 4732
rect 17380 4678 17382 4730
rect 17382 4678 17434 4730
rect 17434 4678 17436 4730
rect 17380 4676 17436 4678
rect 16716 3388 16772 3444
rect 17500 4172 17556 4228
rect 17172 3162 17228 3164
rect 17172 3110 17174 3162
rect 17174 3110 17226 3162
rect 17226 3110 17228 3162
rect 17172 3108 17228 3110
rect 17276 3162 17332 3164
rect 17276 3110 17278 3162
rect 17278 3110 17330 3162
rect 17330 3110 17332 3162
rect 17276 3108 17332 3110
rect 17380 3162 17436 3164
rect 17380 3110 17382 3162
rect 17382 3110 17434 3162
rect 17434 3110 17436 3162
rect 17380 3108 17436 3110
rect 18060 5292 18116 5348
rect 18284 6524 18340 6580
rect 18284 5516 18340 5572
rect 18172 5068 18228 5124
rect 18396 5068 18452 5124
rect 18284 4844 18340 4900
rect 18396 4732 18452 4788
rect 18620 7084 18676 7140
rect 18508 4396 18564 4452
rect 18620 6860 18676 6916
rect 18956 7420 19012 7476
rect 18732 5404 18788 5460
rect 18844 6524 18900 6580
rect 18732 5180 18788 5236
rect 18732 3724 18788 3780
rect 19832 8650 19888 8652
rect 19832 8598 19834 8650
rect 19834 8598 19886 8650
rect 19886 8598 19888 8650
rect 19832 8596 19888 8598
rect 19936 8650 19992 8652
rect 19936 8598 19938 8650
rect 19938 8598 19990 8650
rect 19990 8598 19992 8650
rect 19936 8596 19992 8598
rect 20040 8650 20096 8652
rect 20040 8598 20042 8650
rect 20042 8598 20094 8650
rect 20094 8598 20096 8650
rect 20040 8596 20096 8598
rect 19180 6860 19236 6916
rect 20188 7532 20244 7588
rect 20076 7474 20132 7476
rect 20076 7422 20078 7474
rect 20078 7422 20130 7474
rect 20130 7422 20132 7474
rect 20076 7420 20132 7422
rect 19832 7082 19888 7084
rect 19832 7030 19834 7082
rect 19834 7030 19886 7082
rect 19886 7030 19888 7082
rect 19832 7028 19888 7030
rect 19936 7082 19992 7084
rect 19936 7030 19938 7082
rect 19938 7030 19990 7082
rect 19990 7030 19992 7082
rect 19936 7028 19992 7030
rect 20040 7082 20096 7084
rect 20040 7030 20042 7082
rect 20042 7030 20094 7082
rect 20094 7030 20096 7082
rect 20040 7028 20096 7030
rect 19740 6748 19796 6804
rect 19516 6076 19572 6132
rect 19964 5964 20020 6020
rect 19404 5852 19460 5908
rect 19292 5740 19348 5796
rect 19832 5514 19888 5516
rect 19292 5180 19348 5236
rect 19068 4396 19124 4452
rect 19404 5068 19460 5124
rect 19628 5404 19684 5460
rect 19832 5462 19834 5514
rect 19834 5462 19886 5514
rect 19886 5462 19888 5514
rect 19832 5460 19888 5462
rect 19936 5514 19992 5516
rect 19936 5462 19938 5514
rect 19938 5462 19990 5514
rect 19990 5462 19992 5514
rect 19936 5460 19992 5462
rect 20040 5514 20096 5516
rect 20040 5462 20042 5514
rect 20042 5462 20094 5514
rect 20094 5462 20096 5514
rect 20040 5460 20096 5462
rect 19740 5122 19796 5124
rect 19740 5070 19742 5122
rect 19742 5070 19794 5122
rect 19794 5070 19796 5122
rect 19740 5068 19796 5070
rect 19628 4956 19684 5012
rect 20188 4844 20244 4900
rect 20412 6860 20468 6916
rect 20412 6578 20468 6580
rect 20412 6526 20414 6578
rect 20414 6526 20466 6578
rect 20466 6526 20468 6578
rect 20412 6524 20468 6526
rect 20412 6076 20468 6132
rect 21868 12738 21924 12740
rect 21868 12686 21870 12738
rect 21870 12686 21922 12738
rect 21922 12686 21924 12738
rect 21868 12684 21924 12686
rect 21644 12348 21700 12404
rect 22492 12570 22548 12572
rect 22492 12518 22494 12570
rect 22494 12518 22546 12570
rect 22546 12518 22548 12570
rect 22492 12516 22548 12518
rect 22596 12570 22652 12572
rect 22596 12518 22598 12570
rect 22598 12518 22650 12570
rect 22650 12518 22652 12570
rect 22596 12516 22652 12518
rect 22700 12570 22756 12572
rect 22700 12518 22702 12570
rect 22702 12518 22754 12570
rect 22754 12518 22756 12570
rect 22700 12516 22756 12518
rect 22204 12348 22260 12404
rect 22492 11002 22548 11004
rect 22492 10950 22494 11002
rect 22494 10950 22546 11002
rect 22546 10950 22548 11002
rect 22492 10948 22548 10950
rect 22596 11002 22652 11004
rect 22596 10950 22598 11002
rect 22598 10950 22650 11002
rect 22650 10950 22652 11002
rect 22596 10948 22652 10950
rect 22700 11002 22756 11004
rect 22700 10950 22702 11002
rect 22702 10950 22754 11002
rect 22754 10950 22756 11002
rect 22700 10948 22756 10950
rect 22204 9602 22260 9604
rect 22204 9550 22206 9602
rect 22206 9550 22258 9602
rect 22258 9550 22260 9602
rect 22204 9548 22260 9550
rect 22492 9434 22548 9436
rect 22492 9382 22494 9434
rect 22494 9382 22546 9434
rect 22546 9382 22548 9434
rect 22492 9380 22548 9382
rect 22596 9434 22652 9436
rect 22596 9382 22598 9434
rect 22598 9382 22650 9434
rect 22650 9382 22652 9434
rect 22596 9380 22652 9382
rect 22700 9434 22756 9436
rect 22700 9382 22702 9434
rect 22702 9382 22754 9434
rect 22754 9382 22756 9434
rect 22700 9380 22756 9382
rect 20748 7420 20804 7476
rect 20748 7250 20804 7252
rect 20748 7198 20750 7250
rect 20750 7198 20802 7250
rect 20802 7198 20804 7250
rect 20748 7196 20804 7198
rect 20524 5740 20580 5796
rect 20636 6412 20692 6468
rect 20412 5292 20468 5348
rect 20300 4732 20356 4788
rect 20524 4508 20580 4564
rect 19832 3946 19888 3948
rect 19832 3894 19834 3946
rect 19834 3894 19886 3946
rect 19886 3894 19888 3946
rect 19832 3892 19888 3894
rect 19936 3946 19992 3948
rect 19936 3894 19938 3946
rect 19938 3894 19990 3946
rect 19990 3894 19992 3946
rect 19936 3892 19992 3894
rect 20040 3946 20096 3948
rect 20040 3894 20042 3946
rect 20042 3894 20094 3946
rect 20094 3894 20096 3946
rect 20040 3892 20096 3894
rect 20748 5068 20804 5124
rect 21196 6860 21252 6916
rect 20972 6412 21028 6468
rect 21532 7586 21588 7588
rect 21532 7534 21534 7586
rect 21534 7534 21586 7586
rect 21586 7534 21588 7586
rect 21532 7532 21588 7534
rect 21756 6860 21812 6916
rect 21420 5740 21476 5796
rect 21420 5234 21476 5236
rect 21420 5182 21422 5234
rect 21422 5182 21474 5234
rect 21474 5182 21476 5234
rect 21420 5180 21476 5182
rect 21308 5122 21364 5124
rect 21308 5070 21310 5122
rect 21310 5070 21362 5122
rect 21362 5070 21364 5122
rect 21308 5068 21364 5070
rect 21420 4284 21476 4340
rect 20972 3612 21028 3668
rect 20748 3442 20804 3444
rect 20748 3390 20750 3442
rect 20750 3390 20802 3442
rect 20802 3390 20804 3442
rect 20748 3388 20804 3390
rect 21532 3724 21588 3780
rect 21868 5628 21924 5684
rect 22492 7866 22548 7868
rect 22492 7814 22494 7866
rect 22494 7814 22546 7866
rect 22546 7814 22548 7866
rect 22492 7812 22548 7814
rect 22596 7866 22652 7868
rect 22596 7814 22598 7866
rect 22598 7814 22650 7866
rect 22650 7814 22652 7866
rect 22596 7812 22652 7814
rect 22700 7866 22756 7868
rect 22700 7814 22702 7866
rect 22702 7814 22754 7866
rect 22754 7814 22756 7866
rect 22700 7812 22756 7814
rect 22428 7420 22484 7476
rect 22092 6578 22148 6580
rect 22092 6526 22094 6578
rect 22094 6526 22146 6578
rect 22146 6526 22148 6578
rect 22092 6524 22148 6526
rect 21868 4508 21924 4564
rect 22492 6298 22548 6300
rect 22492 6246 22494 6298
rect 22494 6246 22546 6298
rect 22546 6246 22548 6298
rect 22492 6244 22548 6246
rect 22596 6298 22652 6300
rect 22596 6246 22598 6298
rect 22598 6246 22650 6298
rect 22650 6246 22652 6298
rect 22596 6244 22652 6246
rect 22700 6298 22756 6300
rect 22700 6246 22702 6298
rect 22702 6246 22754 6298
rect 22754 6246 22756 6298
rect 22700 6244 22756 6246
rect 22492 4730 22548 4732
rect 22492 4678 22494 4730
rect 22494 4678 22546 4730
rect 22546 4678 22548 4730
rect 22492 4676 22548 4678
rect 22596 4730 22652 4732
rect 22596 4678 22598 4730
rect 22598 4678 22650 4730
rect 22650 4678 22652 4730
rect 22596 4676 22652 4678
rect 22700 4730 22756 4732
rect 22700 4678 22702 4730
rect 22702 4678 22754 4730
rect 22754 4678 22756 4730
rect 22700 4676 22756 4678
rect 22492 3162 22548 3164
rect 22492 3110 22494 3162
rect 22494 3110 22546 3162
rect 22546 3110 22548 3162
rect 22492 3108 22548 3110
rect 22596 3162 22652 3164
rect 22596 3110 22598 3162
rect 22598 3110 22650 3162
rect 22650 3110 22652 3162
rect 22596 3108 22652 3110
rect 22700 3162 22756 3164
rect 22700 3110 22702 3162
rect 22702 3110 22754 3162
rect 22754 3110 22756 3162
rect 22700 3108 22756 3110
rect 22316 2492 22372 2548
<< metal3 >>
rect 0 17332 800 17360
rect 23200 17332 24000 17360
rect 0 17276 3500 17332
rect 3556 17276 3566 17332
rect 22194 17276 22204 17332
rect 22260 17276 24000 17332
rect 0 17248 800 17276
rect 23200 17248 24000 17276
rect 0 16884 800 16912
rect 0 16828 3612 16884
rect 3668 16828 3678 16884
rect 0 16800 800 16828
rect 0 16436 800 16464
rect 3862 16436 3872 16492
rect 3928 16436 3976 16492
rect 4032 16436 4080 16492
rect 4136 16436 4146 16492
rect 9182 16436 9192 16492
rect 9248 16436 9296 16492
rect 9352 16436 9400 16492
rect 9456 16436 9466 16492
rect 14502 16436 14512 16492
rect 14568 16436 14616 16492
rect 14672 16436 14720 16492
rect 14776 16436 14786 16492
rect 19822 16436 19832 16492
rect 19888 16436 19936 16492
rect 19992 16436 20040 16492
rect 20096 16436 20106 16492
rect 0 16380 3052 16436
rect 3108 16380 3118 16436
rect 0 16352 800 16380
rect 16146 16268 16156 16324
rect 16212 16268 17052 16324
rect 17108 16268 17118 16324
rect 0 15988 800 16016
rect 0 15932 2380 15988
rect 2436 15932 2446 15988
rect 0 15904 800 15932
rect 8754 15820 8764 15876
rect 8820 15820 9436 15876
rect 9492 15820 15932 15876
rect 15988 15820 15998 15876
rect 6522 15652 6532 15708
rect 6588 15652 6636 15708
rect 6692 15652 6740 15708
rect 6796 15652 6806 15708
rect 11842 15652 11852 15708
rect 11908 15652 11956 15708
rect 12012 15652 12060 15708
rect 12116 15652 12126 15708
rect 17162 15652 17172 15708
rect 17228 15652 17276 15708
rect 17332 15652 17380 15708
rect 17436 15652 17446 15708
rect 22482 15652 22492 15708
rect 22548 15652 22596 15708
rect 22652 15652 22700 15708
rect 22756 15652 22766 15708
rect 0 15540 800 15568
rect 0 15484 3388 15540
rect 3444 15484 3454 15540
rect 0 15456 800 15484
rect 0 15092 800 15120
rect 0 15036 2156 15092
rect 2212 15036 2222 15092
rect 0 15008 800 15036
rect 1698 14924 1708 14980
rect 1764 14924 1774 14980
rect 0 14644 800 14672
rect 1708 14644 1764 14924
rect 3862 14868 3872 14924
rect 3928 14868 3976 14924
rect 4032 14868 4080 14924
rect 4136 14868 4146 14924
rect 9182 14868 9192 14924
rect 9248 14868 9296 14924
rect 9352 14868 9400 14924
rect 9456 14868 9466 14924
rect 14502 14868 14512 14924
rect 14568 14868 14616 14924
rect 14672 14868 14720 14924
rect 14776 14868 14786 14924
rect 19822 14868 19832 14924
rect 19888 14868 19936 14924
rect 19992 14868 20040 14924
rect 20096 14868 20106 14924
rect 0 14588 1764 14644
rect 0 14560 800 14588
rect 2146 14252 2156 14308
rect 2212 14252 2222 14308
rect 0 14196 800 14224
rect 2156 14196 2212 14252
rect 0 14140 2212 14196
rect 0 14112 800 14140
rect 6522 14084 6532 14140
rect 6588 14084 6636 14140
rect 6692 14084 6740 14140
rect 6796 14084 6806 14140
rect 11842 14084 11852 14140
rect 11908 14084 11956 14140
rect 12012 14084 12060 14140
rect 12116 14084 12126 14140
rect 17162 14084 17172 14140
rect 17228 14084 17276 14140
rect 17332 14084 17380 14140
rect 17436 14084 17446 14140
rect 22482 14084 22492 14140
rect 22548 14084 22596 14140
rect 22652 14084 22700 14140
rect 22756 14084 22766 14140
rect 1698 14028 1708 14084
rect 1764 14028 1774 14084
rect 0 13748 800 13776
rect 1708 13748 1764 14028
rect 0 13692 1764 13748
rect 0 13664 800 13692
rect 0 13300 800 13328
rect 3862 13300 3872 13356
rect 3928 13300 3976 13356
rect 4032 13300 4080 13356
rect 4136 13300 4146 13356
rect 9182 13300 9192 13356
rect 9248 13300 9296 13356
rect 9352 13300 9400 13356
rect 9456 13300 9466 13356
rect 14502 13300 14512 13356
rect 14568 13300 14616 13356
rect 14672 13300 14720 13356
rect 14776 13300 14786 13356
rect 19822 13300 19832 13356
rect 19888 13300 19936 13356
rect 19992 13300 20040 13356
rect 20096 13300 20106 13356
rect 0 13244 1708 13300
rect 1764 13244 1774 13300
rect 0 13216 800 13244
rect 0 12852 800 12880
rect 0 12796 1708 12852
rect 1764 12796 1774 12852
rect 0 12768 800 12796
rect 2146 12684 2156 12740
rect 2212 12684 2222 12740
rect 21074 12684 21084 12740
rect 21140 12684 21868 12740
rect 21924 12684 21934 12740
rect 0 12404 800 12432
rect 2156 12404 2212 12684
rect 6522 12516 6532 12572
rect 6588 12516 6636 12572
rect 6692 12516 6740 12572
rect 6796 12516 6806 12572
rect 11842 12516 11852 12572
rect 11908 12516 11956 12572
rect 12012 12516 12060 12572
rect 12116 12516 12126 12572
rect 17162 12516 17172 12572
rect 17228 12516 17276 12572
rect 17332 12516 17380 12572
rect 17436 12516 17446 12572
rect 22482 12516 22492 12572
rect 22548 12516 22596 12572
rect 22652 12516 22700 12572
rect 22756 12516 22766 12572
rect 23200 12404 24000 12432
rect 0 12348 2212 12404
rect 21634 12348 21644 12404
rect 21700 12348 22204 12404
rect 22260 12348 24000 12404
rect 0 12320 800 12348
rect 23200 12320 24000 12348
rect 3686 12012 3724 12068
rect 3780 12012 3790 12068
rect 0 11956 800 11984
rect 0 11900 1708 11956
rect 1764 11900 1774 11956
rect 0 11872 800 11900
rect 3862 11732 3872 11788
rect 3928 11732 3976 11788
rect 4032 11732 4080 11788
rect 4136 11732 4146 11788
rect 9182 11732 9192 11788
rect 9248 11732 9296 11788
rect 9352 11732 9400 11788
rect 9456 11732 9466 11788
rect 14502 11732 14512 11788
rect 14568 11732 14616 11788
rect 14672 11732 14720 11788
rect 14776 11732 14786 11788
rect 19822 11732 19832 11788
rect 19888 11732 19936 11788
rect 19992 11732 20040 11788
rect 20096 11732 20106 11788
rect 0 11508 800 11536
rect 0 11452 2156 11508
rect 2212 11452 2222 11508
rect 4834 11452 4844 11508
rect 4900 11452 4956 11508
rect 5012 11452 5022 11508
rect 0 11424 800 11452
rect 1698 11116 1708 11172
rect 1764 11116 1774 11172
rect 2454 11116 2492 11172
rect 2548 11116 2558 11172
rect 3378 11116 3388 11172
rect 3444 11116 3482 11172
rect 9986 11116 9996 11172
rect 10052 11116 15148 11172
rect 15204 11116 16380 11172
rect 16436 11116 20300 11172
rect 20356 11116 20366 11172
rect 0 11060 800 11088
rect 1708 11060 1764 11116
rect 0 11004 1764 11060
rect 0 10976 800 11004
rect 6522 10948 6532 11004
rect 6588 10948 6636 11004
rect 6692 10948 6740 11004
rect 6796 10948 6806 11004
rect 11842 10948 11852 11004
rect 11908 10948 11956 11004
rect 12012 10948 12060 11004
rect 12116 10948 12126 11004
rect 17162 10948 17172 11004
rect 17228 10948 17276 11004
rect 17332 10948 17380 11004
rect 17436 10948 17446 11004
rect 22482 10948 22492 11004
rect 22548 10948 22596 11004
rect 22652 10948 22700 11004
rect 22756 10948 22766 11004
rect 4470 10892 4508 10948
rect 4564 10892 4574 10948
rect 0 10612 800 10640
rect 0 10556 2044 10612
rect 2100 10556 2110 10612
rect 2370 10556 2380 10612
rect 2436 10556 3724 10612
rect 3780 10556 3790 10612
rect 0 10528 800 10556
rect 12114 10444 12124 10500
rect 12180 10444 12460 10500
rect 12516 10444 12526 10500
rect 0 10164 800 10192
rect 3862 10164 3872 10220
rect 3928 10164 3976 10220
rect 4032 10164 4080 10220
rect 4136 10164 4146 10220
rect 9182 10164 9192 10220
rect 9248 10164 9296 10220
rect 9352 10164 9400 10220
rect 9456 10164 9466 10220
rect 14502 10164 14512 10220
rect 14568 10164 14616 10220
rect 14672 10164 14720 10220
rect 14776 10164 14786 10220
rect 19822 10164 19832 10220
rect 19888 10164 19936 10220
rect 19992 10164 20040 10220
rect 20096 10164 20106 10220
rect 0 10108 1708 10164
rect 1764 10108 1774 10164
rect 0 10080 800 10108
rect 0 9716 800 9744
rect 0 9660 1764 9716
rect 0 9632 800 9660
rect 1708 9604 1764 9660
rect 1698 9548 1708 9604
rect 1764 9548 1774 9604
rect 2034 9548 2044 9604
rect 2100 9548 4172 9604
rect 4228 9548 4238 9604
rect 4834 9548 4844 9604
rect 4900 9548 5068 9604
rect 5124 9548 5134 9604
rect 7382 9548 7420 9604
rect 7476 9548 7486 9604
rect 8418 9548 8428 9604
rect 8484 9548 9772 9604
rect 9828 9548 9838 9604
rect 11442 9548 11452 9604
rect 11508 9548 12684 9604
rect 12740 9548 12750 9604
rect 15474 9548 15484 9604
rect 15540 9548 22204 9604
rect 22260 9548 22270 9604
rect 6522 9380 6532 9436
rect 6588 9380 6636 9436
rect 6692 9380 6740 9436
rect 6796 9380 6806 9436
rect 11842 9380 11852 9436
rect 11908 9380 11956 9436
rect 12012 9380 12060 9436
rect 12116 9380 12126 9436
rect 17162 9380 17172 9436
rect 17228 9380 17276 9436
rect 17332 9380 17380 9436
rect 17436 9380 17446 9436
rect 22482 9380 22492 9436
rect 22548 9380 22596 9436
rect 22652 9380 22700 9436
rect 22756 9380 22766 9436
rect 1810 9324 1820 9380
rect 1876 9324 2716 9380
rect 2772 9324 2782 9380
rect 3378 9324 3388 9380
rect 3444 9324 4396 9380
rect 4452 9324 5964 9380
rect 6020 9324 6030 9380
rect 0 9268 800 9296
rect 0 9212 2156 9268
rect 2212 9212 2222 9268
rect 2380 9212 5124 9268
rect 5282 9212 5292 9268
rect 5348 9212 11228 9268
rect 11284 9212 11294 9268
rect 0 9184 800 9212
rect 2380 9156 2436 9212
rect 2034 9100 2044 9156
rect 2100 9100 2436 9156
rect 2678 9100 2716 9156
rect 2772 9100 2782 9156
rect 3266 9100 3276 9156
rect 3332 9100 4844 9156
rect 4900 9100 4910 9156
rect 5068 9044 5124 9212
rect 6066 9100 6076 9156
rect 6132 9100 7084 9156
rect 7140 9100 7150 9156
rect 9986 9100 9996 9156
rect 10052 9100 12124 9156
rect 12180 9100 12190 9156
rect 5068 8988 9044 9044
rect 9202 8988 9212 9044
rect 9268 8988 11564 9044
rect 11620 8988 11630 9044
rect 8988 8932 9044 8988
rect 4946 8876 4956 8932
rect 5012 8876 5852 8932
rect 5908 8876 5918 8932
rect 7074 8876 7084 8932
rect 7140 8876 8428 8932
rect 8484 8876 8494 8932
rect 8988 8876 12908 8932
rect 12964 8876 12974 8932
rect 0 8820 800 8848
rect 0 8764 2492 8820
rect 2548 8764 2558 8820
rect 5366 8764 5404 8820
rect 5460 8764 5470 8820
rect 6178 8764 6188 8820
rect 6244 8764 6860 8820
rect 6916 8764 6926 8820
rect 7084 8764 10108 8820
rect 10164 8764 10174 8820
rect 0 8736 800 8764
rect 7084 8708 7140 8764
rect 4610 8652 4620 8708
rect 4676 8652 7140 8708
rect 8194 8652 8204 8708
rect 8260 8652 8876 8708
rect 8932 8652 8942 8708
rect 3862 8596 3872 8652
rect 3928 8596 3976 8652
rect 4032 8596 4080 8652
rect 4136 8596 4146 8652
rect 9182 8596 9192 8652
rect 9248 8596 9296 8652
rect 9352 8596 9400 8652
rect 9456 8596 9466 8652
rect 14502 8596 14512 8652
rect 14568 8596 14616 8652
rect 14672 8596 14720 8652
rect 14776 8596 14786 8652
rect 19822 8596 19832 8652
rect 19888 8596 19936 8652
rect 19992 8596 20040 8652
rect 20096 8596 20106 8652
rect 1922 8540 1932 8596
rect 1988 8540 2268 8596
rect 2324 8540 2334 8596
rect 6626 8540 6636 8596
rect 6692 8540 8316 8596
rect 8372 8540 8382 8596
rect 1810 8428 1820 8484
rect 1876 8428 1886 8484
rect 2566 8428 2604 8484
rect 2660 8428 2670 8484
rect 2930 8428 2940 8484
rect 2996 8428 3006 8484
rect 4834 8428 4844 8484
rect 4900 8428 4910 8484
rect 0 8372 800 8400
rect 1820 8372 1876 8428
rect 0 8316 1876 8372
rect 0 8288 800 8316
rect 2940 8148 2996 8428
rect 4844 8372 4900 8428
rect 4844 8316 5404 8372
rect 5460 8316 5470 8372
rect 6290 8316 6300 8372
rect 6356 8316 6972 8372
rect 7028 8316 7038 8372
rect 5954 8204 5964 8260
rect 6020 8204 9884 8260
rect 9940 8204 9950 8260
rect 12198 8204 12236 8260
rect 12292 8204 12302 8260
rect 12422 8204 12460 8260
rect 12516 8204 12526 8260
rect 1484 8092 2996 8148
rect 3490 8092 3500 8148
rect 3556 8092 3612 8148
rect 3668 8092 3678 8148
rect 4834 8092 4844 8148
rect 4900 8092 5516 8148
rect 5572 8092 5582 8148
rect 5730 8092 5740 8148
rect 5796 8092 5834 8148
rect 6626 8092 6636 8148
rect 6692 8092 7980 8148
rect 8036 8092 8046 8148
rect 8306 8092 8316 8148
rect 8372 8092 10444 8148
rect 10500 8092 10510 8148
rect 0 7924 800 7952
rect 1484 7924 1540 8092
rect 2706 7980 2716 8036
rect 2772 7980 3388 8036
rect 3444 7980 3454 8036
rect 3602 7980 3612 8036
rect 3668 7980 3724 8036
rect 3780 7980 3790 8036
rect 4050 7980 4060 8036
rect 4116 7980 7868 8036
rect 7924 7980 7934 8036
rect 0 7868 1540 7924
rect 1782 7868 1820 7924
rect 1876 7868 1886 7924
rect 2930 7868 2940 7924
rect 2996 7868 5068 7924
rect 5124 7868 5134 7924
rect 7382 7868 7420 7924
rect 7476 7868 7486 7924
rect 0 7840 800 7868
rect 6522 7812 6532 7868
rect 6588 7812 6636 7868
rect 6692 7812 6740 7868
rect 6796 7812 6806 7868
rect 11842 7812 11852 7868
rect 11908 7812 11956 7868
rect 12012 7812 12060 7868
rect 12116 7812 12126 7868
rect 17162 7812 17172 7868
rect 17228 7812 17276 7868
rect 17332 7812 17380 7868
rect 17436 7812 17446 7868
rect 22482 7812 22492 7868
rect 22548 7812 22596 7868
rect 22652 7812 22700 7868
rect 22756 7812 22766 7868
rect 2342 7756 2380 7812
rect 2436 7756 2446 7812
rect 3332 7756 5460 7812
rect 6290 7756 6300 7812
rect 6356 7756 6366 7812
rect 3332 7700 3388 7756
rect 5404 7700 5460 7756
rect 6300 7700 6356 7756
rect 1810 7644 1820 7700
rect 1876 7644 2604 7700
rect 2660 7644 2670 7700
rect 3042 7644 3052 7700
rect 3108 7644 3388 7700
rect 3490 7644 3500 7700
rect 3556 7644 3566 7700
rect 5394 7644 5404 7700
rect 5460 7644 5470 7700
rect 6300 7644 8204 7700
rect 8260 7644 8270 7700
rect 1698 7532 1708 7588
rect 1764 7532 2492 7588
rect 2548 7532 2558 7588
rect 0 7476 800 7504
rect 3500 7476 3556 7644
rect 3714 7532 3724 7588
rect 3780 7532 6076 7588
rect 6132 7532 6142 7588
rect 6850 7532 6860 7588
rect 6916 7532 9548 7588
rect 9604 7532 9614 7588
rect 10210 7532 10220 7588
rect 10276 7532 12124 7588
rect 12180 7532 12190 7588
rect 20178 7532 20188 7588
rect 20244 7532 21532 7588
rect 21588 7532 21598 7588
rect 10220 7476 10276 7532
rect 23200 7476 24000 7504
rect 0 7420 3556 7476
rect 3826 7420 3836 7476
rect 3892 7420 5180 7476
rect 5236 7420 8036 7476
rect 8306 7420 8316 7476
rect 8372 7420 10276 7476
rect 11218 7420 11228 7476
rect 11284 7420 13020 7476
rect 13076 7420 13086 7476
rect 13654 7420 13692 7476
rect 13748 7420 17948 7476
rect 18004 7420 18014 7476
rect 18946 7420 18956 7476
rect 19012 7420 20076 7476
rect 20132 7420 20748 7476
rect 20804 7420 20814 7476
rect 22418 7420 22428 7476
rect 22484 7420 24000 7476
rect 0 7392 800 7420
rect 7980 7364 8036 7420
rect 23200 7392 24000 7420
rect 2146 7308 2156 7364
rect 2212 7308 7756 7364
rect 7812 7308 7822 7364
rect 7980 7308 8428 7364
rect 8484 7308 8494 7364
rect 8866 7308 8876 7364
rect 8932 7308 13356 7364
rect 13412 7308 13422 7364
rect 15810 7308 15820 7364
rect 15876 7308 17500 7364
rect 17556 7308 17566 7364
rect 3490 7196 3500 7252
rect 3556 7196 3724 7252
rect 3780 7196 3790 7252
rect 5058 7196 5068 7252
rect 5124 7196 14140 7252
rect 14196 7196 14206 7252
rect 16706 7196 16716 7252
rect 16772 7196 20748 7252
rect 20804 7196 20814 7252
rect 3378 7084 3388 7140
rect 3444 7084 3482 7140
rect 4694 7084 4732 7140
rect 4788 7084 4798 7140
rect 5170 7084 5180 7140
rect 5236 7084 6188 7140
rect 6244 7084 6972 7140
rect 7028 7084 7038 7140
rect 18582 7084 18620 7140
rect 18676 7084 18686 7140
rect 0 7028 800 7056
rect 3862 7028 3872 7084
rect 3928 7028 3976 7084
rect 4032 7028 4080 7084
rect 4136 7028 4146 7084
rect 9182 7028 9192 7084
rect 9248 7028 9296 7084
rect 9352 7028 9400 7084
rect 9456 7028 9466 7084
rect 14502 7028 14512 7084
rect 14568 7028 14616 7084
rect 14672 7028 14720 7084
rect 14776 7028 14786 7084
rect 19822 7028 19832 7084
rect 19888 7028 19936 7084
rect 19992 7028 20040 7084
rect 20096 7028 20106 7084
rect 0 6972 2044 7028
rect 2100 6972 2110 7028
rect 4274 6972 4284 7028
rect 4340 6972 7196 7028
rect 7252 6972 7262 7028
rect 0 6944 800 6972
rect 5058 6860 5068 6916
rect 5124 6860 5628 6916
rect 5684 6860 5694 6916
rect 6066 6860 6076 6916
rect 6132 6860 6860 6916
rect 6916 6860 6926 6916
rect 8642 6860 8652 6916
rect 8708 6860 13468 6916
rect 13524 6860 16492 6916
rect 16548 6860 16558 6916
rect 18610 6860 18620 6916
rect 18676 6860 19180 6916
rect 19236 6860 19246 6916
rect 20402 6860 20412 6916
rect 20468 6860 21196 6916
rect 21252 6860 21262 6916
rect 21746 6860 21756 6916
rect 21812 6860 21822 6916
rect 6150 6748 6188 6804
rect 6244 6748 6254 6804
rect 6626 6748 6636 6804
rect 6692 6748 11228 6804
rect 11284 6748 11294 6804
rect 14018 6748 14028 6804
rect 14084 6748 15596 6804
rect 15652 6748 15662 6804
rect 16930 6748 16940 6804
rect 16996 6748 19740 6804
rect 19796 6748 19806 6804
rect 21756 6692 21812 6860
rect 3490 6636 3500 6692
rect 3556 6636 4620 6692
rect 4676 6636 4686 6692
rect 4834 6636 4844 6692
rect 4900 6636 5180 6692
rect 5236 6636 5246 6692
rect 5404 6636 6748 6692
rect 6804 6636 7420 6692
rect 7476 6636 10668 6692
rect 10724 6636 10734 6692
rect 12338 6636 12348 6692
rect 12404 6636 13468 6692
rect 13524 6636 13534 6692
rect 15092 6636 17388 6692
rect 17444 6636 17454 6692
rect 18162 6636 18172 6692
rect 18228 6636 21812 6692
rect 0 6580 800 6608
rect 0 6524 4620 6580
rect 4676 6524 4686 6580
rect 0 6496 800 6524
rect 5404 6468 5460 6636
rect 15092 6580 15148 6636
rect 5618 6524 5628 6580
rect 5684 6524 6524 6580
rect 6580 6524 7308 6580
rect 7364 6524 7374 6580
rect 12786 6524 12796 6580
rect 12852 6524 15148 6580
rect 15922 6524 15932 6580
rect 15988 6524 18284 6580
rect 18340 6524 18350 6580
rect 18834 6524 18844 6580
rect 18900 6524 20412 6580
rect 20468 6524 22092 6580
rect 22148 6524 22158 6580
rect 1922 6412 1932 6468
rect 1988 6412 1998 6468
rect 4274 6412 4284 6468
rect 4340 6412 5460 6468
rect 5618 6412 5628 6468
rect 5684 6412 7420 6468
rect 7476 6412 7486 6468
rect 10098 6412 10108 6468
rect 10164 6412 16716 6468
rect 16772 6412 16782 6468
rect 16940 6412 17276 6468
rect 17332 6412 17342 6468
rect 20626 6412 20636 6468
rect 20692 6412 20972 6468
rect 21028 6412 21038 6468
rect 0 6132 800 6160
rect 0 6076 1708 6132
rect 1764 6076 1774 6132
rect 0 6048 800 6076
rect 0 5684 800 5712
rect 1932 5684 1988 6412
rect 2818 6300 2828 6356
rect 2884 6300 6076 6356
rect 6132 6300 6142 6356
rect 6522 6244 6532 6300
rect 6588 6244 6636 6300
rect 6692 6244 6740 6300
rect 6796 6244 6806 6300
rect 11842 6244 11852 6300
rect 11908 6244 11956 6300
rect 12012 6244 12060 6300
rect 12116 6244 12126 6300
rect 5394 6188 5404 6244
rect 5460 6188 6300 6244
rect 6356 6188 6366 6244
rect 7970 6188 7980 6244
rect 8036 6188 10332 6244
rect 10388 6188 10398 6244
rect 5404 6132 5460 6188
rect 16940 6132 16996 6412
rect 17162 6244 17172 6300
rect 17228 6244 17276 6300
rect 17332 6244 17380 6300
rect 17436 6244 17446 6300
rect 22482 6244 22492 6300
rect 22548 6244 22596 6300
rect 22652 6244 22700 6300
rect 22756 6244 22766 6300
rect 17602 6188 17612 6244
rect 17668 6188 17948 6244
rect 18004 6188 18014 6244
rect 2258 6076 2268 6132
rect 2324 6076 2940 6132
rect 2996 6076 3006 6132
rect 3332 6076 5460 6132
rect 5842 6076 5852 6132
rect 5908 6076 7084 6132
rect 7140 6076 7150 6132
rect 7298 6076 7308 6132
rect 7364 6076 12236 6132
rect 12292 6076 12302 6132
rect 13468 6076 14252 6132
rect 14308 6076 17388 6132
rect 17444 6076 17454 6132
rect 17836 6076 19516 6132
rect 19572 6076 20412 6132
rect 20468 6076 20478 6132
rect 3266 5852 3276 5908
rect 3332 5852 3388 6076
rect 3602 5964 3612 6020
rect 3668 5964 4732 6020
rect 4788 5964 5628 6020
rect 5684 5964 9604 6020
rect 9548 5908 9604 5964
rect 4162 5852 4172 5908
rect 4228 5852 6860 5908
rect 6916 5852 6926 5908
rect 9538 5852 9548 5908
rect 9604 5852 9614 5908
rect 13468 5796 13524 6076
rect 17836 6020 17892 6076
rect 14018 5964 14028 6020
rect 14084 5964 14924 6020
rect 14980 5964 17836 6020
rect 17892 5964 17902 6020
rect 18050 5964 18060 6020
rect 18116 5964 19964 6020
rect 20020 5964 20030 6020
rect 15250 5852 15260 5908
rect 15316 5852 19404 5908
rect 19460 5852 19628 5908
rect 19684 5852 19694 5908
rect 2146 5740 2156 5796
rect 2212 5740 3388 5796
rect 3938 5740 3948 5796
rect 4004 5740 4508 5796
rect 4564 5740 4956 5796
rect 5012 5740 5022 5796
rect 5394 5740 5404 5796
rect 5460 5740 5740 5796
rect 5796 5740 5806 5796
rect 6290 5740 6300 5796
rect 6356 5740 6412 5796
rect 6468 5740 6478 5796
rect 7970 5740 7980 5796
rect 8036 5740 8046 5796
rect 13458 5740 13468 5796
rect 13524 5740 13534 5796
rect 17826 5740 17836 5796
rect 17892 5740 19292 5796
rect 19348 5740 19358 5796
rect 20514 5740 20524 5796
rect 20580 5740 21420 5796
rect 21476 5740 21486 5796
rect 0 5628 1988 5684
rect 3332 5684 3388 5740
rect 7980 5684 8036 5740
rect 3332 5628 4284 5684
rect 4340 5628 8036 5684
rect 8092 5628 9884 5684
rect 9940 5628 9950 5684
rect 10658 5628 10668 5684
rect 10724 5628 14028 5684
rect 14084 5628 14094 5684
rect 14252 5628 21868 5684
rect 21924 5628 21934 5684
rect 0 5600 800 5628
rect 3266 5516 3276 5572
rect 3332 5516 3724 5572
rect 3780 5516 3790 5572
rect 4498 5516 4508 5572
rect 4564 5516 4732 5572
rect 4788 5516 4798 5572
rect 5058 5516 5068 5572
rect 5124 5516 6188 5572
rect 6244 5516 6254 5572
rect 3862 5460 3872 5516
rect 3928 5460 3976 5516
rect 4032 5460 4080 5516
rect 4136 5460 4146 5516
rect 4732 5460 4788 5516
rect 8092 5460 8148 5628
rect 9182 5460 9192 5516
rect 9248 5460 9296 5516
rect 9352 5460 9400 5516
rect 9456 5460 9466 5516
rect 4732 5404 8148 5460
rect 1922 5292 1932 5348
rect 1988 5292 9660 5348
rect 9716 5292 11116 5348
rect 11172 5292 11182 5348
rect 0 5236 800 5264
rect 0 5180 2716 5236
rect 2772 5180 2782 5236
rect 3938 5180 3948 5236
rect 4004 5180 4844 5236
rect 4900 5180 4910 5236
rect 5170 5180 5180 5236
rect 5236 5180 13244 5236
rect 13300 5180 13310 5236
rect 0 5152 800 5180
rect 14252 5124 14308 5628
rect 16482 5516 16492 5572
rect 16548 5516 18284 5572
rect 18340 5516 18350 5572
rect 14502 5460 14512 5516
rect 14568 5460 14616 5516
rect 14672 5460 14720 5516
rect 14776 5460 14786 5516
rect 19822 5460 19832 5516
rect 19888 5460 19936 5516
rect 19992 5460 20040 5516
rect 20096 5460 20106 5516
rect 16594 5404 16604 5460
rect 16660 5404 18732 5460
rect 18788 5404 19628 5460
rect 19684 5404 19694 5460
rect 15026 5292 15036 5348
rect 15092 5292 16716 5348
rect 16772 5292 16782 5348
rect 18050 5292 18060 5348
rect 18116 5292 20412 5348
rect 20468 5292 20478 5348
rect 16370 5180 16380 5236
rect 16436 5180 18732 5236
rect 18788 5180 18798 5236
rect 19282 5180 19292 5236
rect 19348 5180 21420 5236
rect 21476 5180 21486 5236
rect 2706 5068 2716 5124
rect 2772 5068 5852 5124
rect 5908 5068 5918 5124
rect 6076 5068 6524 5124
rect 6580 5068 6590 5124
rect 6850 5068 6860 5124
rect 6916 5068 7756 5124
rect 7812 5068 7822 5124
rect 8306 5068 8316 5124
rect 8372 5068 14308 5124
rect 16146 5068 16156 5124
rect 16212 5068 16884 5124
rect 17490 5068 17500 5124
rect 17556 5068 18172 5124
rect 18228 5068 18238 5124
rect 18386 5068 18396 5124
rect 18452 5068 19404 5124
rect 19460 5068 19470 5124
rect 19618 5068 19628 5124
rect 19684 5068 19740 5124
rect 19796 5068 19806 5124
rect 20738 5068 20748 5124
rect 20804 5068 21308 5124
rect 21364 5068 21374 5124
rect 6076 5012 6132 5068
rect 16828 5012 16884 5068
rect 4834 4956 4844 5012
rect 4900 4956 6132 5012
rect 8978 4956 8988 5012
rect 9044 4956 12236 5012
rect 12292 4956 12302 5012
rect 12898 4956 12908 5012
rect 12964 4956 13356 5012
rect 13412 4956 13804 5012
rect 13860 4956 13870 5012
rect 14130 4956 14140 5012
rect 14196 4956 16268 5012
rect 16324 4956 16334 5012
rect 16828 4956 17164 5012
rect 17220 4956 19628 5012
rect 19684 4956 19694 5012
rect 1810 4844 1820 4900
rect 1876 4844 3388 4900
rect 4162 4844 4172 4900
rect 4228 4844 4732 4900
rect 4788 4844 4798 4900
rect 4946 4844 4956 4900
rect 5012 4844 6860 4900
rect 6916 4844 6926 4900
rect 10546 4844 10556 4900
rect 10612 4844 10622 4900
rect 11106 4844 11116 4900
rect 11172 4844 12628 4900
rect 12786 4844 12796 4900
rect 12852 4844 13468 4900
rect 13524 4844 13534 4900
rect 13682 4844 13692 4900
rect 13748 4844 15148 4900
rect 15204 4844 15214 4900
rect 18274 4844 18284 4900
rect 18340 4844 20188 4900
rect 20244 4844 20254 4900
rect 0 4788 800 4816
rect 3332 4788 3388 4844
rect 10556 4788 10612 4844
rect 0 4732 1820 4788
rect 1876 4732 1886 4788
rect 3332 4732 5460 4788
rect 6962 4732 6972 4788
rect 7028 4732 10612 4788
rect 12572 4788 12628 4844
rect 12572 4732 13132 4788
rect 13188 4732 13198 4788
rect 18386 4732 18396 4788
rect 18452 4732 20300 4788
rect 20356 4732 20366 4788
rect 0 4704 800 4732
rect 5404 4676 5460 4732
rect 6522 4676 6532 4732
rect 6588 4676 6636 4732
rect 6692 4676 6740 4732
rect 6796 4676 6806 4732
rect 11842 4676 11852 4732
rect 11908 4676 11956 4732
rect 12012 4676 12060 4732
rect 12116 4676 12126 4732
rect 17162 4676 17172 4732
rect 17228 4676 17276 4732
rect 17332 4676 17380 4732
rect 17436 4676 17446 4732
rect 22482 4676 22492 4732
rect 22548 4676 22596 4732
rect 22652 4676 22700 4732
rect 22756 4676 22766 4732
rect 2594 4620 2604 4676
rect 2660 4620 3388 4676
rect 5394 4620 5404 4676
rect 5460 4620 5470 4676
rect 7970 4620 7980 4676
rect 8036 4620 8316 4676
rect 8372 4620 8382 4676
rect 3332 4564 3388 4620
rect 1474 4508 1484 4564
rect 1540 4508 1550 4564
rect 3332 4508 6132 4564
rect 7074 4508 7084 4564
rect 7140 4508 7868 4564
rect 7924 4508 7934 4564
rect 9650 4508 9660 4564
rect 9716 4508 13692 4564
rect 13748 4508 13758 4564
rect 20514 4508 20524 4564
rect 20580 4508 21868 4564
rect 21924 4508 21934 4564
rect 0 4340 800 4368
rect 1484 4340 1540 4508
rect 6076 4452 6132 4508
rect 2818 4396 2828 4452
rect 2884 4396 4060 4452
rect 4116 4396 4126 4452
rect 6066 4396 6076 4452
rect 6132 4396 6142 4452
rect 8866 4396 8876 4452
rect 8932 4396 10892 4452
rect 10948 4396 11788 4452
rect 11844 4396 11854 4452
rect 14242 4396 14252 4452
rect 14308 4396 15484 4452
rect 15540 4396 15550 4452
rect 16604 4396 18508 4452
rect 18564 4396 19068 4452
rect 19124 4396 19134 4452
rect 16604 4340 16660 4396
rect 0 4284 1540 4340
rect 2482 4284 2492 4340
rect 2548 4284 3164 4340
rect 3220 4284 3230 4340
rect 3490 4284 3500 4340
rect 3556 4284 13020 4340
rect 13076 4284 13086 4340
rect 14354 4284 14364 4340
rect 14420 4284 16660 4340
rect 16818 4284 16828 4340
rect 16884 4284 21420 4340
rect 21476 4284 21486 4340
rect 0 4256 800 4284
rect 3938 4172 3948 4228
rect 4004 4172 5124 4228
rect 5730 4172 5740 4228
rect 5796 4172 7196 4228
rect 7252 4172 7262 4228
rect 9986 4172 9996 4228
rect 10052 4172 10668 4228
rect 10724 4172 10734 4228
rect 17490 4172 17500 4228
rect 17556 4172 18620 4228
rect 18676 4172 18686 4228
rect 5068 4116 5124 4172
rect 4274 4060 4284 4116
rect 4340 4060 4844 4116
rect 4900 4060 4910 4116
rect 5068 4060 13916 4116
rect 13972 4060 13982 4116
rect 4722 3948 4732 4004
rect 4788 3948 8260 4004
rect 0 3892 800 3920
rect 3862 3892 3872 3948
rect 3928 3892 3976 3948
rect 4032 3892 4080 3948
rect 4136 3892 4146 3948
rect 0 3836 1988 3892
rect 0 3808 800 3836
rect 1932 3780 1988 3836
rect 8204 3780 8260 3948
rect 9182 3892 9192 3948
rect 9248 3892 9296 3948
rect 9352 3892 9400 3948
rect 9456 3892 9466 3948
rect 14502 3892 14512 3948
rect 14568 3892 14616 3948
rect 14672 3892 14720 3948
rect 14776 3892 14786 3948
rect 19822 3892 19832 3948
rect 19888 3892 19936 3948
rect 19992 3892 20040 3948
rect 20096 3892 20106 3948
rect 1922 3724 1932 3780
rect 1988 3724 1998 3780
rect 5954 3724 5964 3780
rect 6020 3724 6972 3780
rect 7028 3724 7038 3780
rect 8204 3724 15148 3780
rect 15204 3724 15214 3780
rect 15922 3724 15932 3780
rect 15988 3724 18732 3780
rect 18788 3724 21532 3780
rect 21588 3724 21598 3780
rect 6290 3612 6300 3668
rect 6356 3612 7084 3668
rect 7140 3612 7150 3668
rect 8642 3612 8652 3668
rect 8708 3612 12572 3668
rect 12628 3612 12638 3668
rect 13570 3612 13580 3668
rect 13636 3612 20972 3668
rect 21028 3612 21038 3668
rect 3490 3500 3500 3556
rect 3556 3500 3724 3556
rect 3780 3500 3790 3556
rect 4274 3500 4284 3556
rect 4340 3500 5628 3556
rect 5684 3500 5694 3556
rect 6402 3500 6412 3556
rect 6468 3500 10164 3556
rect 12674 3500 12684 3556
rect 12740 3500 16828 3556
rect 16884 3500 16894 3556
rect 0 3444 800 3472
rect 10108 3444 10164 3500
rect 0 3388 3052 3444
rect 3108 3388 3118 3444
rect 4722 3388 4732 3444
rect 4788 3388 7980 3444
rect 8036 3388 8046 3444
rect 8306 3388 8316 3444
rect 8372 3388 9884 3444
rect 9940 3388 9950 3444
rect 10098 3388 10108 3444
rect 10164 3388 10174 3444
rect 13010 3388 13020 3444
rect 13076 3388 15708 3444
rect 15764 3388 15774 3444
rect 16706 3388 16716 3444
rect 16772 3388 20748 3444
rect 20804 3388 20814 3444
rect 0 3360 800 3388
rect 6402 3276 6412 3332
rect 6468 3276 9324 3332
rect 9380 3276 9390 3332
rect 13234 3276 13244 3332
rect 13300 3276 13692 3332
rect 13748 3276 13758 3332
rect 6522 3108 6532 3164
rect 6588 3108 6636 3164
rect 6692 3108 6740 3164
rect 6796 3108 6806 3164
rect 11842 3108 11852 3164
rect 11908 3108 11956 3164
rect 12012 3108 12060 3164
rect 12116 3108 12126 3164
rect 17162 3108 17172 3164
rect 17228 3108 17276 3164
rect 17332 3108 17380 3164
rect 17436 3108 17446 3164
rect 22482 3108 22492 3164
rect 22548 3108 22596 3164
rect 22652 3108 22700 3164
rect 22756 3108 22766 3164
rect 0 2996 800 3024
rect 0 2940 2492 2996
rect 2548 2940 2558 2996
rect 0 2912 800 2940
rect 0 2548 800 2576
rect 23200 2548 24000 2576
rect 0 2492 1708 2548
rect 1764 2492 1774 2548
rect 22306 2492 22316 2548
rect 22372 2492 24000 2548
rect 0 2464 800 2492
rect 23200 2464 24000 2492
<< via3 >>
rect 3872 16436 3928 16492
rect 3976 16436 4032 16492
rect 4080 16436 4136 16492
rect 9192 16436 9248 16492
rect 9296 16436 9352 16492
rect 9400 16436 9456 16492
rect 14512 16436 14568 16492
rect 14616 16436 14672 16492
rect 14720 16436 14776 16492
rect 19832 16436 19888 16492
rect 19936 16436 19992 16492
rect 20040 16436 20096 16492
rect 6532 15652 6588 15708
rect 6636 15652 6692 15708
rect 6740 15652 6796 15708
rect 11852 15652 11908 15708
rect 11956 15652 12012 15708
rect 12060 15652 12116 15708
rect 17172 15652 17228 15708
rect 17276 15652 17332 15708
rect 17380 15652 17436 15708
rect 22492 15652 22548 15708
rect 22596 15652 22652 15708
rect 22700 15652 22756 15708
rect 3872 14868 3928 14924
rect 3976 14868 4032 14924
rect 4080 14868 4136 14924
rect 9192 14868 9248 14924
rect 9296 14868 9352 14924
rect 9400 14868 9456 14924
rect 14512 14868 14568 14924
rect 14616 14868 14672 14924
rect 14720 14868 14776 14924
rect 19832 14868 19888 14924
rect 19936 14868 19992 14924
rect 20040 14868 20096 14924
rect 6532 14084 6588 14140
rect 6636 14084 6692 14140
rect 6740 14084 6796 14140
rect 11852 14084 11908 14140
rect 11956 14084 12012 14140
rect 12060 14084 12116 14140
rect 17172 14084 17228 14140
rect 17276 14084 17332 14140
rect 17380 14084 17436 14140
rect 22492 14084 22548 14140
rect 22596 14084 22652 14140
rect 22700 14084 22756 14140
rect 3872 13300 3928 13356
rect 3976 13300 4032 13356
rect 4080 13300 4136 13356
rect 9192 13300 9248 13356
rect 9296 13300 9352 13356
rect 9400 13300 9456 13356
rect 14512 13300 14568 13356
rect 14616 13300 14672 13356
rect 14720 13300 14776 13356
rect 19832 13300 19888 13356
rect 19936 13300 19992 13356
rect 20040 13300 20096 13356
rect 6532 12516 6588 12572
rect 6636 12516 6692 12572
rect 6740 12516 6796 12572
rect 11852 12516 11908 12572
rect 11956 12516 12012 12572
rect 12060 12516 12116 12572
rect 17172 12516 17228 12572
rect 17276 12516 17332 12572
rect 17380 12516 17436 12572
rect 22492 12516 22548 12572
rect 22596 12516 22652 12572
rect 22700 12516 22756 12572
rect 3724 12012 3780 12068
rect 3872 11732 3928 11788
rect 3976 11732 4032 11788
rect 4080 11732 4136 11788
rect 9192 11732 9248 11788
rect 9296 11732 9352 11788
rect 9400 11732 9456 11788
rect 14512 11732 14568 11788
rect 14616 11732 14672 11788
rect 14720 11732 14776 11788
rect 19832 11732 19888 11788
rect 19936 11732 19992 11788
rect 20040 11732 20096 11788
rect 4844 11452 4900 11508
rect 2492 11116 2548 11172
rect 3388 11116 3444 11172
rect 6532 10948 6588 11004
rect 6636 10948 6692 11004
rect 6740 10948 6796 11004
rect 11852 10948 11908 11004
rect 11956 10948 12012 11004
rect 12060 10948 12116 11004
rect 17172 10948 17228 11004
rect 17276 10948 17332 11004
rect 17380 10948 17436 11004
rect 22492 10948 22548 11004
rect 22596 10948 22652 11004
rect 22700 10948 22756 11004
rect 4508 10892 4564 10948
rect 2380 10556 2436 10612
rect 12460 10444 12516 10500
rect 3872 10164 3928 10220
rect 3976 10164 4032 10220
rect 4080 10164 4136 10220
rect 9192 10164 9248 10220
rect 9296 10164 9352 10220
rect 9400 10164 9456 10220
rect 14512 10164 14568 10220
rect 14616 10164 14672 10220
rect 14720 10164 14776 10220
rect 19832 10164 19888 10220
rect 19936 10164 19992 10220
rect 20040 10164 20096 10220
rect 2044 9548 2100 9604
rect 5068 9548 5124 9604
rect 7420 9548 7476 9604
rect 6532 9380 6588 9436
rect 6636 9380 6692 9436
rect 6740 9380 6796 9436
rect 11852 9380 11908 9436
rect 11956 9380 12012 9436
rect 12060 9380 12116 9436
rect 17172 9380 17228 9436
rect 17276 9380 17332 9436
rect 17380 9380 17436 9436
rect 22492 9380 22548 9436
rect 22596 9380 22652 9436
rect 22700 9380 22756 9436
rect 1820 9324 1876 9380
rect 2716 9100 2772 9156
rect 6076 9100 6132 9156
rect 5404 8764 5460 8820
rect 4620 8652 4676 8708
rect 3872 8596 3928 8652
rect 3976 8596 4032 8652
rect 4080 8596 4136 8652
rect 9192 8596 9248 8652
rect 9296 8596 9352 8652
rect 9400 8596 9456 8652
rect 14512 8596 14568 8652
rect 14616 8596 14672 8652
rect 14720 8596 14776 8652
rect 19832 8596 19888 8652
rect 19936 8596 19992 8652
rect 20040 8596 20096 8652
rect 8316 8540 8372 8596
rect 2604 8428 2660 8484
rect 12236 8204 12292 8260
rect 12460 8204 12516 8260
rect 3500 8092 3556 8148
rect 5740 8092 5796 8148
rect 3388 7980 3444 8036
rect 3612 7980 3668 8036
rect 1820 7868 1876 7924
rect 5068 7868 5124 7924
rect 7420 7868 7476 7924
rect 6532 7812 6588 7868
rect 6636 7812 6692 7868
rect 6740 7812 6796 7868
rect 11852 7812 11908 7868
rect 11956 7812 12012 7868
rect 12060 7812 12116 7868
rect 17172 7812 17228 7868
rect 17276 7812 17332 7868
rect 17380 7812 17436 7868
rect 22492 7812 22548 7868
rect 22596 7812 22652 7868
rect 22700 7812 22756 7868
rect 2380 7756 2436 7812
rect 2604 7644 2660 7700
rect 3500 7644 3556 7700
rect 2492 7532 2548 7588
rect 13692 7420 13748 7476
rect 3500 7196 3556 7252
rect 3388 7084 3444 7140
rect 4732 7084 4788 7140
rect 6188 7084 6244 7140
rect 18620 7084 18676 7140
rect 3872 7028 3928 7084
rect 3976 7028 4032 7084
rect 4080 7028 4136 7084
rect 9192 7028 9248 7084
rect 9296 7028 9352 7084
rect 9400 7028 9456 7084
rect 14512 7028 14568 7084
rect 14616 7028 14672 7084
rect 14720 7028 14776 7084
rect 19832 7028 19888 7084
rect 19936 7028 19992 7084
rect 20040 7028 20096 7084
rect 2044 6972 2100 7028
rect 5628 6860 5684 6916
rect 6188 6748 6244 6804
rect 4620 6636 4676 6692
rect 7420 6636 7476 6692
rect 5628 6524 5684 6580
rect 6076 6300 6132 6356
rect 6532 6244 6588 6300
rect 6636 6244 6692 6300
rect 6740 6244 6796 6300
rect 11852 6244 11908 6300
rect 11956 6244 12012 6300
rect 12060 6244 12116 6300
rect 5404 6188 5460 6244
rect 6300 6188 6356 6244
rect 17172 6244 17228 6300
rect 17276 6244 17332 6300
rect 17380 6244 17436 6300
rect 22492 6244 22548 6300
rect 22596 6244 22652 6300
rect 22700 6244 22756 6300
rect 3612 5964 3668 6020
rect 19628 5852 19684 5908
rect 4508 5740 4564 5796
rect 4956 5740 5012 5796
rect 6300 5740 6356 5796
rect 3724 5516 3780 5572
rect 4732 5516 4788 5572
rect 5068 5516 5124 5572
rect 3872 5460 3928 5516
rect 3976 5460 4032 5516
rect 4080 5460 4136 5516
rect 9192 5460 9248 5516
rect 9296 5460 9352 5516
rect 9400 5460 9456 5516
rect 2716 5180 2772 5236
rect 4844 5180 4900 5236
rect 14512 5460 14568 5516
rect 14616 5460 14672 5516
rect 14720 5460 14776 5516
rect 19832 5460 19888 5516
rect 19936 5460 19992 5516
rect 20040 5460 20096 5516
rect 8316 5068 8372 5124
rect 19628 5068 19684 5124
rect 12236 4956 12292 5012
rect 1820 4844 1876 4900
rect 4732 4844 4788 4900
rect 4956 4844 5012 4900
rect 6532 4676 6588 4732
rect 6636 4676 6692 4732
rect 6740 4676 6796 4732
rect 11852 4676 11908 4732
rect 11956 4676 12012 4732
rect 12060 4676 12116 4732
rect 17172 4676 17228 4732
rect 17276 4676 17332 4732
rect 17380 4676 17436 4732
rect 22492 4676 22548 4732
rect 22596 4676 22652 4732
rect 22700 4676 22756 4732
rect 8316 4620 8372 4676
rect 5740 4172 5796 4228
rect 18620 4172 18676 4228
rect 4732 3948 4788 4004
rect 3872 3892 3928 3948
rect 3976 3892 4032 3948
rect 4080 3892 4136 3948
rect 9192 3892 9248 3948
rect 9296 3892 9352 3948
rect 9400 3892 9456 3948
rect 14512 3892 14568 3948
rect 14616 3892 14672 3948
rect 14720 3892 14776 3948
rect 19832 3892 19888 3948
rect 19936 3892 19992 3948
rect 20040 3892 20096 3948
rect 3500 3500 3556 3556
rect 13692 3276 13748 3332
rect 6532 3108 6588 3164
rect 6636 3108 6692 3164
rect 6740 3108 6796 3164
rect 11852 3108 11908 3164
rect 11956 3108 12012 3164
rect 12060 3108 12116 3164
rect 17172 3108 17228 3164
rect 17276 3108 17332 3164
rect 17380 3108 17436 3164
rect 22492 3108 22548 3164
rect 22596 3108 22652 3164
rect 22700 3108 22756 3164
<< metal4 >>
rect 3844 16492 4164 16524
rect 3844 16436 3872 16492
rect 3928 16436 3976 16492
rect 4032 16436 4080 16492
rect 4136 16436 4164 16492
rect 3844 14924 4164 16436
rect 3844 14868 3872 14924
rect 3928 14868 3976 14924
rect 4032 14868 4080 14924
rect 4136 14868 4164 14924
rect 3844 13356 4164 14868
rect 3844 13300 3872 13356
rect 3928 13300 3976 13356
rect 4032 13300 4080 13356
rect 4136 13300 4164 13356
rect 3724 12068 3780 12078
rect 2492 11172 2548 11182
rect 2380 10612 2436 10622
rect 2044 9604 2100 9614
rect 1820 9380 1876 9390
rect 1820 7924 1876 9324
rect 1820 4900 1876 7868
rect 2044 7028 2100 9548
rect 2380 7812 2436 10556
rect 2380 7746 2436 7756
rect 2492 7588 2548 11116
rect 3388 11172 3444 11182
rect 2716 9156 2772 9166
rect 2604 8484 2660 8494
rect 2604 7700 2660 8428
rect 2604 7634 2660 7644
rect 2492 7522 2548 7532
rect 2044 6962 2100 6972
rect 2716 5236 2772 9100
rect 3388 8036 3444 11116
rect 3388 7140 3444 7980
rect 3500 8148 3556 8158
rect 3500 7700 3556 8092
rect 3500 7634 3556 7644
rect 3612 8036 3668 8046
rect 3388 7074 3444 7084
rect 3500 7252 3556 7262
rect 2716 5170 2772 5180
rect 1820 4834 1876 4844
rect 3500 3556 3556 7196
rect 3612 6020 3668 7980
rect 3612 5954 3668 5964
rect 3724 5572 3780 12012
rect 3724 5506 3780 5516
rect 3844 11788 4164 13300
rect 3844 11732 3872 11788
rect 3928 11732 3976 11788
rect 4032 11732 4080 11788
rect 4136 11732 4164 11788
rect 3844 10220 4164 11732
rect 6504 15708 6824 16524
rect 6504 15652 6532 15708
rect 6588 15652 6636 15708
rect 6692 15652 6740 15708
rect 6796 15652 6824 15708
rect 6504 14140 6824 15652
rect 6504 14084 6532 14140
rect 6588 14084 6636 14140
rect 6692 14084 6740 14140
rect 6796 14084 6824 14140
rect 6504 12572 6824 14084
rect 6504 12516 6532 12572
rect 6588 12516 6636 12572
rect 6692 12516 6740 12572
rect 6796 12516 6824 12572
rect 4844 11508 4900 11518
rect 3844 10164 3872 10220
rect 3928 10164 3976 10220
rect 4032 10164 4080 10220
rect 4136 10164 4164 10220
rect 3844 8652 4164 10164
rect 3844 8596 3872 8652
rect 3928 8596 3976 8652
rect 4032 8596 4080 8652
rect 4136 8596 4164 8652
rect 3844 7084 4164 8596
rect 3844 7028 3872 7084
rect 3928 7028 3976 7084
rect 4032 7028 4080 7084
rect 4136 7028 4164 7084
rect 3844 5516 4164 7028
rect 4508 10948 4564 10958
rect 4508 5796 4564 10892
rect 4620 8708 4676 8718
rect 4620 6692 4676 8652
rect 4620 6626 4676 6636
rect 4732 7140 4788 7150
rect 4508 5730 4564 5740
rect 3500 3490 3556 3500
rect 3844 5460 3872 5516
rect 3928 5460 3976 5516
rect 4032 5460 4080 5516
rect 4136 5460 4164 5516
rect 4732 5572 4788 7084
rect 4732 5506 4788 5516
rect 3844 3948 4164 5460
rect 4844 5236 4900 11452
rect 6504 11004 6824 12516
rect 6504 10948 6532 11004
rect 6588 10948 6636 11004
rect 6692 10948 6740 11004
rect 6796 10948 6824 11004
rect 5068 9604 5124 9614
rect 5068 7924 5124 9548
rect 6504 9436 6824 10948
rect 9164 16492 9484 16524
rect 9164 16436 9192 16492
rect 9248 16436 9296 16492
rect 9352 16436 9400 16492
rect 9456 16436 9484 16492
rect 9164 14924 9484 16436
rect 9164 14868 9192 14924
rect 9248 14868 9296 14924
rect 9352 14868 9400 14924
rect 9456 14868 9484 14924
rect 9164 13356 9484 14868
rect 9164 13300 9192 13356
rect 9248 13300 9296 13356
rect 9352 13300 9400 13356
rect 9456 13300 9484 13356
rect 9164 11788 9484 13300
rect 9164 11732 9192 11788
rect 9248 11732 9296 11788
rect 9352 11732 9400 11788
rect 9456 11732 9484 11788
rect 9164 10220 9484 11732
rect 9164 10164 9192 10220
rect 9248 10164 9296 10220
rect 9352 10164 9400 10220
rect 9456 10164 9484 10220
rect 6504 9380 6532 9436
rect 6588 9380 6636 9436
rect 6692 9380 6740 9436
rect 6796 9380 6824 9436
rect 6076 9156 6132 9166
rect 4844 5170 4900 5180
rect 4956 5796 5012 5806
rect 3844 3892 3872 3948
rect 3928 3892 3976 3948
rect 4032 3892 4080 3948
rect 4136 3892 4164 3948
rect 4732 4900 4788 4910
rect 4732 4004 4788 4844
rect 4956 4900 5012 5740
rect 5068 5572 5124 7868
rect 5404 8820 5460 8830
rect 5404 6244 5460 8764
rect 5740 8148 5796 8158
rect 5628 6916 5684 6926
rect 5628 6580 5684 6860
rect 5628 6514 5684 6524
rect 5404 6178 5460 6188
rect 5068 5506 5124 5516
rect 4956 4834 5012 4844
rect 5740 4228 5796 8092
rect 6076 6356 6132 9100
rect 6504 7868 6824 9380
rect 6504 7812 6532 7868
rect 6588 7812 6636 7868
rect 6692 7812 6740 7868
rect 6796 7812 6824 7868
rect 6188 7140 6244 7150
rect 6188 6804 6244 7084
rect 6188 6738 6244 6748
rect 6076 6290 6132 6300
rect 6504 6300 6824 7812
rect 7420 9604 7476 9614
rect 7420 7924 7476 9548
rect 9164 8652 9484 10164
rect 7420 6692 7476 7868
rect 7420 6626 7476 6636
rect 8316 8596 8372 8606
rect 6300 6244 6356 6254
rect 6300 5796 6356 6188
rect 6300 5730 6356 5740
rect 6504 6244 6532 6300
rect 6588 6244 6636 6300
rect 6692 6244 6740 6300
rect 6796 6244 6824 6300
rect 5740 4162 5796 4172
rect 6504 4732 6824 6244
rect 6504 4676 6532 4732
rect 6588 4676 6636 4732
rect 6692 4676 6740 4732
rect 6796 4676 6824 4732
rect 4732 3938 4788 3948
rect 3844 3076 4164 3892
rect 6504 3164 6824 4676
rect 8316 5124 8372 8540
rect 8316 4676 8372 5068
rect 8316 4610 8372 4620
rect 9164 8596 9192 8652
rect 9248 8596 9296 8652
rect 9352 8596 9400 8652
rect 9456 8596 9484 8652
rect 9164 7084 9484 8596
rect 9164 7028 9192 7084
rect 9248 7028 9296 7084
rect 9352 7028 9400 7084
rect 9456 7028 9484 7084
rect 9164 5516 9484 7028
rect 9164 5460 9192 5516
rect 9248 5460 9296 5516
rect 9352 5460 9400 5516
rect 9456 5460 9484 5516
rect 6504 3108 6532 3164
rect 6588 3108 6636 3164
rect 6692 3108 6740 3164
rect 6796 3108 6824 3164
rect 6504 3076 6824 3108
rect 9164 3948 9484 5460
rect 9164 3892 9192 3948
rect 9248 3892 9296 3948
rect 9352 3892 9400 3948
rect 9456 3892 9484 3948
rect 9164 3076 9484 3892
rect 11824 15708 12144 16524
rect 11824 15652 11852 15708
rect 11908 15652 11956 15708
rect 12012 15652 12060 15708
rect 12116 15652 12144 15708
rect 11824 14140 12144 15652
rect 11824 14084 11852 14140
rect 11908 14084 11956 14140
rect 12012 14084 12060 14140
rect 12116 14084 12144 14140
rect 11824 12572 12144 14084
rect 11824 12516 11852 12572
rect 11908 12516 11956 12572
rect 12012 12516 12060 12572
rect 12116 12516 12144 12572
rect 11824 11004 12144 12516
rect 11824 10948 11852 11004
rect 11908 10948 11956 11004
rect 12012 10948 12060 11004
rect 12116 10948 12144 11004
rect 11824 9436 12144 10948
rect 14484 16492 14804 16524
rect 14484 16436 14512 16492
rect 14568 16436 14616 16492
rect 14672 16436 14720 16492
rect 14776 16436 14804 16492
rect 14484 14924 14804 16436
rect 14484 14868 14512 14924
rect 14568 14868 14616 14924
rect 14672 14868 14720 14924
rect 14776 14868 14804 14924
rect 14484 13356 14804 14868
rect 14484 13300 14512 13356
rect 14568 13300 14616 13356
rect 14672 13300 14720 13356
rect 14776 13300 14804 13356
rect 14484 11788 14804 13300
rect 14484 11732 14512 11788
rect 14568 11732 14616 11788
rect 14672 11732 14720 11788
rect 14776 11732 14804 11788
rect 11824 9380 11852 9436
rect 11908 9380 11956 9436
rect 12012 9380 12060 9436
rect 12116 9380 12144 9436
rect 11824 7868 12144 9380
rect 12460 10500 12516 10510
rect 11824 7812 11852 7868
rect 11908 7812 11956 7868
rect 12012 7812 12060 7868
rect 12116 7812 12144 7868
rect 11824 6300 12144 7812
rect 11824 6244 11852 6300
rect 11908 6244 11956 6300
rect 12012 6244 12060 6300
rect 12116 6244 12144 6300
rect 11824 4732 12144 6244
rect 12236 8260 12292 8270
rect 12236 5012 12292 8204
rect 12460 8260 12516 10444
rect 12460 8194 12516 8204
rect 14484 10220 14804 11732
rect 14484 10164 14512 10220
rect 14568 10164 14616 10220
rect 14672 10164 14720 10220
rect 14776 10164 14804 10220
rect 14484 8652 14804 10164
rect 14484 8596 14512 8652
rect 14568 8596 14616 8652
rect 14672 8596 14720 8652
rect 14776 8596 14804 8652
rect 12236 4946 12292 4956
rect 13692 7476 13748 7486
rect 11824 4676 11852 4732
rect 11908 4676 11956 4732
rect 12012 4676 12060 4732
rect 12116 4676 12144 4732
rect 11824 3164 12144 4676
rect 13692 3332 13748 7420
rect 13692 3266 13748 3276
rect 14484 7084 14804 8596
rect 14484 7028 14512 7084
rect 14568 7028 14616 7084
rect 14672 7028 14720 7084
rect 14776 7028 14804 7084
rect 14484 5516 14804 7028
rect 14484 5460 14512 5516
rect 14568 5460 14616 5516
rect 14672 5460 14720 5516
rect 14776 5460 14804 5516
rect 14484 3948 14804 5460
rect 14484 3892 14512 3948
rect 14568 3892 14616 3948
rect 14672 3892 14720 3948
rect 14776 3892 14804 3948
rect 11824 3108 11852 3164
rect 11908 3108 11956 3164
rect 12012 3108 12060 3164
rect 12116 3108 12144 3164
rect 11824 3076 12144 3108
rect 14484 3076 14804 3892
rect 17144 15708 17464 16524
rect 17144 15652 17172 15708
rect 17228 15652 17276 15708
rect 17332 15652 17380 15708
rect 17436 15652 17464 15708
rect 17144 14140 17464 15652
rect 17144 14084 17172 14140
rect 17228 14084 17276 14140
rect 17332 14084 17380 14140
rect 17436 14084 17464 14140
rect 17144 12572 17464 14084
rect 17144 12516 17172 12572
rect 17228 12516 17276 12572
rect 17332 12516 17380 12572
rect 17436 12516 17464 12572
rect 17144 11004 17464 12516
rect 17144 10948 17172 11004
rect 17228 10948 17276 11004
rect 17332 10948 17380 11004
rect 17436 10948 17464 11004
rect 17144 9436 17464 10948
rect 17144 9380 17172 9436
rect 17228 9380 17276 9436
rect 17332 9380 17380 9436
rect 17436 9380 17464 9436
rect 17144 7868 17464 9380
rect 17144 7812 17172 7868
rect 17228 7812 17276 7868
rect 17332 7812 17380 7868
rect 17436 7812 17464 7868
rect 17144 6300 17464 7812
rect 19804 16492 20124 16524
rect 19804 16436 19832 16492
rect 19888 16436 19936 16492
rect 19992 16436 20040 16492
rect 20096 16436 20124 16492
rect 19804 14924 20124 16436
rect 19804 14868 19832 14924
rect 19888 14868 19936 14924
rect 19992 14868 20040 14924
rect 20096 14868 20124 14924
rect 19804 13356 20124 14868
rect 19804 13300 19832 13356
rect 19888 13300 19936 13356
rect 19992 13300 20040 13356
rect 20096 13300 20124 13356
rect 19804 11788 20124 13300
rect 19804 11732 19832 11788
rect 19888 11732 19936 11788
rect 19992 11732 20040 11788
rect 20096 11732 20124 11788
rect 19804 10220 20124 11732
rect 19804 10164 19832 10220
rect 19888 10164 19936 10220
rect 19992 10164 20040 10220
rect 20096 10164 20124 10220
rect 19804 8652 20124 10164
rect 19804 8596 19832 8652
rect 19888 8596 19936 8652
rect 19992 8596 20040 8652
rect 20096 8596 20124 8652
rect 17144 6244 17172 6300
rect 17228 6244 17276 6300
rect 17332 6244 17380 6300
rect 17436 6244 17464 6300
rect 17144 4732 17464 6244
rect 17144 4676 17172 4732
rect 17228 4676 17276 4732
rect 17332 4676 17380 4732
rect 17436 4676 17464 4732
rect 17144 3164 17464 4676
rect 18620 7140 18676 7150
rect 18620 4228 18676 7084
rect 19804 7084 20124 8596
rect 19804 7028 19832 7084
rect 19888 7028 19936 7084
rect 19992 7028 20040 7084
rect 20096 7028 20124 7084
rect 19628 5908 19684 5918
rect 19628 5124 19684 5852
rect 19628 5058 19684 5068
rect 19804 5516 20124 7028
rect 19804 5460 19832 5516
rect 19888 5460 19936 5516
rect 19992 5460 20040 5516
rect 20096 5460 20124 5516
rect 18620 4162 18676 4172
rect 17144 3108 17172 3164
rect 17228 3108 17276 3164
rect 17332 3108 17380 3164
rect 17436 3108 17464 3164
rect 17144 3076 17464 3108
rect 19804 3948 20124 5460
rect 19804 3892 19832 3948
rect 19888 3892 19936 3948
rect 19992 3892 20040 3948
rect 20096 3892 20124 3948
rect 19804 3076 20124 3892
rect 22464 15708 22784 16524
rect 22464 15652 22492 15708
rect 22548 15652 22596 15708
rect 22652 15652 22700 15708
rect 22756 15652 22784 15708
rect 22464 14140 22784 15652
rect 22464 14084 22492 14140
rect 22548 14084 22596 14140
rect 22652 14084 22700 14140
rect 22756 14084 22784 14140
rect 22464 12572 22784 14084
rect 22464 12516 22492 12572
rect 22548 12516 22596 12572
rect 22652 12516 22700 12572
rect 22756 12516 22784 12572
rect 22464 11004 22784 12516
rect 22464 10948 22492 11004
rect 22548 10948 22596 11004
rect 22652 10948 22700 11004
rect 22756 10948 22784 11004
rect 22464 9436 22784 10948
rect 22464 9380 22492 9436
rect 22548 9380 22596 9436
rect 22652 9380 22700 9436
rect 22756 9380 22784 9436
rect 22464 7868 22784 9380
rect 22464 7812 22492 7868
rect 22548 7812 22596 7868
rect 22652 7812 22700 7868
rect 22756 7812 22784 7868
rect 22464 6300 22784 7812
rect 22464 6244 22492 6300
rect 22548 6244 22596 6300
rect 22652 6244 22700 6300
rect 22756 6244 22784 6300
rect 22464 4732 22784 6244
rect 22464 4676 22492 4732
rect 22548 4676 22596 4732
rect 22652 4676 22700 4732
rect 22756 4676 22784 4732
rect 22464 3164 22784 4676
rect 22464 3108 22492 3164
rect 22548 3108 22596 3164
rect 22652 3108 22700 3164
rect 22756 3108 22784 3164
rect 22464 3076 22784 3108
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _042_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 16464 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _043_
timestamp 1698431365
transform 1 0 12544 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _044_
timestamp 1698431365
transform -1 0 7280 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _045_
timestamp 1698431365
transform -1 0 22288 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _046_
timestamp 1698431365
transform -1 0 21056 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _047_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 21392 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _048_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 9184 0 -1 4704
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _049_
timestamp 1698431365
transform 1 0 9408 0 -1 9408
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _050_
timestamp 1698431365
transform 1 0 7728 0 1 7840
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  _051_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 9968 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _052_
timestamp 1698431365
transform -1 0 18592 0 1 4704
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _053_
timestamp 1698431365
transform -1 0 17024 0 -1 4704
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  _054_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 15344 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _055_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 21168 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _056_
timestamp 1698431365
transform -1 0 21392 0 -1 4704
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _057_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 20384 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _058_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 7392 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _059_
timestamp 1698431365
transform 1 0 5040 0 -1 6272
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _060_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5488 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _061_
timestamp 1698431365
transform 1 0 9408 0 -1 7840
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _062_
timestamp 1698431365
transform -1 0 7392 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _063_
timestamp 1698431365
transform 1 0 5040 0 -1 7840
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _064_
timestamp 1698431365
transform -1 0 2352 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _065_
timestamp 1698431365
transform -1 0 3584 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _066_
timestamp 1698431365
transform -1 0 3584 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _067_
timestamp 1698431365
transform -1 0 5152 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _068_
timestamp 1698431365
transform 1 0 4368 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _069_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 5152 0 1 3136
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _070_
timestamp 1698431365
transform 1 0 12992 0 1 3136
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _071_
timestamp 1698431365
transform 1 0 9184 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _072_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 6048 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _073_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 5264 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _074_
timestamp 1698431365
transform -1 0 10528 0 -1 6272
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _075_
timestamp 1698431365
transform -1 0 9968 0 -1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _076_
timestamp 1698431365
transform 1 0 6832 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _077_
timestamp 1698431365
transform -1 0 9184 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _078_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 6832 0 1 3136
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _079_
timestamp 1698431365
transform 1 0 8960 0 1 4704
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _080_
timestamp 1698431365
transform 1 0 17248 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _081_
timestamp 1698431365
transform 1 0 17248 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _082_
timestamp 1698431365
transform 1 0 13328 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _083_
timestamp 1698431365
transform -1 0 14448 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _084_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 5040 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _085_
timestamp 1698431365
transform -1 0 6832 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _086_
timestamp 1698431365
transform -1 0 8960 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _087_
timestamp 1698431365
transform -1 0 16800 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _088_
timestamp 1698431365
transform 1 0 13328 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _089_
timestamp 1698431365
transform -1 0 21392 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _090_
timestamp 1698431365
transform -1 0 5264 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__065__A2 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 4368 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__069__A1
timestamp 1698431365
transform -1 0 6608 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__072__B
timestamp 1698431365
transform 1 0 6944 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__075__A1
timestamp 1698431365
transform 1 0 9968 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__076__B
timestamp 1698431365
transform 1 0 7392 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__080__B
timestamp 1698431365
transform 1 0 19488 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__082__A1
timestamp 1698431365
transform 1 0 15120 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__082__B
timestamp 1698431365
transform 1 0 14672 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__089__D
timestamp 1698431365
transform 1 0 22176 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__090__D
timestamp 1698431365
transform 1 0 5936 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I
timestamp 1698431365
transform -1 0 17472 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1698431365
transform -1 0 22400 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1698431365
transform -1 0 21728 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1698431365
transform -1 0 21616 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1698431365
transform 1 0 4592 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1698431365
transform -1 0 5712 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1698431365
transform 1 0 10640 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input7_I
timestamp 1698431365
transform 1 0 11088 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input8_I
timestamp 1698431365
transform 1 0 12656 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input9_I
timestamp 1698431365
transform -1 0 11760 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input10_I
timestamp 1698431365
transform -1 0 12208 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input11_I
timestamp 1698431365
transform -1 0 3920 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input12_I
timestamp 1698431365
transform 1 0 22176 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input13_I
timestamp 1698431365
transform -1 0 20608 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input14_I
timestamp 1698431365
transform -1 0 5040 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input15_I
timestamp 1698431365
transform -1 0 2912 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input16_I
timestamp 1698431365
transform -1 0 18592 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input17_I
timestamp 1698431365
transform 1 0 16800 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input18_I
timestamp 1698431365
transform 1 0 19824 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input19_I
timestamp 1698431365
transform -1 0 20160 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input20_I
timestamp 1698431365
transform -1 0 18144 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input21_I
timestamp 1698431365
transform -1 0 19152 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input22_I
timestamp 1698431365
transform -1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input23_I
timestamp 1698431365
transform 1 0 19040 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input24_I
timestamp 1698431365
transform -1 0 19600 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input25_I
timestamp 1698431365
transform -1 0 20496 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input26_I
timestamp 1698431365
transform -1 0 3360 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input27_I
timestamp 1698431365
transform 1 0 22064 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input28_I
timestamp 1698431365
transform 1 0 20720 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input29_I
timestamp 1698431365
transform -1 0 4592 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input30_I
timestamp 1698431365
transform -1 0 6384 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input31_I
timestamp 1698431365
transform 1 0 7840 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input32_I
timestamp 1698431365
transform -1 0 7056 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input33_I
timestamp 1698431365
transform -1 0 5264 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input34_I
timestamp 1698431365
transform 1 0 8960 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input35_I
timestamp 1698431365
transform -1 0 8512 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input36_I
timestamp 1698431365
transform 1 0 3696 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input37_I
timestamp 1698431365
transform -1 0 2912 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input38_I
timestamp 1698431365
transform -1 0 5936 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input39_I
timestamp 1698431365
transform -1 0 3472 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input40_I
timestamp 1698431365
transform -1 0 4144 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input41_I
timestamp 1698431365
transform -1 0 21168 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output43_I
timestamp 1698431365
transform -1 0 20384 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output48_I
timestamp 1698431365
transform 1 0 9408 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 16352 0 -1 6272
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1698431365
transform -1 0 12544 0 1 6272
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1698431365
transform 1 0 13328 0 1 6272
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_2 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_53 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 7280 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_135
timestamp 1698431365
transform 1 0 16464 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_184
timestamp 1698431365
transform 1 0 21952 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_2
timestamp 1698431365
transform 1 0 1568 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_185
timestamp 1698431365
transform 1 0 22064 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_187
timestamp 1698431365
transform 1 0 22288 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_12
timestamp 1698431365
transform 1 0 2688 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_14
timestamp 1698431365
transform 1 0 2912 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_37
timestamp 1698431365
transform 1 0 5488 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_115
timestamp 1698431365
transform 1 0 14224 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_172
timestamp 1698431365
transform 1 0 20608 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_174
timestamp 1698431365
transform 1 0 20832 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_187
timestamp 1698431365
transform 1 0 22288 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_2
timestamp 1698431365
transform 1 0 1568 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_82
timestamp 1698431365
transform 1 0 10528 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_185
timestamp 1698431365
transform 1 0 22064 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_187
timestamp 1698431365
transform 1 0 22288 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_104
timestamp 1698431365
transform 1 0 12992 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_183
timestamp 1698431365
transform 1 0 21840 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_187
timestamp 1698431365
transform 1 0 22288 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_26
timestamp 1698431365
transform 1 0 4256 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_32
timestamp 1698431365
transform 1 0 4928 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_138
timestamp 1698431365
transform 1 0 16800 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_156
timestamp 1698431365
transform 1 0 18816 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_160
timestamp 1698431365
transform 1 0 19264 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_164
timestamp 1698431365
transform 1 0 19712 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_2
timestamp 1698431365
transform 1 0 1568 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_9
timestamp 1698431365
transform 1 0 2352 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_94
timestamp 1698431365
transform 1 0 11872 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_96
timestamp 1698431365
transform 1 0 12096 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_103
timestamp 1698431365
transform 1 0 12880 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_136
timestamp 1698431365
transform 1 0 16576 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_140
timestamp 1698431365
transform 1 0 17024 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_144 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17472 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_150
timestamp 1698431365
transform 1 0 18144 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_154
timestamp 1698431365
transform 1 0 18592 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_156
timestamp 1698431365
transform 1 0 18816 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_159
timestamp 1698431365
transform 1 0 19152 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_163
timestamp 1698431365
transform 1 0 19600 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_167
timestamp 1698431365
transform 1 0 20048 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_171
timestamp 1698431365
transform 1 0 20496 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_177
timestamp 1698431365
transform 1 0 21168 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_2
timestamp 1698431365
transform 1 0 1568 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_54
timestamp 1698431365
transform 1 0 7392 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_117
timestamp 1698431365
transform 1 0 14448 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_121
timestamp 1698431365
transform 1 0 14896 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_125 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 15344 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_133
timestamp 1698431365
transform 1 0 16240 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_137
timestamp 1698431365
transform 1 0 16688 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_139
timestamp 1698431365
transform 1 0 16912 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_142 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17248 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_158
timestamp 1698431365
transform 1 0 19040 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_168
timestamp 1698431365
transform 1 0 20160 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_172
timestamp 1698431365
transform 1 0 20608 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_174
timestamp 1698431365
transform 1 0 20832 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_177
timestamp 1698431365
transform 1 0 21168 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_181
timestamp 1698431365
transform 1 0 21616 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_185
timestamp 1698431365
transform 1 0 22064 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_18
timestamp 1698431365
transform 1 0 3360 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_28
timestamp 1698431365
transform 1 0 4480 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698431365
transform 1 0 5152 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_37
timestamp 1698431365
transform 1 0 5488 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_41
timestamp 1698431365
transform 1 0 5936 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_45
timestamp 1698431365
transform 1 0 6384 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_51
timestamp 1698431365
transform 1 0 7056 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_53
timestamp 1698431365
transform 1 0 7280 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_56
timestamp 1698431365
transform 1 0 7616 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_60
timestamp 1698431365
transform 1 0 8064 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_70
timestamp 1698431365
transform 1 0 9184 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_72
timestamp 1698431365
transform 1 0 9408 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_79
timestamp 1698431365
transform 1 0 10192 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_99
timestamp 1698431365
transform 1 0 12432 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_103
timestamp 1698431365
transform 1 0 12880 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_107 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13328 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_171
timestamp 1698431365
transform 1 0 20496 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_177
timestamp 1698431365
transform 1 0 21168 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_185
timestamp 1698431365
transform 1 0 22064 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_18
timestamp 1698431365
transform 1 0 3360 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_22
timestamp 1698431365
transform 1 0 3808 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_25
timestamp 1698431365
transform 1 0 4144 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_31
timestamp 1698431365
transform 1 0 4816 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_35
timestamp 1698431365
transform 1 0 5264 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_39
timestamp 1698431365
transform 1 0 5712 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_43
timestamp 1698431365
transform 1 0 6160 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_47
timestamp 1698431365
transform 1 0 6608 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_49
timestamp 1698431365
transform 1 0 6832 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_52
timestamp 1698431365
transform 1 0 7168 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_72
timestamp 1698431365
transform 1 0 9408 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_74
timestamp 1698431365
transform 1 0 9632 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_81
timestamp 1698431365
transform 1 0 10416 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_85
timestamp 1698431365
transform 1 0 10864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_89
timestamp 1698431365
transform 1 0 11312 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_93
timestamp 1698431365
transform 1 0 11760 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_9_97 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 12208 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_129
timestamp 1698431365
transform 1 0 15792 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_137
timestamp 1698431365
transform 1 0 16688 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_139
timestamp 1698431365
transform 1 0 16912 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_9_142
timestamp 1698431365
transform 1 0 17248 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_174
timestamp 1698431365
transform 1 0 20832 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_182
timestamp 1698431365
transform 1 0 21728 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_186
timestamp 1698431365
transform 1 0 22176 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_10
timestamp 1698431365
transform 1 0 2464 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_14
timestamp 1698431365
transform 1 0 2912 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_16
timestamp 1698431365
transform 1 0 3136 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_19
timestamp 1698431365
transform 1 0 3472 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_23
timestamp 1698431365
transform 1 0 3920 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_29
timestamp 1698431365
transform 1 0 4592 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_33
timestamp 1698431365
transform 1 0 5040 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_37
timestamp 1698431365
transform 1 0 5488 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_69
timestamp 1698431365
transform 1 0 9072 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_79
timestamp 1698431365
transform 1 0 10192 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_95
timestamp 1698431365
transform 1 0 11984 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_103
timestamp 1698431365
transform 1 0 12880 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_107
timestamp 1698431365
transform 1 0 13328 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_171
timestamp 1698431365
transform 1 0 20496 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_177
timestamp 1698431365
transform 1 0 21168 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_185
timestamp 1698431365
transform 1 0 22064 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_187
timestamp 1698431365
transform 1 0 22288 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_10
timestamp 1698431365
transform 1 0 2464 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_14
timestamp 1698431365
transform 1 0 2912 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_18
timestamp 1698431365
transform 1 0 3360 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_20
timestamp 1698431365
transform 1 0 3584 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_23
timestamp 1698431365
transform 1 0 3920 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_11_27
timestamp 1698431365
transform 1 0 4368 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_59
timestamp 1698431365
transform 1 0 7952 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_67
timestamp 1698431365
transform 1 0 8848 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_69
timestamp 1698431365
transform 1 0 9072 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_72
timestamp 1698431365
transform 1 0 9408 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_136
timestamp 1698431365
transform 1 0 16576 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_11_142
timestamp 1698431365
transform 1 0 17248 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_174
timestamp 1698431365
transform 1 0 20832 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_182
timestamp 1698431365
transform 1 0 21728 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_186
timestamp 1698431365
transform 1 0 22176 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_10
timestamp 1698431365
transform 1 0 2464 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_26
timestamp 1698431365
transform 1 0 4256 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698431365
transform 1 0 5152 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_37
timestamp 1698431365
transform 1 0 5488 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_101
timestamp 1698431365
transform 1 0 12656 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_107
timestamp 1698431365
transform 1 0 13328 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_171
timestamp 1698431365
transform 1 0 20496 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_177
timestamp 1698431365
transform 1 0 21168 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_179
timestamp 1698431365
transform 1 0 21392 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_6
timestamp 1698431365
transform 1 0 2016 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_72
timestamp 1698431365
transform 1 0 9408 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_136
timestamp 1698431365
transform 1 0 16576 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_142
timestamp 1698431365
transform 1 0 17248 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_174
timestamp 1698431365
transform 1 0 20832 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_182
timestamp 1698431365
transform 1 0 21728 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_186
timestamp 1698431365
transform 1 0 22176 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_10
timestamp 1698431365
transform 1 0 2464 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_26
timestamp 1698431365
transform 1 0 4256 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698431365
transform 1 0 5152 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_37
timestamp 1698431365
transform 1 0 5488 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_101
timestamp 1698431365
transform 1 0 12656 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_107
timestamp 1698431365
transform 1 0 13328 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_171
timestamp 1698431365
transform 1 0 20496 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_177
timestamp 1698431365
transform 1 0 21168 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_185
timestamp 1698431365
transform 1 0 22064 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_187
timestamp 1698431365
transform 1 0 22288 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_22
timestamp 1698431365
transform 1 0 3808 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_54
timestamp 1698431365
transform 1 0 7392 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_72
timestamp 1698431365
transform 1 0 9408 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_136
timestamp 1698431365
transform 1 0 16576 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_142
timestamp 1698431365
transform 1 0 17248 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_174
timestamp 1698431365
transform 1 0 20832 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_182
timestamp 1698431365
transform 1 0 21728 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_2
timestamp 1698431365
transform 1 0 1568 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_13
timestamp 1698431365
transform 1 0 2800 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_25
timestamp 1698431365
transform 1 0 4144 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_33
timestamp 1698431365
transform 1 0 5040 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_36
timestamp 1698431365
transform 1 0 5376 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_52
timestamp 1698431365
transform 1 0 7168 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_70
timestamp 1698431365
transform 1 0 9184 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_74
timestamp 1698431365
transform 1 0 9632 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_78
timestamp 1698431365
transform 1 0 10080 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_80
timestamp 1698431365
transform 1 0 10304 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_85
timestamp 1698431365
transform 1 0 10864 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_101
timestamp 1698431365
transform 1 0 12656 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_104
timestamp 1698431365
transform 1 0 12992 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_106
timestamp 1698431365
transform 1 0 13216 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_111
timestamp 1698431365
transform 1 0 13776 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_127
timestamp 1698431365
transform 1 0 15568 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_135
timestamp 1698431365
transform 1 0 16464 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_148
timestamp 1698431365
transform 1 0 17920 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_156
timestamp 1698431365
transform 1 0 18816 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_158
timestamp 1698431365
transform 1 0 19040 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_163
timestamp 1698431365
transform 1 0 19600 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_167
timestamp 1698431365
transform 1 0 20048 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_172
timestamp 1698431365
transform 1 0 20608 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_184
timestamp 1698431365
transform 1 0 21952 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input1 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 22400 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input2
timestamp 1698431365
transform -1 0 22400 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input3
timestamp 1698431365
transform -1 0 22064 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input4 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 3920 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input5
timestamp 1698431365
transform 1 0 3024 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input6
timestamp 1698431365
transform 1 0 9744 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input7
timestamp 1698431365
transform -1 0 11088 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input8
timestamp 1698431365
transform -1 0 11760 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input9
timestamp 1698431365
transform -1 0 12432 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input10
timestamp 1698431365
transform -1 0 12880 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input11
timestamp 1698431365
transform 1 0 3024 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input12
timestamp 1698431365
transform -1 0 16016 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input13
timestamp 1698431365
transform -1 0 21280 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input14
timestamp 1698431365
transform 1 0 3696 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input15
timestamp 1698431365
transform 1 0 1680 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input16
timestamp 1698431365
transform -1 0 19264 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input17
timestamp 1698431365
transform -1 0 17024 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input18
timestamp 1698431365
transform -1 0 19936 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input19
timestamp 1698431365
transform -1 0 21952 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input20
timestamp 1698431365
transform 1 0 18144 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input21
timestamp 1698431365
transform 1 0 19936 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input22
timestamp 1698431365
transform -1 0 21952 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input23
timestamp 1698431365
transform -1 0 19600 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input24
timestamp 1698431365
transform -1 0 20272 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input25
timestamp 1698431365
transform -1 0 21728 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input26
timestamp 1698431365
transform 1 0 2352 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input27
timestamp 1698431365
transform 1 0 20272 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input28
timestamp 1698431365
transform 1 0 19936 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input29
timestamp 1698431365
transform 1 0 3696 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input30
timestamp 1698431365
transform 1 0 5488 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input31
timestamp 1698431365
transform 1 0 7616 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input32
timestamp 1698431365
transform 1 0 6160 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input33
timestamp 1698431365
transform 1 0 3584 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input34
timestamp 1698431365
transform 1 0 8512 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input35
timestamp 1698431365
transform 1 0 9520 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input36
timestamp 1698431365
transform 1 0 2240 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input37
timestamp 1698431365
transform 1 0 1568 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input38
timestamp 1698431365
transform 1 0 4592 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input39
timestamp 1698431365
transform 1 0 2576 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input40
timestamp 1698431365
transform 1 0 3248 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input41
timestamp 1698431365
transform 1 0 21168 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output42 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 17920 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output43
timestamp 1698431365
transform 1 0 20832 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output44
timestamp 1698431365
transform -1 0 2688 0 1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output45
timestamp 1698431365
transform -1 0 4032 0 1 3136
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output46
timestamp 1698431365
transform -1 0 2912 0 1 3136
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output47
timestamp 1698431365
transform -1 0 2800 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output48 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 8960 0 1 15680
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_17 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698431365
transform -1 0 22624 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_18
timestamp 1698431365
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698431365
transform -1 0 22624 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_19
timestamp 1698431365
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698431365
transform -1 0 22624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_20
timestamp 1698431365
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698431365
transform -1 0 22624 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_21
timestamp 1698431365
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698431365
transform -1 0 22624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_22
timestamp 1698431365
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698431365
transform -1 0 22624 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_23
timestamp 1698431365
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698431365
transform -1 0 22624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_24
timestamp 1698431365
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698431365
transform -1 0 22624 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_25
timestamp 1698431365
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698431365
transform -1 0 22624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_26
timestamp 1698431365
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698431365
transform -1 0 22624 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_27
timestamp 1698431365
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698431365
transform -1 0 22624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_28
timestamp 1698431365
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698431365
transform -1 0 22624 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_29
timestamp 1698431365
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698431365
transform -1 0 22624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_30
timestamp 1698431365
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698431365
transform -1 0 22624 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_31
timestamp 1698431365
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698431365
transform -1 0 22624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_32
timestamp 1698431365
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698431365
transform -1 0 22624 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_33
timestamp 1698431365
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698431365
transform -1 0 22624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_34 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_35
timestamp 1698431365
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_36
timestamp 1698431365
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_37
timestamp 1698431365
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_38
timestamp 1698431365
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_39
timestamp 1698431365
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_40
timestamp 1698431365
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_41
timestamp 1698431365
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_42
timestamp 1698431365
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_43
timestamp 1698431365
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_44
timestamp 1698431365
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_45
timestamp 1698431365
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_46
timestamp 1698431365
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_47
timestamp 1698431365
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_48
timestamp 1698431365
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_49
timestamp 1698431365
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_50
timestamp 1698431365
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_51
timestamp 1698431365
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_52
timestamp 1698431365
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_53
timestamp 1698431365
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_54
timestamp 1698431365
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_55
timestamp 1698431365
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_56
timestamp 1698431365
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_57
timestamp 1698431365
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_58
timestamp 1698431365
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_59
timestamp 1698431365
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_60
timestamp 1698431365
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_61
timestamp 1698431365
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_62
timestamp 1698431365
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_63
timestamp 1698431365
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_64
timestamp 1698431365
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_65
timestamp 1698431365
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_66
timestamp 1698431365
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_67
timestamp 1698431365
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_68
timestamp 1698431365
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_69
timestamp 1698431365
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_70
timestamp 1698431365
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_71
timestamp 1698431365
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_72
timestamp 1698431365
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_73
timestamp 1698431365
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_74
timestamp 1698431365
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_75
timestamp 1698431365
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_76
timestamp 1698431365
transform 1 0 5152 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_77
timestamp 1698431365
transform 1 0 8960 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_78
timestamp 1698431365
transform 1 0 12768 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_79
timestamp 1698431365
transform 1 0 16576 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_80
timestamp 1698431365
transform 1 0 20384 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_49 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 21952 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_50
timestamp 1698431365
transform -1 0 13776 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_51
timestamp 1698431365
transform -1 0 19600 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_52
timestamp 1698431365
transform -1 0 2464 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_53
timestamp 1698431365
transform -1 0 2912 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_54
timestamp 1698431365
transform -1 0 3024 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_55
timestamp 1698431365
transform -1 0 2576 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_56
timestamp 1698431365
transform -1 0 2016 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_57
timestamp 1698431365
transform -1 0 4928 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_58
timestamp 1698431365
transform -1 0 4480 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_59
timestamp 1698431365
transform -1 0 4032 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_60
timestamp 1698431365
transform -1 0 3360 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_61
timestamp 1698431365
transform -1 0 2128 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_62
timestamp 1698431365
transform -1 0 2912 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_63
timestamp 1698431365
transform -1 0 2464 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_64
timestamp 1698431365
transform -1 0 2016 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_65
timestamp 1698431365
transform -1 0 2016 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_66
timestamp 1698431365
transform -1 0 2464 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_67
timestamp 1698431365
transform -1 0 2016 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_68
timestamp 1698431365
transform -1 0 2464 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_69
timestamp 1698431365
transform -1 0 2016 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_70
timestamp 1698431365
transform -1 0 2464 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_71
timestamp 1698431365
transform -1 0 2016 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_72
timestamp 1698431365
transform -1 0 2016 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_73
timestamp 1698431365
transform -1 0 2016 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_74
timestamp 1698431365
transform -1 0 2464 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_75
timestamp 1698431365
transform -1 0 2016 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_76
timestamp 1698431365
transform -1 0 2464 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_77
timestamp 1698431365
transform -1 0 3696 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_78
timestamp 1698431365
transform -1 0 2912 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_79
timestamp 1698431365
transform -1 0 3360 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_80
timestamp 1698431365
transform -1 0 4144 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_81
timestamp 1698431365
transform -1 0 3808 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_82
timestamp 1698431365
transform -1 0 3360 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_83
timestamp 1698431365
transform -1 0 5040 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_84
timestamp 1698431365
transform -1 0 10864 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  wb_buttons_leds_85 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 21952 0 -1 15680
box -86 -86 534 870
<< labels >>
flabel metal3 s 23200 2464 24000 2576 0 FreeSans 448 0 0 0 buttons[0]
port 0 nsew signal input
flabel metal3 s 23200 12320 24000 12432 0 FreeSans 448 0 0 0 buttons[1]
port 1 nsew signal input
flabel metal3 s 23200 17248 24000 17360 0 FreeSans 448 0 0 0 buttons_enb[0]
port 2 nsew signal tristate
flabel metal3 s 23200 7392 24000 7504 0 FreeSans 448 0 0 0 buttons_enb[1]
port 3 nsew signal tristate
flabel metal2 s 19712 0 19824 800 0 FreeSans 448 90 0 0 clk
port 4 nsew signal input
flabel metal2 s 20160 0 20272 800 0 FreeSans 448 90 0 0 clk2
port 5 nsew signal input
flabel metal2 s 4480 0 4592 800 0 FreeSans 448 90 0 0 i_wb_addr[0]
port 6 nsew signal input
flabel metal2 s 9856 0 9968 800 0 FreeSans 448 90 0 0 i_wb_addr[10]
port 7 nsew signal input
flabel metal2 s 10304 0 10416 800 0 FreeSans 448 90 0 0 i_wb_addr[11]
port 8 nsew signal input
flabel metal2 s 10752 0 10864 800 0 FreeSans 448 90 0 0 i_wb_addr[12]
port 9 nsew signal input
flabel metal2 s 11200 0 11312 800 0 FreeSans 448 90 0 0 i_wb_addr[13]
port 10 nsew signal input
flabel metal2 s 11648 0 11760 800 0 FreeSans 448 90 0 0 i_wb_addr[14]
port 11 nsew signal input
flabel metal2 s 12096 0 12208 800 0 FreeSans 448 90 0 0 i_wb_addr[15]
port 12 nsew signal input
flabel metal2 s 12544 0 12656 800 0 FreeSans 448 90 0 0 i_wb_addr[16]
port 13 nsew signal input
flabel metal2 s 12992 0 13104 800 0 FreeSans 448 90 0 0 i_wb_addr[17]
port 14 nsew signal input
flabel metal2 s 13440 0 13552 800 0 FreeSans 448 90 0 0 i_wb_addr[18]
port 15 nsew signal input
flabel metal2 s 13888 0 14000 800 0 FreeSans 448 90 0 0 i_wb_addr[19]
port 16 nsew signal input
flabel metal2 s 5376 0 5488 800 0 FreeSans 448 90 0 0 i_wb_addr[1]
port 17 nsew signal input
flabel metal2 s 14336 0 14448 800 0 FreeSans 448 90 0 0 i_wb_addr[20]
port 18 nsew signal input
flabel metal2 s 14784 0 14896 800 0 FreeSans 448 90 0 0 i_wb_addr[21]
port 19 nsew signal input
flabel metal2 s 15232 0 15344 800 0 FreeSans 448 90 0 0 i_wb_addr[22]
port 20 nsew signal input
flabel metal2 s 15680 0 15792 800 0 FreeSans 448 90 0 0 i_wb_addr[23]
port 21 nsew signal input
flabel metal2 s 16128 0 16240 800 0 FreeSans 448 90 0 0 i_wb_addr[24]
port 22 nsew signal input
flabel metal2 s 16576 0 16688 800 0 FreeSans 448 90 0 0 i_wb_addr[25]
port 23 nsew signal input
flabel metal2 s 17024 0 17136 800 0 FreeSans 448 90 0 0 i_wb_addr[26]
port 24 nsew signal input
flabel metal2 s 17472 0 17584 800 0 FreeSans 448 90 0 0 i_wb_addr[27]
port 25 nsew signal input
flabel metal2 s 17920 0 18032 800 0 FreeSans 448 90 0 0 i_wb_addr[28]
port 26 nsew signal input
flabel metal2 s 18368 0 18480 800 0 FreeSans 448 90 0 0 i_wb_addr[29]
port 27 nsew signal input
flabel metal2 s 6272 0 6384 800 0 FreeSans 448 90 0 0 i_wb_addr[2]
port 28 nsew signal input
flabel metal2 s 18816 0 18928 800 0 FreeSans 448 90 0 0 i_wb_addr[30]
port 29 nsew signal input
flabel metal2 s 19264 0 19376 800 0 FreeSans 448 90 0 0 i_wb_addr[31]
port 30 nsew signal input
flabel metal2 s 6720 0 6832 800 0 FreeSans 448 90 0 0 i_wb_addr[3]
port 31 nsew signal input
flabel metal2 s 7168 0 7280 800 0 FreeSans 448 90 0 0 i_wb_addr[4]
port 32 nsew signal input
flabel metal2 s 7616 0 7728 800 0 FreeSans 448 90 0 0 i_wb_addr[5]
port 33 nsew signal input
flabel metal2 s 8064 0 8176 800 0 FreeSans 448 90 0 0 i_wb_addr[6]
port 34 nsew signal input
flabel metal2 s 8512 0 8624 800 0 FreeSans 448 90 0 0 i_wb_addr[7]
port 35 nsew signal input
flabel metal2 s 8960 0 9072 800 0 FreeSans 448 90 0 0 i_wb_addr[8]
port 36 nsew signal input
flabel metal2 s 9408 0 9520 800 0 FreeSans 448 90 0 0 i_wb_addr[9]
port 37 nsew signal input
flabel metal2 s 3136 0 3248 800 0 FreeSans 448 90 0 0 i_wb_cyc
port 38 nsew signal input
flabel metal2 s 4928 0 5040 800 0 FreeSans 448 90 0 0 i_wb_data[0]
port 39 nsew signal input
flabel metal2 s 5824 0 5936 800 0 FreeSans 448 90 0 0 i_wb_data[1]
port 40 nsew signal input
flabel metal2 s 3584 0 3696 800 0 FreeSans 448 90 0 0 i_wb_stb
port 41 nsew signal input
flabel metal2 s 4032 0 4144 800 0 FreeSans 448 90 0 0 i_wb_we
port 42 nsew signal input
flabel metal2 s 13216 19200 13328 20000 0 FreeSans 448 90 0 0 led_enb[0]
port 43 nsew signal tristate
flabel metal2 s 19040 19200 19152 20000 0 FreeSans 448 90 0 0 led_enb[1]
port 44 nsew signal tristate
flabel metal2 s 16128 19200 16240 20000 0 FreeSans 448 90 0 0 leds[0]
port 45 nsew signal tristate
flabel metal2 s 21952 19200 22064 20000 0 FreeSans 448 90 0 0 leds[1]
port 46 nsew signal tristate
flabel metal3 s 0 2464 800 2576 0 FreeSans 448 0 0 0 o_wb_ack
port 47 nsew signal tristate
flabel metal3 s 0 3360 800 3472 0 FreeSans 448 0 0 0 o_wb_data[0]
port 48 nsew signal tristate
flabel metal3 s 0 7840 800 7952 0 FreeSans 448 0 0 0 o_wb_data[10]
port 49 nsew signal tristate
flabel metal3 s 0 8288 800 8400 0 FreeSans 448 0 0 0 o_wb_data[11]
port 50 nsew signal tristate
flabel metal3 s 0 8736 800 8848 0 FreeSans 448 0 0 0 o_wb_data[12]
port 51 nsew signal tristate
flabel metal3 s 0 9184 800 9296 0 FreeSans 448 0 0 0 o_wb_data[13]
port 52 nsew signal tristate
flabel metal3 s 0 9632 800 9744 0 FreeSans 448 0 0 0 o_wb_data[14]
port 53 nsew signal tristate
flabel metal3 s 0 10080 800 10192 0 FreeSans 448 0 0 0 o_wb_data[15]
port 54 nsew signal tristate
flabel metal3 s 0 10528 800 10640 0 FreeSans 448 0 0 0 o_wb_data[16]
port 55 nsew signal tristate
flabel metal3 s 0 10976 800 11088 0 FreeSans 448 0 0 0 o_wb_data[17]
port 56 nsew signal tristate
flabel metal3 s 0 11424 800 11536 0 FreeSans 448 0 0 0 o_wb_data[18]
port 57 nsew signal tristate
flabel metal3 s 0 11872 800 11984 0 FreeSans 448 0 0 0 o_wb_data[19]
port 58 nsew signal tristate
flabel metal3 s 0 3808 800 3920 0 FreeSans 448 0 0 0 o_wb_data[1]
port 59 nsew signal tristate
flabel metal3 s 0 12320 800 12432 0 FreeSans 448 0 0 0 o_wb_data[20]
port 60 nsew signal tristate
flabel metal3 s 0 12768 800 12880 0 FreeSans 448 0 0 0 o_wb_data[21]
port 61 nsew signal tristate
flabel metal3 s 0 13216 800 13328 0 FreeSans 448 0 0 0 o_wb_data[22]
port 62 nsew signal tristate
flabel metal3 s 0 13664 800 13776 0 FreeSans 448 0 0 0 o_wb_data[23]
port 63 nsew signal tristate
flabel metal3 s 0 14112 800 14224 0 FreeSans 448 0 0 0 o_wb_data[24]
port 64 nsew signal tristate
flabel metal3 s 0 14560 800 14672 0 FreeSans 448 0 0 0 o_wb_data[25]
port 65 nsew signal tristate
flabel metal3 s 0 15008 800 15120 0 FreeSans 448 0 0 0 o_wb_data[26]
port 66 nsew signal tristate
flabel metal3 s 0 15456 800 15568 0 FreeSans 448 0 0 0 o_wb_data[27]
port 67 nsew signal tristate
flabel metal3 s 0 15904 800 16016 0 FreeSans 448 0 0 0 o_wb_data[28]
port 68 nsew signal tristate
flabel metal3 s 0 16352 800 16464 0 FreeSans 448 0 0 0 o_wb_data[29]
port 69 nsew signal tristate
flabel metal3 s 0 4256 800 4368 0 FreeSans 448 0 0 0 o_wb_data[2]
port 70 nsew signal tristate
flabel metal3 s 0 16800 800 16912 0 FreeSans 448 0 0 0 o_wb_data[30]
port 71 nsew signal tristate
flabel metal3 s 0 17248 800 17360 0 FreeSans 448 0 0 0 o_wb_data[31]
port 72 nsew signal tristate
flabel metal3 s 0 4704 800 4816 0 FreeSans 448 0 0 0 o_wb_data[3]
port 73 nsew signal tristate
flabel metal3 s 0 5152 800 5264 0 FreeSans 448 0 0 0 o_wb_data[4]
port 74 nsew signal tristate
flabel metal3 s 0 5600 800 5712 0 FreeSans 448 0 0 0 o_wb_data[5]
port 75 nsew signal tristate
flabel metal3 s 0 6048 800 6160 0 FreeSans 448 0 0 0 o_wb_data[6]
port 76 nsew signal tristate
flabel metal3 s 0 6496 800 6608 0 FreeSans 448 0 0 0 o_wb_data[7]
port 77 nsew signal tristate
flabel metal3 s 0 6944 800 7056 0 FreeSans 448 0 0 0 o_wb_data[8]
port 78 nsew signal tristate
flabel metal3 s 0 7392 800 7504 0 FreeSans 448 0 0 0 o_wb_data[9]
port 79 nsew signal tristate
flabel metal3 s 0 2912 800 3024 0 FreeSans 448 0 0 0 o_wb_stall
port 80 nsew signal tristate
flabel metal2 s 20608 0 20720 800 0 FreeSans 448 90 0 0 reset
port 81 nsew signal input
flabel metal4 s 3844 3076 4164 16524 0 FreeSans 1280 90 0 0 vdd
port 82 nsew power bidirectional
flabel metal4 s 9164 3076 9484 16524 0 FreeSans 1280 90 0 0 vdd
port 82 nsew power bidirectional
flabel metal4 s 14484 3076 14804 16524 0 FreeSans 1280 90 0 0 vdd
port 82 nsew power bidirectional
flabel metal4 s 19804 3076 20124 16524 0 FreeSans 1280 90 0 0 vdd
port 82 nsew power bidirectional
flabel metal4 s 6504 3076 6824 16524 0 FreeSans 1280 90 0 0 vss
port 83 nsew ground bidirectional
flabel metal4 s 11824 3076 12144 16524 0 FreeSans 1280 90 0 0 vss
port 83 nsew ground bidirectional
flabel metal4 s 17144 3076 17464 16524 0 FreeSans 1280 90 0 0 vss
port 83 nsew ground bidirectional
flabel metal4 s 22464 3076 22784 16524 0 FreeSans 1280 90 0 0 vss
port 83 nsew ground bidirectional
flabel metal2 s 4480 19200 4592 20000 0 FreeSans 448 90 0 0 xtal_clk[0]
port 84 nsew signal tristate
flabel metal2 s 10304 19200 10416 20000 0 FreeSans 448 90 0 0 xtal_clk[1]
port 85 nsew signal tristate
flabel metal2 s 1568 19200 1680 20000 0 FreeSans 448 90 0 0 xtal_clk_enb[0]
port 86 nsew signal tristate
flabel metal2 s 7392 19200 7504 20000 0 FreeSans 448 90 0 0 xtal_clk_enb[1]
port 87 nsew signal tristate
rlabel metal1 11984 16464 11984 16464 0 vdd
rlabel via1 12064 15680 12064 15680 0 vss
rlabel metal2 20440 6048 20440 6048 0 _000_
rlabel metal2 2856 5096 2856 5096 0 _001_
rlabel metal2 4984 6888 4984 6888 0 _002_
rlabel metal2 8064 5208 8064 5208 0 _003_
rlabel metal3 16688 7336 16688 7336 0 _004_
rlabel metal2 14224 8344 14224 8344 0 _005_
rlabel metal2 16184 4256 16184 4256 0 _006_
rlabel metal2 17416 6776 17416 6776 0 _007_
rlabel metal3 6496 3752 6496 3752 0 _008_
rlabel metal2 22008 5040 22008 5040 0 _009_
rlabel metal2 16744 6832 16744 6832 0 _010_
rlabel metal2 10920 3920 10920 3920 0 _011_
rlabel metal2 11368 6608 11368 6608 0 _012_
rlabel metal2 10696 4312 10696 4312 0 _013_
rlabel metal3 11200 7560 11200 7560 0 _014_
rlabel metal2 14952 4200 14952 4200 0 _015_
rlabel metal2 14168 3808 14168 3808 0 _016_
rlabel via2 13384 4984 13384 4984 0 _017_
rlabel metal2 19208 4368 19208 4368 0 _018_
rlabel metal2 19320 3808 19320 3808 0 _019_
rlabel metal2 12768 5096 12768 5096 0 _020_
rlabel metal2 5656 6496 5656 6496 0 _021_
rlabel metal3 9128 3416 9128 3416 0 _022_
rlabel metal2 6048 6664 6048 6664 0 _023_
rlabel metal2 1960 5656 1960 5656 0 _024_
rlabel metal2 6888 8904 6888 8904 0 _025_
rlabel metal3 2772 5768 2772 5768 0 _026_
rlabel metal2 2184 6104 2184 6104 0 _027_
rlabel metal2 3304 8176 3304 8176 0 _028_
rlabel metal2 4536 5600 4536 5600 0 _029_
rlabel metal2 4872 6216 4872 6216 0 _030_
rlabel metal2 4816 3640 4816 3640 0 _031_
rlabel metal2 13272 4480 13272 4480 0 _032_
rlabel metal2 10584 4144 10584 4144 0 _033_
rlabel metal2 4648 5152 4648 5152 0 _034_
rlabel metal2 8792 7560 8792 7560 0 _035_
rlabel metal2 9464 4928 9464 4928 0 _036_
rlabel metal2 7112 8624 7112 8624 0 _037_
rlabel metal3 7896 3304 7896 3304 0 _038_
rlabel metal2 17304 6944 17304 6944 0 _039_
rlabel metal2 17528 6272 17528 6272 0 _040_
rlabel metal2 13608 7112 13608 7112 0 _041_
rlabel metal3 22778 2520 22778 2520 0 buttons[0]
rlabel metal2 22232 12600 22232 12600 0 buttons[1]
rlabel metal2 19768 2058 19768 2058 0 clk
rlabel metal1 21000 2968 21000 2968 0 clk2
rlabel metal2 13496 6328 13496 6328 0 clknet_0_clk
rlabel metal2 5096 6776 5096 6776 0 clknet_1_0__leaf_clk
rlabel metal2 16520 7112 16520 7112 0 clknet_1_1__leaf_clk
rlabel metal2 4480 3304 4480 3304 0 i_wb_addr[0]
rlabel metal2 9912 1470 9912 1470 0 i_wb_addr[10]
rlabel metal2 10360 2030 10360 2030 0 i_wb_addr[11]
rlabel metal2 11032 10584 11032 10584 0 i_wb_addr[12]
rlabel metal2 11256 2058 11256 2058 0 i_wb_addr[13]
rlabel metal2 11704 5614 11704 5614 0 i_wb_addr[14]
rlabel metal2 12544 8232 12544 8232 0 i_wb_addr[15]
rlabel metal2 3864 12096 3864 12096 0 i_wb_addr[16]
rlabel metal2 15736 4088 15736 4088 0 i_wb_addr[17]
rlabel metal2 13496 1302 13496 1302 0 i_wb_addr[18]
rlabel metal2 3976 4648 3976 4648 0 i_wb_addr[19]
rlabel metal2 1848 7952 1848 7952 0 i_wb_addr[1]
rlabel metal2 19096 4760 19096 4760 0 i_wb_addr[20]
rlabel metal2 14952 3304 14952 3304 0 i_wb_addr[21]
rlabel metal3 19712 5096 19712 5096 0 i_wb_addr[22]
rlabel metal2 15792 3192 15792 3192 0 i_wb_addr[23]
rlabel metal2 16352 3192 16352 3192 0 i_wb_addr[24]
rlabel metal2 20104 5208 20104 5208 0 i_wb_addr[25]
rlabel metal2 17080 2030 17080 2030 0 i_wb_addr[26]
rlabel metal2 17528 2058 17528 2058 0 i_wb_addr[27]
rlabel metal2 19992 6328 19992 6328 0 i_wb_addr[28]
rlabel metal2 18424 1582 18424 1582 0 i_wb_addr[29]
rlabel metal2 6216 3192 6216 3192 0 i_wb_addr[2]
rlabel metal3 19656 6552 19656 6552 0 i_wb_addr[30]
rlabel metal2 19152 3192 19152 3192 0 i_wb_addr[31]
rlabel metal2 6832 2968 6832 2968 0 i_wb_addr[3]
rlabel metal2 5768 8176 5768 8176 0 i_wb_addr[4]
rlabel metal2 7728 9016 7728 9016 0 i_wb_addr[5]
rlabel metal2 6328 7952 6328 7952 0 i_wb_addr[6]
rlabel metal3 5936 7448 5936 7448 0 i_wb_addr[7]
rlabel metal2 9016 2058 9016 2058 0 i_wb_addr[8]
rlabel metal2 9464 2058 9464 2058 0 i_wb_addr[9]
rlabel metal2 2464 7448 2464 7448 0 i_wb_cyc
rlabel metal2 2744 12040 2744 12040 0 i_wb_data[0]
rlabel metal2 5712 3192 5712 3192 0 i_wb_data[1]
rlabel metal2 3640 2058 3640 2058 0 i_wb_stb
rlabel metal2 3528 7560 3528 7560 0 i_wb_we
rlabel metal2 17080 16240 17080 16240 0 leds[0]
rlabel metal2 21896 16296 21896 16296 0 leds[1]
rlabel metal2 22064 5208 22064 5208 0 net1
rlabel metal2 7336 5208 7336 5208 0 net10
rlabel metal2 3528 4592 3528 4592 0 net11
rlabel metal2 15512 3920 15512 3920 0 net12
rlabel metal2 16744 3920 16744 3920 0 net13
rlabel metal2 15176 4032 15176 4032 0 net14
rlabel metal2 2184 7672 2184 7672 0 net15
rlabel metal2 16408 5152 16408 5152 0 net16
rlabel metal2 15848 5544 15848 5544 0 net17
rlabel metal2 18424 5040 18424 5040 0 net18
rlabel metal2 16856 4704 16856 4704 0 net19
rlabel metal2 20944 7560 20944 7560 0 net2
rlabel metal2 18648 7336 18648 7336 0 net20
rlabel metal2 20440 5152 20440 5152 0 net21
rlabel metal2 21056 4424 21056 4424 0 net22
rlabel metal2 19096 5936 19096 5936 0 net23
rlabel metal2 16968 5152 16968 5152 0 net24
rlabel metal2 18424 4088 18424 4088 0 net25
rlabel metal2 6272 5992 6272 5992 0 net26
rlabel metal3 21056 5096 21056 5096 0 net27
rlabel metal2 21560 5376 21560 5376 0 net28
rlabel metal2 6888 5488 6888 5488 0 net29
rlabel metal2 21224 5936 21224 5936 0 net3
rlabel metal2 5992 8176 5992 8176 0 net30
rlabel metal2 8232 9128 8232 9128 0 net31
rlabel metal3 7336 8120 7336 8120 0 net32
rlabel metal2 4088 7840 4088 7840 0 net33
rlabel metal2 9072 9576 9072 9576 0 net34
rlabel metal2 10024 9352 10024 9352 0 net35
rlabel metal3 4984 9576 4984 9576 0 net36
rlabel metal2 2072 8400 2072 8400 0 net37
rlabel metal2 16296 4312 16296 4312 0 net38
rlabel metal2 3080 7840 3080 7840 0 net39
rlabel metal2 7224 6440 7224 6440 0 net4
rlabel metal3 7168 5992 7168 5992 0 net40
rlabel metal2 21672 5376 21672 5376 0 net41
rlabel metal2 17752 13804 17752 13804 0 net42
rlabel metal2 20664 15848 20664 15848 0 net43
rlabel metal2 1960 4648 1960 4648 0 net44
rlabel metal2 3752 8568 3752 8568 0 net45
rlabel metal2 5880 5152 5880 5152 0 net46
rlabel metal2 2688 15848 2688 15848 0 net47
rlabel metal3 12712 15848 12712 15848 0 net48
rlabel metal2 22288 8008 22288 8008 0 net49
rlabel metal2 3528 6384 3528 6384 0 net5
rlabel metal2 13384 15960 13384 15960 0 net50
rlabel metal2 19208 15960 19208 15960 0 net51
rlabel metal3 1134 4312 1134 4312 0 net52
rlabel metal3 1302 4760 1302 4760 0 net53
rlabel metal3 1750 5208 1750 5208 0 net54
rlabel metal3 1358 5656 1358 5656 0 net55
rlabel metal3 1246 6104 1246 6104 0 net56
rlabel metal2 4648 7056 4648 7056 0 net57
rlabel metal3 1414 7000 1414 7000 0 net58
rlabel metal3 3528 7560 3528 7560 0 net59
rlabel metal2 10248 10528 10248 10528 0 net6
rlabel metal3 1134 7896 1134 7896 0 net60
rlabel metal3 1302 8344 1302 8344 0 net61
rlabel metal3 1638 8792 1638 8792 0 net62
rlabel metal3 1470 9240 1470 9240 0 net63
rlabel metal3 1736 9632 1736 9632 0 net64
rlabel metal3 1246 10136 1246 10136 0 net65
rlabel metal3 1414 10584 1414 10584 0 net66
rlabel metal3 1246 11032 1246 11032 0 net67
rlabel metal3 1470 11480 1470 11480 0 net68
rlabel metal3 1246 11928 1246 11928 0 net69
rlabel metal2 7000 4536 7000 4536 0 net7
rlabel metal3 1470 12376 1470 12376 0 net70
rlabel metal3 1246 12824 1246 12824 0 net71
rlabel metal3 1246 13272 1246 13272 0 net72
rlabel metal3 1246 13720 1246 13720 0 net73
rlabel metal3 1470 14168 1470 14168 0 net74
rlabel metal3 1246 14616 1246 14616 0 net75
rlabel metal3 1470 15064 1470 15064 0 net76
rlabel metal3 2086 15512 2086 15512 0 net77
rlabel metal2 2576 15512 2576 15512 0 net78
rlabel metal2 3080 15960 3080 15960 0 net79
rlabel metal2 11256 9408 11256 9408 0 net8
rlabel metal2 3808 15960 3808 15960 0 net80
rlabel metal2 3528 16408 3528 16408 0 net81
rlabel metal3 1638 2968 1638 2968 0 net82
rlabel metal2 4648 15960 4648 15960 0 net83
rlabel metal2 10472 15960 10472 15960 0 net84
rlabel metal3 22722 17304 22722 17304 0 net85
rlabel metal2 9016 4704 9016 4704 0 net9
rlabel metal3 1246 2520 1246 2520 0 o_wb_ack
rlabel metal3 1918 3416 1918 3416 0 o_wb_data[0]
rlabel metal3 1358 3864 1358 3864 0 o_wb_data[1]
rlabel metal2 21336 6496 21336 6496 0 reset
rlabel metal2 1736 16296 1736 16296 0 xtal_clk_enb[0]
rlabel metal2 7784 16912 7784 16912 0 xtal_clk_enb[1]
<< properties >>
string FIXED_BBOX 0 0 24000 20000
<< end >>
