magic
tech gf180mcuD
magscale 1 5
timestamp 1700704991
<< obsm1 >>
rect 672 1538 89320 98422
<< metal2 >>
rect 1904 99600 1960 100000
rect 5488 99600 5544 100000
rect 9072 99600 9128 100000
rect 12656 99600 12712 100000
rect 16240 99600 16296 100000
rect 19824 99600 19880 100000
rect 23408 99600 23464 100000
rect 26992 99600 27048 100000
rect 30576 99600 30632 100000
rect 34160 99600 34216 100000
rect 37744 99600 37800 100000
rect 41328 99600 41384 100000
rect 44912 99600 44968 100000
rect 48496 99600 48552 100000
rect 52080 99600 52136 100000
rect 55664 99600 55720 100000
rect 59248 99600 59304 100000
rect 62832 99600 62888 100000
rect 66416 99600 66472 100000
rect 70000 99600 70056 100000
rect 73584 99600 73640 100000
rect 77168 99600 77224 100000
rect 80752 99600 80808 100000
rect 84336 99600 84392 100000
rect 87920 99600 87976 100000
rect 4592 0 4648 400
rect 5488 0 5544 400
rect 6384 0 6440 400
rect 7280 0 7336 400
rect 8176 0 8232 400
rect 9072 0 9128 400
rect 9968 0 10024 400
rect 10864 0 10920 400
rect 11760 0 11816 400
rect 12656 0 12712 400
rect 13552 0 13608 400
rect 14448 0 14504 400
rect 15344 0 15400 400
rect 16240 0 16296 400
rect 17136 0 17192 400
rect 18032 0 18088 400
rect 18928 0 18984 400
rect 19824 0 19880 400
rect 20720 0 20776 400
rect 21616 0 21672 400
rect 22512 0 22568 400
rect 23408 0 23464 400
rect 24304 0 24360 400
rect 25200 0 25256 400
rect 26096 0 26152 400
rect 26992 0 27048 400
rect 27888 0 27944 400
rect 28784 0 28840 400
rect 29680 0 29736 400
rect 30576 0 30632 400
rect 31472 0 31528 400
rect 32368 0 32424 400
rect 33264 0 33320 400
rect 34160 0 34216 400
rect 35056 0 35112 400
rect 35952 0 36008 400
rect 36848 0 36904 400
rect 37744 0 37800 400
rect 38640 0 38696 400
rect 39536 0 39592 400
rect 40432 0 40488 400
rect 41328 0 41384 400
rect 42224 0 42280 400
rect 43120 0 43176 400
rect 44016 0 44072 400
rect 44912 0 44968 400
rect 45808 0 45864 400
rect 46704 0 46760 400
rect 47600 0 47656 400
rect 48496 0 48552 400
rect 49392 0 49448 400
rect 50288 0 50344 400
rect 51184 0 51240 400
rect 52080 0 52136 400
rect 52976 0 53032 400
rect 53872 0 53928 400
rect 54768 0 54824 400
rect 55664 0 55720 400
rect 56560 0 56616 400
rect 57456 0 57512 400
rect 58352 0 58408 400
rect 59248 0 59304 400
rect 60144 0 60200 400
rect 61040 0 61096 400
rect 61936 0 61992 400
rect 62832 0 62888 400
rect 63728 0 63784 400
rect 64624 0 64680 400
rect 65520 0 65576 400
rect 66416 0 66472 400
rect 67312 0 67368 400
rect 68208 0 68264 400
rect 69104 0 69160 400
rect 70000 0 70056 400
rect 70896 0 70952 400
rect 71792 0 71848 400
rect 72688 0 72744 400
rect 73584 0 73640 400
rect 74480 0 74536 400
rect 75376 0 75432 400
rect 76272 0 76328 400
rect 77168 0 77224 400
rect 78064 0 78120 400
rect 78960 0 79016 400
rect 79856 0 79912 400
rect 80752 0 80808 400
rect 81648 0 81704 400
rect 82544 0 82600 400
rect 83440 0 83496 400
rect 84336 0 84392 400
rect 85232 0 85288 400
<< obsm2 >>
rect 854 99570 1874 99666
rect 1990 99570 5458 99666
rect 5574 99570 9042 99666
rect 9158 99570 12626 99666
rect 12742 99570 16210 99666
rect 16326 99570 19794 99666
rect 19910 99570 23378 99666
rect 23494 99570 26962 99666
rect 27078 99570 30546 99666
rect 30662 99570 34130 99666
rect 34246 99570 37714 99666
rect 37830 99570 41298 99666
rect 41414 99570 44882 99666
rect 44998 99570 48466 99666
rect 48582 99570 52050 99666
rect 52166 99570 55634 99666
rect 55750 99570 59218 99666
rect 59334 99570 62802 99666
rect 62918 99570 66386 99666
rect 66502 99570 69970 99666
rect 70086 99570 73554 99666
rect 73670 99570 77138 99666
rect 77254 99570 80722 99666
rect 80838 99570 84306 99666
rect 84422 99570 87890 99666
rect 88006 99570 89418 99666
rect 854 430 89418 99570
rect 854 350 4562 430
rect 4678 350 5458 430
rect 5574 350 6354 430
rect 6470 350 7250 430
rect 7366 350 8146 430
rect 8262 350 9042 430
rect 9158 350 9938 430
rect 10054 350 10834 430
rect 10950 350 11730 430
rect 11846 350 12626 430
rect 12742 350 13522 430
rect 13638 350 14418 430
rect 14534 350 15314 430
rect 15430 350 16210 430
rect 16326 350 17106 430
rect 17222 350 18002 430
rect 18118 350 18898 430
rect 19014 350 19794 430
rect 19910 350 20690 430
rect 20806 350 21586 430
rect 21702 350 22482 430
rect 22598 350 23378 430
rect 23494 350 24274 430
rect 24390 350 25170 430
rect 25286 350 26066 430
rect 26182 350 26962 430
rect 27078 350 27858 430
rect 27974 350 28754 430
rect 28870 350 29650 430
rect 29766 350 30546 430
rect 30662 350 31442 430
rect 31558 350 32338 430
rect 32454 350 33234 430
rect 33350 350 34130 430
rect 34246 350 35026 430
rect 35142 350 35922 430
rect 36038 350 36818 430
rect 36934 350 37714 430
rect 37830 350 38610 430
rect 38726 350 39506 430
rect 39622 350 40402 430
rect 40518 350 41298 430
rect 41414 350 42194 430
rect 42310 350 43090 430
rect 43206 350 43986 430
rect 44102 350 44882 430
rect 44998 350 45778 430
rect 45894 350 46674 430
rect 46790 350 47570 430
rect 47686 350 48466 430
rect 48582 350 49362 430
rect 49478 350 50258 430
rect 50374 350 51154 430
rect 51270 350 52050 430
rect 52166 350 52946 430
rect 53062 350 53842 430
rect 53958 350 54738 430
rect 54854 350 55634 430
rect 55750 350 56530 430
rect 56646 350 57426 430
rect 57542 350 58322 430
rect 58438 350 59218 430
rect 59334 350 60114 430
rect 60230 350 61010 430
rect 61126 350 61906 430
rect 62022 350 62802 430
rect 62918 350 63698 430
rect 63814 350 64594 430
rect 64710 350 65490 430
rect 65606 350 66386 430
rect 66502 350 67282 430
rect 67398 350 68178 430
rect 68294 350 69074 430
rect 69190 350 69970 430
rect 70086 350 70866 430
rect 70982 350 71762 430
rect 71878 350 72658 430
rect 72774 350 73554 430
rect 73670 350 74450 430
rect 74566 350 75346 430
rect 75462 350 76242 430
rect 76358 350 77138 430
rect 77254 350 78034 430
rect 78150 350 78930 430
rect 79046 350 79826 430
rect 79942 350 80722 430
rect 80838 350 81618 430
rect 81734 350 82514 430
rect 82630 350 83410 430
rect 83526 350 84306 430
rect 84422 350 85202 430
rect 85318 350 89418 430
<< metal3 >>
rect 0 97552 400 97608
rect 0 95648 400 95704
rect 89600 95312 90000 95368
rect 89600 94304 90000 94360
rect 0 93744 400 93800
rect 89600 93296 90000 93352
rect 89600 92288 90000 92344
rect 0 91840 400 91896
rect 89600 91280 90000 91336
rect 89600 90272 90000 90328
rect 0 89936 400 89992
rect 89600 89264 90000 89320
rect 89600 88256 90000 88312
rect 0 88032 400 88088
rect 89600 87248 90000 87304
rect 89600 86240 90000 86296
rect 0 86128 400 86184
rect 89600 85232 90000 85288
rect 0 84224 400 84280
rect 89600 84224 90000 84280
rect 89600 83216 90000 83272
rect 0 82320 400 82376
rect 89600 82208 90000 82264
rect 89600 81200 90000 81256
rect 0 80416 400 80472
rect 89600 80192 90000 80248
rect 89600 79184 90000 79240
rect 0 78512 400 78568
rect 89600 78176 90000 78232
rect 89600 77168 90000 77224
rect 0 76608 400 76664
rect 89600 76160 90000 76216
rect 89600 75152 90000 75208
rect 0 74704 400 74760
rect 89600 74144 90000 74200
rect 89600 73136 90000 73192
rect 0 72800 400 72856
rect 89600 72128 90000 72184
rect 89600 71120 90000 71176
rect 0 70896 400 70952
rect 89600 70112 90000 70168
rect 89600 69104 90000 69160
rect 0 68992 400 69048
rect 89600 68096 90000 68152
rect 0 67088 400 67144
rect 89600 67088 90000 67144
rect 89600 66080 90000 66136
rect 0 65184 400 65240
rect 89600 65072 90000 65128
rect 89600 64064 90000 64120
rect 0 63280 400 63336
rect 89600 63056 90000 63112
rect 89600 62048 90000 62104
rect 0 61376 400 61432
rect 89600 61040 90000 61096
rect 89600 60032 90000 60088
rect 0 59472 400 59528
rect 89600 59024 90000 59080
rect 89600 58016 90000 58072
rect 0 57568 400 57624
rect 89600 57008 90000 57064
rect 89600 56000 90000 56056
rect 0 55664 400 55720
rect 89600 54992 90000 55048
rect 89600 53984 90000 54040
rect 0 53760 400 53816
rect 89600 52976 90000 53032
rect 89600 51968 90000 52024
rect 0 51856 400 51912
rect 89600 50960 90000 51016
rect 0 49952 400 50008
rect 89600 49952 90000 50008
rect 89600 48944 90000 49000
rect 0 48048 400 48104
rect 89600 47936 90000 47992
rect 89600 46928 90000 46984
rect 0 46144 400 46200
rect 89600 45920 90000 45976
rect 89600 44912 90000 44968
rect 0 44240 400 44296
rect 89600 43904 90000 43960
rect 89600 42896 90000 42952
rect 0 42336 400 42392
rect 89600 41888 90000 41944
rect 89600 40880 90000 40936
rect 0 40432 400 40488
rect 89600 39872 90000 39928
rect 89600 38864 90000 38920
rect 0 38528 400 38584
rect 89600 37856 90000 37912
rect 89600 36848 90000 36904
rect 0 36624 400 36680
rect 89600 35840 90000 35896
rect 89600 34832 90000 34888
rect 0 34720 400 34776
rect 89600 33824 90000 33880
rect 0 32816 400 32872
rect 89600 32816 90000 32872
rect 89600 31808 90000 31864
rect 0 30912 400 30968
rect 89600 30800 90000 30856
rect 89600 29792 90000 29848
rect 0 29008 400 29064
rect 89600 28784 90000 28840
rect 89600 27776 90000 27832
rect 0 27104 400 27160
rect 89600 26768 90000 26824
rect 89600 25760 90000 25816
rect 0 25200 400 25256
rect 89600 24752 90000 24808
rect 89600 23744 90000 23800
rect 0 23296 400 23352
rect 89600 22736 90000 22792
rect 89600 21728 90000 21784
rect 0 21392 400 21448
rect 89600 20720 90000 20776
rect 89600 19712 90000 19768
rect 0 19488 400 19544
rect 89600 18704 90000 18760
rect 89600 17696 90000 17752
rect 0 17584 400 17640
rect 89600 16688 90000 16744
rect 0 15680 400 15736
rect 89600 15680 90000 15736
rect 89600 14672 90000 14728
rect 0 13776 400 13832
rect 89600 13664 90000 13720
rect 89600 12656 90000 12712
rect 0 11872 400 11928
rect 89600 11648 90000 11704
rect 89600 10640 90000 10696
rect 0 9968 400 10024
rect 89600 9632 90000 9688
rect 89600 8624 90000 8680
rect 0 8064 400 8120
rect 89600 7616 90000 7672
rect 89600 6608 90000 6664
rect 0 6160 400 6216
rect 89600 5600 90000 5656
rect 89600 4592 90000 4648
rect 0 4256 400 4312
rect 0 2352 400 2408
<< obsm3 >>
rect 400 97638 89600 98406
rect 430 97522 89600 97638
rect 400 95734 89600 97522
rect 430 95618 89600 95734
rect 400 95398 89600 95618
rect 400 95282 89570 95398
rect 400 94390 89600 95282
rect 400 94274 89570 94390
rect 400 93830 89600 94274
rect 430 93714 89600 93830
rect 400 93382 89600 93714
rect 400 93266 89570 93382
rect 400 92374 89600 93266
rect 400 92258 89570 92374
rect 400 91926 89600 92258
rect 430 91810 89600 91926
rect 400 91366 89600 91810
rect 400 91250 89570 91366
rect 400 90358 89600 91250
rect 400 90242 89570 90358
rect 400 90022 89600 90242
rect 430 89906 89600 90022
rect 400 89350 89600 89906
rect 400 89234 89570 89350
rect 400 88342 89600 89234
rect 400 88226 89570 88342
rect 400 88118 89600 88226
rect 430 88002 89600 88118
rect 400 87334 89600 88002
rect 400 87218 89570 87334
rect 400 86326 89600 87218
rect 400 86214 89570 86326
rect 430 86210 89570 86214
rect 430 86098 89600 86210
rect 400 85318 89600 86098
rect 400 85202 89570 85318
rect 400 84310 89600 85202
rect 430 84194 89570 84310
rect 400 83302 89600 84194
rect 400 83186 89570 83302
rect 400 82406 89600 83186
rect 430 82294 89600 82406
rect 430 82290 89570 82294
rect 400 82178 89570 82290
rect 400 81286 89600 82178
rect 400 81170 89570 81286
rect 400 80502 89600 81170
rect 430 80386 89600 80502
rect 400 80278 89600 80386
rect 400 80162 89570 80278
rect 400 79270 89600 80162
rect 400 79154 89570 79270
rect 400 78598 89600 79154
rect 430 78482 89600 78598
rect 400 78262 89600 78482
rect 400 78146 89570 78262
rect 400 77254 89600 78146
rect 400 77138 89570 77254
rect 400 76694 89600 77138
rect 430 76578 89600 76694
rect 400 76246 89600 76578
rect 400 76130 89570 76246
rect 400 75238 89600 76130
rect 400 75122 89570 75238
rect 400 74790 89600 75122
rect 430 74674 89600 74790
rect 400 74230 89600 74674
rect 400 74114 89570 74230
rect 400 73222 89600 74114
rect 400 73106 89570 73222
rect 400 72886 89600 73106
rect 430 72770 89600 72886
rect 400 72214 89600 72770
rect 400 72098 89570 72214
rect 400 71206 89600 72098
rect 400 71090 89570 71206
rect 400 70982 89600 71090
rect 430 70866 89600 70982
rect 400 70198 89600 70866
rect 400 70082 89570 70198
rect 400 69190 89600 70082
rect 400 69078 89570 69190
rect 430 69074 89570 69078
rect 430 68962 89600 69074
rect 400 68182 89600 68962
rect 400 68066 89570 68182
rect 400 67174 89600 68066
rect 430 67058 89570 67174
rect 400 66166 89600 67058
rect 400 66050 89570 66166
rect 400 65270 89600 66050
rect 430 65158 89600 65270
rect 430 65154 89570 65158
rect 400 65042 89570 65154
rect 400 64150 89600 65042
rect 400 64034 89570 64150
rect 400 63366 89600 64034
rect 430 63250 89600 63366
rect 400 63142 89600 63250
rect 400 63026 89570 63142
rect 400 62134 89600 63026
rect 400 62018 89570 62134
rect 400 61462 89600 62018
rect 430 61346 89600 61462
rect 400 61126 89600 61346
rect 400 61010 89570 61126
rect 400 60118 89600 61010
rect 400 60002 89570 60118
rect 400 59558 89600 60002
rect 430 59442 89600 59558
rect 400 59110 89600 59442
rect 400 58994 89570 59110
rect 400 58102 89600 58994
rect 400 57986 89570 58102
rect 400 57654 89600 57986
rect 430 57538 89600 57654
rect 400 57094 89600 57538
rect 400 56978 89570 57094
rect 400 56086 89600 56978
rect 400 55970 89570 56086
rect 400 55750 89600 55970
rect 430 55634 89600 55750
rect 400 55078 89600 55634
rect 400 54962 89570 55078
rect 400 54070 89600 54962
rect 400 53954 89570 54070
rect 400 53846 89600 53954
rect 430 53730 89600 53846
rect 400 53062 89600 53730
rect 400 52946 89570 53062
rect 400 52054 89600 52946
rect 400 51942 89570 52054
rect 430 51938 89570 51942
rect 430 51826 89600 51938
rect 400 51046 89600 51826
rect 400 50930 89570 51046
rect 400 50038 89600 50930
rect 430 49922 89570 50038
rect 400 49030 89600 49922
rect 400 48914 89570 49030
rect 400 48134 89600 48914
rect 430 48022 89600 48134
rect 430 48018 89570 48022
rect 400 47906 89570 48018
rect 400 47014 89600 47906
rect 400 46898 89570 47014
rect 400 46230 89600 46898
rect 430 46114 89600 46230
rect 400 46006 89600 46114
rect 400 45890 89570 46006
rect 400 44998 89600 45890
rect 400 44882 89570 44998
rect 400 44326 89600 44882
rect 430 44210 89600 44326
rect 400 43990 89600 44210
rect 400 43874 89570 43990
rect 400 42982 89600 43874
rect 400 42866 89570 42982
rect 400 42422 89600 42866
rect 430 42306 89600 42422
rect 400 41974 89600 42306
rect 400 41858 89570 41974
rect 400 40966 89600 41858
rect 400 40850 89570 40966
rect 400 40518 89600 40850
rect 430 40402 89600 40518
rect 400 39958 89600 40402
rect 400 39842 89570 39958
rect 400 38950 89600 39842
rect 400 38834 89570 38950
rect 400 38614 89600 38834
rect 430 38498 89600 38614
rect 400 37942 89600 38498
rect 400 37826 89570 37942
rect 400 36934 89600 37826
rect 400 36818 89570 36934
rect 400 36710 89600 36818
rect 430 36594 89600 36710
rect 400 35926 89600 36594
rect 400 35810 89570 35926
rect 400 34918 89600 35810
rect 400 34806 89570 34918
rect 430 34802 89570 34806
rect 430 34690 89600 34802
rect 400 33910 89600 34690
rect 400 33794 89570 33910
rect 400 32902 89600 33794
rect 430 32786 89570 32902
rect 400 31894 89600 32786
rect 400 31778 89570 31894
rect 400 30998 89600 31778
rect 430 30886 89600 30998
rect 430 30882 89570 30886
rect 400 30770 89570 30882
rect 400 29878 89600 30770
rect 400 29762 89570 29878
rect 400 29094 89600 29762
rect 430 28978 89600 29094
rect 400 28870 89600 28978
rect 400 28754 89570 28870
rect 400 27862 89600 28754
rect 400 27746 89570 27862
rect 400 27190 89600 27746
rect 430 27074 89600 27190
rect 400 26854 89600 27074
rect 400 26738 89570 26854
rect 400 25846 89600 26738
rect 400 25730 89570 25846
rect 400 25286 89600 25730
rect 430 25170 89600 25286
rect 400 24838 89600 25170
rect 400 24722 89570 24838
rect 400 23830 89600 24722
rect 400 23714 89570 23830
rect 400 23382 89600 23714
rect 430 23266 89600 23382
rect 400 22822 89600 23266
rect 400 22706 89570 22822
rect 400 21814 89600 22706
rect 400 21698 89570 21814
rect 400 21478 89600 21698
rect 430 21362 89600 21478
rect 400 20806 89600 21362
rect 400 20690 89570 20806
rect 400 19798 89600 20690
rect 400 19682 89570 19798
rect 400 19574 89600 19682
rect 430 19458 89600 19574
rect 400 18790 89600 19458
rect 400 18674 89570 18790
rect 400 17782 89600 18674
rect 400 17670 89570 17782
rect 430 17666 89570 17670
rect 430 17554 89600 17666
rect 400 16774 89600 17554
rect 400 16658 89570 16774
rect 400 15766 89600 16658
rect 430 15650 89570 15766
rect 400 14758 89600 15650
rect 400 14642 89570 14758
rect 400 13862 89600 14642
rect 430 13750 89600 13862
rect 430 13746 89570 13750
rect 400 13634 89570 13746
rect 400 12742 89600 13634
rect 400 12626 89570 12742
rect 400 11958 89600 12626
rect 430 11842 89600 11958
rect 400 11734 89600 11842
rect 400 11618 89570 11734
rect 400 10726 89600 11618
rect 400 10610 89570 10726
rect 400 10054 89600 10610
rect 430 9938 89600 10054
rect 400 9718 89600 9938
rect 400 9602 89570 9718
rect 400 8710 89600 9602
rect 400 8594 89570 8710
rect 400 8150 89600 8594
rect 430 8034 89600 8150
rect 400 7702 89600 8034
rect 400 7586 89570 7702
rect 400 6694 89600 7586
rect 400 6578 89570 6694
rect 400 6246 89600 6578
rect 430 6130 89600 6246
rect 400 5686 89600 6130
rect 400 5570 89570 5686
rect 400 4678 89600 5570
rect 400 4562 89570 4678
rect 400 4342 89600 4562
rect 430 4226 89600 4342
rect 400 2438 89600 4226
rect 430 2322 89600 2438
rect 400 1554 89600 2322
<< metal4 >>
rect 2224 1538 2384 98422
rect 9904 1538 10064 98422
rect 17584 1538 17744 98422
rect 25264 1538 25424 98422
rect 32944 1538 33104 98422
rect 40624 1538 40784 98422
rect 48304 1538 48464 98422
rect 55984 1538 56144 98422
rect 63664 1538 63824 98422
rect 71344 1538 71504 98422
rect 79024 1538 79184 98422
rect 86704 1538 86864 98422
<< obsm4 >>
rect 1526 1731 2194 93511
rect 2414 1731 9874 93511
rect 10094 1731 17554 93511
rect 17774 1731 25234 93511
rect 25454 1731 32914 93511
rect 33134 1731 40594 93511
rect 40814 1731 48274 93511
rect 48494 1731 55954 93511
rect 56174 1731 63634 93511
rect 63854 1731 71314 93511
rect 71534 1731 78994 93511
rect 79214 1731 86674 93511
rect 86894 1731 89138 93511
<< obsm5 >>
rect 4374 1733 88642 79087
<< labels >>
rlabel metal3 s 0 93744 400 93800 6 digital_io_in[21]
port 1 nsew signal input
rlabel metal3 s 0 88032 400 88088 6 digital_io_in[22]
port 2 nsew signal input
rlabel metal3 s 0 82320 400 82376 6 digital_io_in[23]
port 3 nsew signal input
rlabel metal3 s 0 80416 400 80472 6 digital_io_in[24]
port 4 nsew signal input
rlabel metal3 s 0 74704 400 74760 6 digital_io_in[25]
port 5 nsew signal input
rlabel metal3 s 0 68992 400 69048 6 digital_io_in[26]
port 6 nsew signal input
rlabel metal3 s 0 63280 400 63336 6 digital_io_in[27]
port 7 nsew signal input
rlabel metal3 s 0 57568 400 57624 6 digital_io_in[28]
port 8 nsew signal input
rlabel metal3 s 0 51856 400 51912 6 digital_io_in[29]
port 9 nsew signal input
rlabel metal3 s 0 46144 400 46200 6 digital_io_in[30]
port 10 nsew signal input
rlabel metal3 s 0 40432 400 40488 6 digital_io_in[31]
port 11 nsew signal input
rlabel metal3 s 0 34720 400 34776 6 digital_io_in[32]
port 12 nsew signal input
rlabel metal3 s 0 29008 400 29064 6 digital_io_in[33]
port 13 nsew signal input
rlabel metal3 s 0 23296 400 23352 6 digital_io_in[34]
port 14 nsew signal input
rlabel metal3 s 0 17584 400 17640 6 digital_io_in[35]
port 15 nsew signal input
rlabel metal3 s 0 11872 400 11928 6 digital_io_in[36]
port 16 nsew signal input
rlabel metal3 s 0 6160 400 6216 6 digital_io_in[37]
port 17 nsew signal input
rlabel metal3 s 0 97552 400 97608 6 digital_io_oen[21]
port 18 nsew signal output
rlabel metal3 s 0 91840 400 91896 6 digital_io_oen[22]
port 19 nsew signal output
rlabel metal3 s 0 86128 400 86184 6 digital_io_oen[23]
port 20 nsew signal output
rlabel metal3 s 0 76608 400 76664 6 digital_io_oen[24]
port 21 nsew signal output
rlabel metal3 s 0 70896 400 70952 6 digital_io_oen[25]
port 22 nsew signal output
rlabel metal3 s 0 65184 400 65240 6 digital_io_oen[26]
port 23 nsew signal output
rlabel metal3 s 0 59472 400 59528 6 digital_io_oen[27]
port 24 nsew signal output
rlabel metal3 s 0 53760 400 53816 6 digital_io_oen[28]
port 25 nsew signal output
rlabel metal3 s 0 48048 400 48104 6 digital_io_oen[29]
port 26 nsew signal output
rlabel metal3 s 0 42336 400 42392 6 digital_io_oen[30]
port 27 nsew signal output
rlabel metal3 s 0 36624 400 36680 6 digital_io_oen[31]
port 28 nsew signal output
rlabel metal3 s 0 30912 400 30968 6 digital_io_oen[32]
port 29 nsew signal output
rlabel metal3 s 0 25200 400 25256 6 digital_io_oen[33]
port 30 nsew signal output
rlabel metal3 s 0 19488 400 19544 6 digital_io_oen[34]
port 31 nsew signal output
rlabel metal3 s 0 13776 400 13832 6 digital_io_oen[35]
port 32 nsew signal output
rlabel metal3 s 0 8064 400 8120 6 digital_io_oen[36]
port 33 nsew signal output
rlabel metal3 s 0 2352 400 2408 6 digital_io_oen[37]
port 34 nsew signal output
rlabel metal3 s 0 95648 400 95704 6 digital_io_out[21]
port 35 nsew signal output
rlabel metal3 s 0 89936 400 89992 6 digital_io_out[22]
port 36 nsew signal output
rlabel metal3 s 0 84224 400 84280 6 digital_io_out[23]
port 37 nsew signal output
rlabel metal3 s 0 78512 400 78568 6 digital_io_out[24]
port 38 nsew signal output
rlabel metal3 s 0 72800 400 72856 6 digital_io_out[25]
port 39 nsew signal output
rlabel metal3 s 0 67088 400 67144 6 digital_io_out[26]
port 40 nsew signal output
rlabel metal3 s 0 61376 400 61432 6 digital_io_out[27]
port 41 nsew signal output
rlabel metal3 s 0 55664 400 55720 6 digital_io_out[28]
port 42 nsew signal output
rlabel metal3 s 0 49952 400 50008 6 digital_io_out[29]
port 43 nsew signal output
rlabel metal3 s 0 44240 400 44296 6 digital_io_out[30]
port 44 nsew signal output
rlabel metal3 s 0 38528 400 38584 6 digital_io_out[31]
port 45 nsew signal output
rlabel metal3 s 0 32816 400 32872 6 digital_io_out[32]
port 46 nsew signal output
rlabel metal3 s 0 27104 400 27160 6 digital_io_out[33]
port 47 nsew signal output
rlabel metal3 s 0 21392 400 21448 6 digital_io_out[34]
port 48 nsew signal output
rlabel metal3 s 0 15680 400 15736 6 digital_io_out[35]
port 49 nsew signal output
rlabel metal3 s 0 9968 400 10024 6 digital_io_out[36]
port 50 nsew signal output
rlabel metal3 s 0 4256 400 4312 6 digital_io_out[37]
port 51 nsew signal output
rlabel metal2 s 8176 0 8232 400 6 e_reset_n
port 52 nsew signal input
rlabel metal2 s 48496 99600 48552 100000 6 i2cm_clk_i
port 53 nsew signal output
rlabel metal2 s 44912 99600 44968 100000 6 i2cm_clk_o
port 54 nsew signal input
rlabel metal2 s 52080 99600 52136 100000 6 i2cm_clk_oen
port 55 nsew signal input
rlabel metal2 s 62832 99600 62888 100000 6 i2cm_data_i
port 56 nsew signal output
rlabel metal2 s 59248 99600 59304 100000 6 i2cm_data_o
port 57 nsew signal input
rlabel metal2 s 55664 99600 55720 100000 6 i2cm_data_oen
port 58 nsew signal input
rlabel metal2 s 34160 99600 34216 100000 6 i2cm_intr
port 59 nsew signal input
rlabel metal2 s 12656 99600 12712 100000 6 i2cm_rst_n
port 60 nsew signal output
rlabel metal2 s 4592 0 4648 400 6 mclk
port 61 nsew signal input
rlabel metal2 s 7280 0 7336 400 6 p_reset_n
port 62 nsew signal input
rlabel metal2 s 41328 99600 41384 100000 6 pulse1m_mclk
port 63 nsew signal output
rlabel metal2 s 82544 0 82600 400 6 reg_ack
port 64 nsew signal output
rlabel metal2 s 20720 0 20776 400 6 reg_addr[0]
port 65 nsew signal input
rlabel metal2 s 11760 0 11816 400 6 reg_addr[10]
port 66 nsew signal input
rlabel metal2 s 19824 0 19880 400 6 reg_addr[1]
port 67 nsew signal input
rlabel metal2 s 18928 0 18984 400 6 reg_addr[2]
port 68 nsew signal input
rlabel metal2 s 18032 0 18088 400 6 reg_addr[3]
port 69 nsew signal input
rlabel metal2 s 17136 0 17192 400 6 reg_addr[4]
port 70 nsew signal input
rlabel metal2 s 16240 0 16296 400 6 reg_addr[5]
port 71 nsew signal input
rlabel metal2 s 15344 0 15400 400 6 reg_addr[6]
port 72 nsew signal input
rlabel metal2 s 14448 0 14504 400 6 reg_addr[7]
port 73 nsew signal input
rlabel metal2 s 13552 0 13608 400 6 reg_addr[8]
port 74 nsew signal input
rlabel metal2 s 12656 0 12712 400 6 reg_addr[9]
port 75 nsew signal input
rlabel metal2 s 24304 0 24360 400 6 reg_be[0]
port 76 nsew signal input
rlabel metal2 s 23408 0 23464 400 6 reg_be[1]
port 77 nsew signal input
rlabel metal2 s 22512 0 22568 400 6 reg_be[2]
port 78 nsew signal input
rlabel metal2 s 21616 0 21672 400 6 reg_be[3]
port 79 nsew signal input
rlabel metal2 s 9968 0 10024 400 6 reg_cs
port 80 nsew signal input
rlabel metal3 s 89600 95312 90000 95368 6 reg_peri_ack
port 81 nsew signal input
rlabel metal3 s 89600 25760 90000 25816 6 reg_peri_addr[0]
port 82 nsew signal output
rlabel metal3 s 89600 15680 90000 15736 6 reg_peri_addr[10]
port 83 nsew signal output
rlabel metal3 s 89600 24752 90000 24808 6 reg_peri_addr[1]
port 84 nsew signal output
rlabel metal3 s 89600 23744 90000 23800 6 reg_peri_addr[2]
port 85 nsew signal output
rlabel metal3 s 89600 22736 90000 22792 6 reg_peri_addr[3]
port 86 nsew signal output
rlabel metal3 s 89600 21728 90000 21784 6 reg_peri_addr[4]
port 87 nsew signal output
rlabel metal3 s 89600 20720 90000 20776 6 reg_peri_addr[5]
port 88 nsew signal output
rlabel metal3 s 89600 19712 90000 19768 6 reg_peri_addr[6]
port 89 nsew signal output
rlabel metal3 s 89600 18704 90000 18760 6 reg_peri_addr[7]
port 90 nsew signal output
rlabel metal3 s 89600 17696 90000 17752 6 reg_peri_addr[8]
port 91 nsew signal output
rlabel metal3 s 89600 16688 90000 16744 6 reg_peri_addr[9]
port 92 nsew signal output
rlabel metal3 s 89600 29792 90000 29848 6 reg_peri_be[0]
port 93 nsew signal output
rlabel metal3 s 89600 28784 90000 28840 6 reg_peri_be[1]
port 94 nsew signal output
rlabel metal3 s 89600 27776 90000 27832 6 reg_peri_be[2]
port 95 nsew signal output
rlabel metal3 s 89600 26768 90000 26824 6 reg_peri_be[3]
port 96 nsew signal output
rlabel metal3 s 89600 13664 90000 13720 6 reg_peri_cs
port 97 nsew signal output
rlabel metal3 s 89600 94304 90000 94360 6 reg_peri_rdata[0]
port 98 nsew signal input
rlabel metal3 s 89600 84224 90000 84280 6 reg_peri_rdata[10]
port 99 nsew signal input
rlabel metal3 s 89600 83216 90000 83272 6 reg_peri_rdata[11]
port 100 nsew signal input
rlabel metal3 s 89600 82208 90000 82264 6 reg_peri_rdata[12]
port 101 nsew signal input
rlabel metal3 s 89600 81200 90000 81256 6 reg_peri_rdata[13]
port 102 nsew signal input
rlabel metal3 s 89600 80192 90000 80248 6 reg_peri_rdata[14]
port 103 nsew signal input
rlabel metal3 s 89600 79184 90000 79240 6 reg_peri_rdata[15]
port 104 nsew signal input
rlabel metal3 s 89600 78176 90000 78232 6 reg_peri_rdata[16]
port 105 nsew signal input
rlabel metal3 s 89600 77168 90000 77224 6 reg_peri_rdata[17]
port 106 nsew signal input
rlabel metal3 s 89600 76160 90000 76216 6 reg_peri_rdata[18]
port 107 nsew signal input
rlabel metal3 s 89600 75152 90000 75208 6 reg_peri_rdata[19]
port 108 nsew signal input
rlabel metal3 s 89600 93296 90000 93352 6 reg_peri_rdata[1]
port 109 nsew signal input
rlabel metal3 s 89600 74144 90000 74200 6 reg_peri_rdata[20]
port 110 nsew signal input
rlabel metal3 s 89600 73136 90000 73192 6 reg_peri_rdata[21]
port 111 nsew signal input
rlabel metal3 s 89600 72128 90000 72184 6 reg_peri_rdata[22]
port 112 nsew signal input
rlabel metal3 s 89600 71120 90000 71176 6 reg_peri_rdata[23]
port 113 nsew signal input
rlabel metal3 s 89600 70112 90000 70168 6 reg_peri_rdata[24]
port 114 nsew signal input
rlabel metal3 s 89600 69104 90000 69160 6 reg_peri_rdata[25]
port 115 nsew signal input
rlabel metal3 s 89600 68096 90000 68152 6 reg_peri_rdata[26]
port 116 nsew signal input
rlabel metal3 s 89600 67088 90000 67144 6 reg_peri_rdata[27]
port 117 nsew signal input
rlabel metal3 s 89600 66080 90000 66136 6 reg_peri_rdata[28]
port 118 nsew signal input
rlabel metal3 s 89600 65072 90000 65128 6 reg_peri_rdata[29]
port 119 nsew signal input
rlabel metal3 s 89600 92288 90000 92344 6 reg_peri_rdata[2]
port 120 nsew signal input
rlabel metal3 s 89600 64064 90000 64120 6 reg_peri_rdata[30]
port 121 nsew signal input
rlabel metal3 s 89600 63056 90000 63112 6 reg_peri_rdata[31]
port 122 nsew signal input
rlabel metal3 s 89600 91280 90000 91336 6 reg_peri_rdata[3]
port 123 nsew signal input
rlabel metal3 s 89600 90272 90000 90328 6 reg_peri_rdata[4]
port 124 nsew signal input
rlabel metal3 s 89600 89264 90000 89320 6 reg_peri_rdata[5]
port 125 nsew signal input
rlabel metal3 s 89600 88256 90000 88312 6 reg_peri_rdata[6]
port 126 nsew signal input
rlabel metal3 s 89600 87248 90000 87304 6 reg_peri_rdata[7]
port 127 nsew signal input
rlabel metal3 s 89600 86240 90000 86296 6 reg_peri_rdata[8]
port 128 nsew signal input
rlabel metal3 s 89600 85232 90000 85288 6 reg_peri_rdata[9]
port 129 nsew signal input
rlabel metal3 s 89600 62048 90000 62104 6 reg_peri_wdata[0]
port 130 nsew signal output
rlabel metal3 s 89600 51968 90000 52024 6 reg_peri_wdata[10]
port 131 nsew signal output
rlabel metal3 s 89600 50960 90000 51016 6 reg_peri_wdata[11]
port 132 nsew signal output
rlabel metal3 s 89600 49952 90000 50008 6 reg_peri_wdata[12]
port 133 nsew signal output
rlabel metal3 s 89600 48944 90000 49000 6 reg_peri_wdata[13]
port 134 nsew signal output
rlabel metal3 s 89600 47936 90000 47992 6 reg_peri_wdata[14]
port 135 nsew signal output
rlabel metal3 s 89600 46928 90000 46984 6 reg_peri_wdata[15]
port 136 nsew signal output
rlabel metal3 s 89600 45920 90000 45976 6 reg_peri_wdata[16]
port 137 nsew signal output
rlabel metal3 s 89600 44912 90000 44968 6 reg_peri_wdata[17]
port 138 nsew signal output
rlabel metal3 s 89600 43904 90000 43960 6 reg_peri_wdata[18]
port 139 nsew signal output
rlabel metal3 s 89600 42896 90000 42952 6 reg_peri_wdata[19]
port 140 nsew signal output
rlabel metal3 s 89600 61040 90000 61096 6 reg_peri_wdata[1]
port 141 nsew signal output
rlabel metal3 s 89600 41888 90000 41944 6 reg_peri_wdata[20]
port 142 nsew signal output
rlabel metal3 s 89600 40880 90000 40936 6 reg_peri_wdata[21]
port 143 nsew signal output
rlabel metal3 s 89600 39872 90000 39928 6 reg_peri_wdata[22]
port 144 nsew signal output
rlabel metal3 s 89600 38864 90000 38920 6 reg_peri_wdata[23]
port 145 nsew signal output
rlabel metal3 s 89600 37856 90000 37912 6 reg_peri_wdata[24]
port 146 nsew signal output
rlabel metal3 s 89600 36848 90000 36904 6 reg_peri_wdata[25]
port 147 nsew signal output
rlabel metal3 s 89600 35840 90000 35896 6 reg_peri_wdata[26]
port 148 nsew signal output
rlabel metal3 s 89600 34832 90000 34888 6 reg_peri_wdata[27]
port 149 nsew signal output
rlabel metal3 s 89600 33824 90000 33880 6 reg_peri_wdata[28]
port 150 nsew signal output
rlabel metal3 s 89600 32816 90000 32872 6 reg_peri_wdata[29]
port 151 nsew signal output
rlabel metal3 s 89600 60032 90000 60088 6 reg_peri_wdata[2]
port 152 nsew signal output
rlabel metal3 s 89600 31808 90000 31864 6 reg_peri_wdata[30]
port 153 nsew signal output
rlabel metal3 s 89600 30800 90000 30856 6 reg_peri_wdata[31]
port 154 nsew signal output
rlabel metal3 s 89600 59024 90000 59080 6 reg_peri_wdata[3]
port 155 nsew signal output
rlabel metal3 s 89600 58016 90000 58072 6 reg_peri_wdata[4]
port 156 nsew signal output
rlabel metal3 s 89600 57008 90000 57064 6 reg_peri_wdata[5]
port 157 nsew signal output
rlabel metal3 s 89600 56000 90000 56056 6 reg_peri_wdata[6]
port 158 nsew signal output
rlabel metal3 s 89600 54992 90000 55048 6 reg_peri_wdata[7]
port 159 nsew signal output
rlabel metal3 s 89600 53984 90000 54040 6 reg_peri_wdata[8]
port 160 nsew signal output
rlabel metal3 s 89600 52976 90000 53032 6 reg_peri_wdata[9]
port 161 nsew signal output
rlabel metal3 s 89600 14672 90000 14728 6 reg_peri_wr
port 162 nsew signal output
rlabel metal2 s 81648 0 81704 400 6 reg_rdata[0]
port 163 nsew signal output
rlabel metal2 s 72688 0 72744 400 6 reg_rdata[10]
port 164 nsew signal output
rlabel metal2 s 71792 0 71848 400 6 reg_rdata[11]
port 165 nsew signal output
rlabel metal2 s 70896 0 70952 400 6 reg_rdata[12]
port 166 nsew signal output
rlabel metal2 s 70000 0 70056 400 6 reg_rdata[13]
port 167 nsew signal output
rlabel metal2 s 69104 0 69160 400 6 reg_rdata[14]
port 168 nsew signal output
rlabel metal2 s 68208 0 68264 400 6 reg_rdata[15]
port 169 nsew signal output
rlabel metal2 s 67312 0 67368 400 6 reg_rdata[16]
port 170 nsew signal output
rlabel metal2 s 66416 0 66472 400 6 reg_rdata[17]
port 171 nsew signal output
rlabel metal2 s 65520 0 65576 400 6 reg_rdata[18]
port 172 nsew signal output
rlabel metal2 s 64624 0 64680 400 6 reg_rdata[19]
port 173 nsew signal output
rlabel metal2 s 80752 0 80808 400 6 reg_rdata[1]
port 174 nsew signal output
rlabel metal2 s 63728 0 63784 400 6 reg_rdata[20]
port 175 nsew signal output
rlabel metal2 s 62832 0 62888 400 6 reg_rdata[21]
port 176 nsew signal output
rlabel metal2 s 61936 0 61992 400 6 reg_rdata[22]
port 177 nsew signal output
rlabel metal2 s 61040 0 61096 400 6 reg_rdata[23]
port 178 nsew signal output
rlabel metal2 s 60144 0 60200 400 6 reg_rdata[24]
port 179 nsew signal output
rlabel metal2 s 59248 0 59304 400 6 reg_rdata[25]
port 180 nsew signal output
rlabel metal2 s 58352 0 58408 400 6 reg_rdata[26]
port 181 nsew signal output
rlabel metal2 s 57456 0 57512 400 6 reg_rdata[27]
port 182 nsew signal output
rlabel metal2 s 56560 0 56616 400 6 reg_rdata[28]
port 183 nsew signal output
rlabel metal2 s 55664 0 55720 400 6 reg_rdata[29]
port 184 nsew signal output
rlabel metal2 s 79856 0 79912 400 6 reg_rdata[2]
port 185 nsew signal output
rlabel metal2 s 54768 0 54824 400 6 reg_rdata[30]
port 186 nsew signal output
rlabel metal2 s 53872 0 53928 400 6 reg_rdata[31]
port 187 nsew signal output
rlabel metal2 s 78960 0 79016 400 6 reg_rdata[3]
port 188 nsew signal output
rlabel metal2 s 78064 0 78120 400 6 reg_rdata[4]
port 189 nsew signal output
rlabel metal2 s 77168 0 77224 400 6 reg_rdata[5]
port 190 nsew signal output
rlabel metal2 s 76272 0 76328 400 6 reg_rdata[6]
port 191 nsew signal output
rlabel metal2 s 75376 0 75432 400 6 reg_rdata[7]
port 192 nsew signal output
rlabel metal2 s 74480 0 74536 400 6 reg_rdata[8]
port 193 nsew signal output
rlabel metal2 s 73584 0 73640 400 6 reg_rdata[9]
port 194 nsew signal output
rlabel metal2 s 52976 0 53032 400 6 reg_wdata[0]
port 195 nsew signal input
rlabel metal2 s 44016 0 44072 400 6 reg_wdata[10]
port 196 nsew signal input
rlabel metal2 s 43120 0 43176 400 6 reg_wdata[11]
port 197 nsew signal input
rlabel metal2 s 42224 0 42280 400 6 reg_wdata[12]
port 198 nsew signal input
rlabel metal2 s 41328 0 41384 400 6 reg_wdata[13]
port 199 nsew signal input
rlabel metal2 s 40432 0 40488 400 6 reg_wdata[14]
port 200 nsew signal input
rlabel metal2 s 39536 0 39592 400 6 reg_wdata[15]
port 201 nsew signal input
rlabel metal2 s 38640 0 38696 400 6 reg_wdata[16]
port 202 nsew signal input
rlabel metal2 s 37744 0 37800 400 6 reg_wdata[17]
port 203 nsew signal input
rlabel metal2 s 36848 0 36904 400 6 reg_wdata[18]
port 204 nsew signal input
rlabel metal2 s 35952 0 36008 400 6 reg_wdata[19]
port 205 nsew signal input
rlabel metal2 s 52080 0 52136 400 6 reg_wdata[1]
port 206 nsew signal input
rlabel metal2 s 35056 0 35112 400 6 reg_wdata[20]
port 207 nsew signal input
rlabel metal2 s 34160 0 34216 400 6 reg_wdata[21]
port 208 nsew signal input
rlabel metal2 s 33264 0 33320 400 6 reg_wdata[22]
port 209 nsew signal input
rlabel metal2 s 32368 0 32424 400 6 reg_wdata[23]
port 210 nsew signal input
rlabel metal2 s 31472 0 31528 400 6 reg_wdata[24]
port 211 nsew signal input
rlabel metal2 s 30576 0 30632 400 6 reg_wdata[25]
port 212 nsew signal input
rlabel metal2 s 29680 0 29736 400 6 reg_wdata[26]
port 213 nsew signal input
rlabel metal2 s 28784 0 28840 400 6 reg_wdata[27]
port 214 nsew signal input
rlabel metal2 s 27888 0 27944 400 6 reg_wdata[28]
port 215 nsew signal input
rlabel metal2 s 26992 0 27048 400 6 reg_wdata[29]
port 216 nsew signal input
rlabel metal2 s 51184 0 51240 400 6 reg_wdata[2]
port 217 nsew signal input
rlabel metal2 s 26096 0 26152 400 6 reg_wdata[30]
port 218 nsew signal input
rlabel metal2 s 25200 0 25256 400 6 reg_wdata[31]
port 219 nsew signal input
rlabel metal2 s 50288 0 50344 400 6 reg_wdata[3]
port 220 nsew signal input
rlabel metal2 s 49392 0 49448 400 6 reg_wdata[4]
port 221 nsew signal input
rlabel metal2 s 48496 0 48552 400 6 reg_wdata[5]
port 222 nsew signal input
rlabel metal2 s 47600 0 47656 400 6 reg_wdata[6]
port 223 nsew signal input
rlabel metal2 s 46704 0 46760 400 6 reg_wdata[7]
port 224 nsew signal input
rlabel metal2 s 45808 0 45864 400 6 reg_wdata[8]
port 225 nsew signal input
rlabel metal2 s 44912 0 44968 400 6 reg_wdata[9]
port 226 nsew signal input
rlabel metal2 s 10864 0 10920 400 6 reg_wr
port 227 nsew signal input
rlabel metal2 s 26992 99600 27048 100000 6 rtc_clk
port 228 nsew signal output
rlabel metal2 s 30576 99600 30632 100000 6 rtc_intr
port 229 nsew signal input
rlabel metal2 s 9072 0 9128 400 6 s_reset_n
port 230 nsew signal input
rlabel metal2 s 84336 99600 84392 100000 6 spim_miso
port 231 nsew signal input
rlabel metal2 s 87920 99600 87976 100000 6 spim_mosi
port 232 nsew signal output
rlabel metal2 s 66416 99600 66472 100000 6 spim_sck
port 233 nsew signal input
rlabel metal2 s 80752 99600 80808 100000 6 spim_ssn[0]
port 234 nsew signal input
rlabel metal2 s 77168 99600 77224 100000 6 spim_ssn[1]
port 235 nsew signal input
rlabel metal2 s 73584 99600 73640 100000 6 spim_ssn[2]
port 236 nsew signal input
rlabel metal2 s 70000 99600 70056 100000 6 spim_ssn[3]
port 237 nsew signal input
rlabel metal2 s 1904 99600 1960 100000 6 sspim_rst_n
port 238 nsew signal output
rlabel metal2 s 9072 99600 9128 100000 6 uart_rst_n[0]
port 239 nsew signal output
rlabel metal2 s 5488 99600 5544 100000 6 uart_rst_n[1]
port 240 nsew signal output
rlabel metal3 s 89600 12656 90000 12712 6 uart_rxd[0]
port 241 nsew signal output
rlabel metal3 s 89600 10640 90000 10696 6 uart_rxd[1]
port 242 nsew signal output
rlabel metal3 s 89600 11648 90000 11704 6 uart_txd[0]
port 243 nsew signal input
rlabel metal3 s 89600 9632 90000 9688 6 uart_txd[1]
port 244 nsew signal input
rlabel metal2 s 23408 99600 23464 100000 6 usb_clk
port 245 nsew signal output
rlabel metal3 s 89600 8624 90000 8680 6 usb_dn_i
port 246 nsew signal output
rlabel metal3 s 89600 5600 90000 5656 6 usb_dn_o
port 247 nsew signal input
rlabel metal3 s 89600 7616 90000 7672 6 usb_dp_i
port 248 nsew signal output
rlabel metal3 s 89600 4592 90000 4648 6 usb_dp_o
port 249 nsew signal input
rlabel metal2 s 37744 99600 37800 100000 6 usb_intr
port 250 nsew signal input
rlabel metal3 s 89600 6608 90000 6664 6 usb_oen
port 251 nsew signal input
rlabel metal2 s 16240 99600 16296 100000 6 usb_rst_n
port 252 nsew signal output
rlabel metal2 s 5488 0 5544 400 6 user_clock1
port 253 nsew signal input
rlabel metal2 s 6384 0 6440 400 6 user_clock2
port 254 nsew signal input
rlabel metal2 s 83440 0 83496 400 6 user_irq[0]
port 255 nsew signal output
rlabel metal2 s 84336 0 84392 400 6 user_irq[1]
port 256 nsew signal output
rlabel metal2 s 85232 0 85288 400 6 user_irq[2]
port 257 nsew signal output
rlabel metal4 s 2224 1538 2384 98422 6 vdd
port 258 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 98422 6 vdd
port 258 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 98422 6 vdd
port 258 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 98422 6 vdd
port 258 nsew power bidirectional
rlabel metal4 s 63664 1538 63824 98422 6 vdd
port 258 nsew power bidirectional
rlabel metal4 s 79024 1538 79184 98422 6 vdd
port 258 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 98422 6 vss
port 259 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 98422 6 vss
port 259 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 98422 6 vss
port 259 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 98422 6 vss
port 259 nsew ground bidirectional
rlabel metal4 s 71344 1538 71504 98422 6 vss
port 259 nsew ground bidirectional
rlabel metal4 s 86704 1538 86864 98422 6 vss
port 259 nsew ground bidirectional
rlabel metal2 s 19824 99600 19880 100000 6 xtal_clk
port 260 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 90000 100000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 27211058
string GDS_FILE /home/farag/carvel_riscv_soc/gf180mcu_riscv_soc/openlane/pinmux_top/runs/23_11_23_03_33/results/signoff/pinmux_top.magic.gds
string GDS_START 604018
<< end >>

