* NGSPICE file created from serv_rf_top.ext - technology: gf180mcuD

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_4 A1 A2 B1 B2 C1 C2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_4 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_2 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_2 A1 A2 B1 B2 C1 C2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_4 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_4 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_8 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_4 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_12 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_12 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_2 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_2 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_4 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_3 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_4 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_4 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_1 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_1 A1 A2 B1 B2 C1 C2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_4 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_3 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_4 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_2 A1 A2 A3 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_4 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_4 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_2 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_2 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_4 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_1 A1 A2 A3 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_4 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_2 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_2 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_4 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_2 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_4 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_4 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_2 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_12 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_12 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_2 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_2 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyb_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyb_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_2 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_3 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_2 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_4 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tiel abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tiel ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_4 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_1 I0 I1 I2 I3 S0 S1 Z VDD VNW VPW VSS
.ends

.subckt serv_rf_top clk i_dbus_ack i_dbus_rdt[0] i_dbus_rdt[10] i_dbus_rdt[11] i_dbus_rdt[12]
+ i_dbus_rdt[13] i_dbus_rdt[14] i_dbus_rdt[15] i_dbus_rdt[16] i_dbus_rdt[17] i_dbus_rdt[18]
+ i_dbus_rdt[19] i_dbus_rdt[1] i_dbus_rdt[20] i_dbus_rdt[21] i_dbus_rdt[22] i_dbus_rdt[23]
+ i_dbus_rdt[24] i_dbus_rdt[25] i_dbus_rdt[26] i_dbus_rdt[27] i_dbus_rdt[28] i_dbus_rdt[29]
+ i_dbus_rdt[2] i_dbus_rdt[30] i_dbus_rdt[31] i_dbus_rdt[3] i_dbus_rdt[4] i_dbus_rdt[5]
+ i_dbus_rdt[6] i_dbus_rdt[7] i_dbus_rdt[8] i_dbus_rdt[9] i_ext_rd[0] i_ext_rd[10]
+ i_ext_rd[11] i_ext_rd[12] i_ext_rd[13] i_ext_rd[14] i_ext_rd[15] i_ext_rd[16] i_ext_rd[17]
+ i_ext_rd[18] i_ext_rd[19] i_ext_rd[1] i_ext_rd[20] i_ext_rd[21] i_ext_rd[22] i_ext_rd[23]
+ i_ext_rd[24] i_ext_rd[25] i_ext_rd[26] i_ext_rd[27] i_ext_rd[28] i_ext_rd[29] i_ext_rd[2]
+ i_ext_rd[30] i_ext_rd[31] i_ext_rd[3] i_ext_rd[4] i_ext_rd[5] i_ext_rd[6] i_ext_rd[7]
+ i_ext_rd[8] i_ext_rd[9] i_ext_ready i_ibus_ack i_ibus_rdt[0] i_ibus_rdt[10] i_ibus_rdt[11]
+ i_ibus_rdt[12] i_ibus_rdt[13] i_ibus_rdt[14] i_ibus_rdt[15] i_ibus_rdt[16] i_ibus_rdt[17]
+ i_ibus_rdt[18] i_ibus_rdt[19] i_ibus_rdt[1] i_ibus_rdt[20] i_ibus_rdt[21] i_ibus_rdt[22]
+ i_ibus_rdt[23] i_ibus_rdt[24] i_ibus_rdt[25] i_ibus_rdt[26] i_ibus_rdt[27] i_ibus_rdt[28]
+ i_ibus_rdt[29] i_ibus_rdt[2] i_ibus_rdt[30] i_ibus_rdt[31] i_ibus_rdt[3] i_ibus_rdt[4]
+ i_ibus_rdt[5] i_ibus_rdt[6] i_ibus_rdt[7] i_ibus_rdt[8] i_ibus_rdt[9] i_rst i_timer_irq
+ o_dbus_adr[10] o_dbus_adr[11] o_dbus_adr[12] o_dbus_adr[13] o_dbus_adr[14] o_dbus_adr[15]
+ o_dbus_adr[16] o_dbus_adr[17] o_dbus_adr[18] o_dbus_adr[19] o_dbus_adr[1] o_dbus_adr[20]
+ o_dbus_adr[21] o_dbus_adr[22] o_dbus_adr[23] o_dbus_adr[24] o_dbus_adr[25] o_dbus_adr[26]
+ o_dbus_adr[27] o_dbus_adr[28] o_dbus_adr[29] o_dbus_adr[2] o_dbus_adr[30] o_dbus_adr[31]
+ o_dbus_adr[3] o_dbus_adr[4] o_dbus_adr[5] o_dbus_adr[6] o_dbus_adr[7] o_dbus_adr[8]
+ o_dbus_adr[9] o_dbus_cyc o_dbus_dat[0] o_dbus_dat[10] o_dbus_dat[11] o_dbus_dat[12]
+ o_dbus_dat[13] o_dbus_dat[14] o_dbus_dat[15] o_dbus_dat[16] o_dbus_dat[17] o_dbus_dat[18]
+ o_dbus_dat[19] o_dbus_dat[1] o_dbus_dat[20] o_dbus_dat[21] o_dbus_dat[22] o_dbus_dat[23]
+ o_dbus_dat[24] o_dbus_dat[25] o_dbus_dat[26] o_dbus_dat[27] o_dbus_dat[28] o_dbus_dat[29]
+ o_dbus_dat[2] o_dbus_dat[30] o_dbus_dat[31] o_dbus_dat[3] o_dbus_dat[4] o_dbus_dat[5]
+ o_dbus_dat[6] o_dbus_dat[7] o_dbus_dat[8] o_dbus_dat[9] o_dbus_sel[0] o_dbus_sel[1]
+ o_dbus_sel[2] o_dbus_sel[3] o_dbus_we o_ext_funct3[0] o_ext_funct3[1] o_ext_funct3[2]
+ o_ext_rs1[0] o_ext_rs1[10] o_ext_rs1[11] o_ext_rs1[12] o_ext_rs1[13] o_ext_rs1[14]
+ o_ext_rs1[15] o_ext_rs1[16] o_ext_rs1[17] o_ext_rs1[18] o_ext_rs1[19] o_ext_rs1[1]
+ o_ext_rs1[20] o_ext_rs1[21] o_ext_rs1[22] o_ext_rs1[23] o_ext_rs1[24] o_ext_rs1[25]
+ o_ext_rs1[26] o_ext_rs1[27] o_ext_rs1[28] o_ext_rs1[29] o_ext_rs1[2] o_ext_rs1[30]
+ o_ext_rs1[31] o_ext_rs1[3] o_ext_rs1[4] o_ext_rs1[5] o_ext_rs1[6] o_ext_rs1[7] o_ext_rs1[8]
+ o_ext_rs1[9] o_ext_rs2[0] o_ext_rs2[10] o_ext_rs2[11] o_ext_rs2[12] o_ext_rs2[13]
+ o_ext_rs2[14] o_ext_rs2[15] o_ext_rs2[16] o_ext_rs2[17] o_ext_rs2[18] o_ext_rs2[19]
+ o_ext_rs2[1] o_ext_rs2[20] o_ext_rs2[21] o_ext_rs2[22] o_ext_rs2[23] o_ext_rs2[24]
+ o_ext_rs2[25] o_ext_rs2[26] o_ext_rs2[27] o_ext_rs2[28] o_ext_rs2[29] o_ext_rs2[2]
+ o_ext_rs2[30] o_ext_rs2[31] o_ext_rs2[3] o_ext_rs2[4] o_ext_rs2[5] o_ext_rs2[6]
+ o_ext_rs2[7] o_ext_rs2[8] o_ext_rs2[9] o_ibus_adr[0] o_ibus_adr[10] o_ibus_adr[11]
+ o_ibus_adr[12] o_ibus_adr[13] o_ibus_adr[14] o_ibus_adr[15] o_ibus_adr[16] o_ibus_adr[17]
+ o_ibus_adr[18] o_ibus_adr[19] o_ibus_adr[1] o_ibus_adr[20] o_ibus_adr[21] o_ibus_adr[22]
+ o_ibus_adr[23] o_ibus_adr[24] o_ibus_adr[25] o_ibus_adr[26] o_ibus_adr[27] o_ibus_adr[28]
+ o_ibus_adr[29] o_ibus_adr[2] o_ibus_adr[30] o_ibus_adr[31] o_ibus_adr[3] o_ibus_adr[4]
+ o_ibus_adr[5] o_ibus_adr[6] o_ibus_adr[7] o_ibus_adr[8] o_ibus_adr[9] o_ibus_cyc
+ vdd vss o_mdu_valid o_dbus_adr[0]
XFILLER_0_59_1220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09523__A2 net45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05903_ rf_ram.memory\[82\]\[0\] _01652_ _01654_ rf_ram.memory\[83\]\[0\] _01715_
+ rf_ram.memory\[81\]\[0\] _02099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_06883_ _02750_ _02811_ _02983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_09671_ net1 net27 _04755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_98_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06337__A2 _01755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08622_ _04058_ _04085_ _04086_ _00729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05834_ rf_ram.memory\[222\]\[0\] _01501_ _02030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_118_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05545__B1 _01688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05765_ rf_ram.memory\[154\]\[0\] _01958_ _01959_ rf_ram.memory\[155\]\[0\] _01960_
+ _01961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_08553_ net249 _03158_ _04042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11633__I net83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07504_ rf_ram.memory\[363\]\[0\] _03377_ _03378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_159_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08484_ rf_ram.memory\[379\]\[0\] _03995_ _03996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06727__I _02819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05696_ rf_ram.memory\[390\]\[0\] _01777_ _01773_ rf_ram.memory\[391\]\[0\] _01848_
+ rf_ram.memory\[389\]\[0\] _01892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_49_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_64_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07435_ rf_ram.memory\[332\]\[0\] _03334_ _03335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_64_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09039__A1 _04334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_135_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_21_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_135_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07366_ _03289_ _03290_ _03291_ _00268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_162_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_165_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06317_ rf_ram.memory\[182\]\[1\] _01631_ _01505_ _02512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09105_ rf_ram.memory\[95\]\[1\] _04384_ _04386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05787__B _01923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07297_ _03222_ _03247_ _03248_ _00242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_116_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09036_ rf_ram.memory\[105\]\[0\] _04343_ _04344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_14_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_96_2181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06248_ _02440_ _02442_ _01928_ _02443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_14_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_4_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_142_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06179_ _02370_ _02371_ _02372_ _02373_ _01670_ _02374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XANTENNA__09211__A1 _04431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_57_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_57_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_1000 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09762__A2 _04766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_1133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09938_ _04921_ _04926_ _04928_ _01204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_42_1290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_70_1697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09869_ _04884_ _04885_ _04886_ _01177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07525__A1 _02752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06328__A2 _01537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_1206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_29_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_178_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_166_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10713_ _00457_ clknet_leaf_131_clk rf_ram.memory\[42\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_113_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_165_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_153_3230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_180_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10644_ _00388_ clknet_leaf_107_clk rf_ram.memory\[383\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_153_3241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10575_ _00319_ clknet_leaf_169_clk rf_ram.memory\[324\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_134_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06264__A1 _01674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_77_1829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_114_2513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_114_2524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_146_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06016__A1 _01351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09753__A2 _04766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_1099 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_311_clk_I clknet_5_5__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07764__A1 _03521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11127_ _00863_ clknet_leaf_72_clk rf_ram.memory\[117\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05716__I _01626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11058_ _00795_ clknet_leaf_10_clk rf_ram.memory\[139\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_155_1318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06319__A2 _01922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10009_ rf_ram.memory\[277\]\[1\] _04970_ _04972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_326_clk_I clknet_5_4__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_188_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_149_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09269__A1 cpu.genblk3.csr.o_new_irq vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05550_ _01563_ _01746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_47_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_173_3606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_1194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05481_ _01633_ _01677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_15_1178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_157_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07220_ _03193_ _03198_ _03200_ _00213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_15_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_184_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_132_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07151_ _03013_ _03157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_42_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06102_ rf_ram.memory\[274\]\[1\] _01623_ _01625_ rf_ram.memory\[275\]\[1\] _02296_
+ _02297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_14_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_89_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07082_ _02781_ _02911_ _03114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_140_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_125_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06033_ rf_ram.memory\[574\]\[1\] _01502_ _01505_ _02228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_188_3882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_188_3893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_140_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11628__I net78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_35_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_35_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06231__B _01504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07984_ _03672_ _02866_ _03676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_52_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09723_ _04793_ _01123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06935_ _03018_ _03015_ _03019_ _00109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07507__A1 _03360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09654_ net109 _04737_ _04738_ _04740_ _04741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06866_ _02971_ _02972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__07841__I _03355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08605_ _04058_ _04074_ _04075_ _00723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05817_ rf_ram.memory\[178\]\[0\] _01856_ _01911_ rf_ram.memory\[179\]\[0\] _01931_
+ rf_ram.memory\[177\]\[0\] _02013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_09585_ _04651_ _04696_ _04697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06797_ rf_ram.memory\[50\]\[0\] _02924_ _02925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06191__B1 _01786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_1250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05748_ rf_ram.memory\[418\]\[0\] _01662_ _01646_ rf_ram.memory\[419\]\[0\] _01645_
+ rf_ram.memory\[417\]\[0\] _01944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_38_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08536_ _02865_ _03945_ _04031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_78_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_182_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05679_ rf_ram.memory\[450\]\[0\] _01801_ _01646_ rf_ram.memory\[451\]\[0\] _01810_
+ rf_ram.memory\[449\]\[0\] _01875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_147_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08467_ _03981_ _03982_ _03983_ _03984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_92_423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_108_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08483__A2 _03496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_98_2210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_162_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06494__A1 _01371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_98_2221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_174_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07418_ _02866_ _03101_ _03324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08398_ rf_ram.memory\[17\]\[1\] _03933_ _03935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_5_31__f_clk_I clknet_3_7_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07349_ rf_ram.memory\[26\]\[0\] _03280_ _03281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_116_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_59_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_162_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10360_ _00104_ clknet_leaf_133_clk rf_ram.memory\[298\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07994__A1 _03672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09019_ rf_ram.memory\[108\]\[0\] _04332_ _04333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10291_ _00035_ clknet_leaf_318_clk rf_ram.memory\[525\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_66_1098 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_1217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_72_1737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07746__A1 _03524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_38_1112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_1123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_1134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_107_2383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_1178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_107_2394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_158_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_69_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_96_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09671__A1 net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_153_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_84_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05288__A2 _01341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06485__A1 rf_ram.memory\[4\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_181_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10627_ _00371_ clknet_leaf_114_clk rf_ram.memory\[406\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_148_1144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08226__A2 _03135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_183_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_153_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06237__A1 _01768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_1075 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10033__A2 _02815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_1139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10558_ _00302_ clknet_leaf_158_clk rf_ram.memory\[330\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_161_1322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06788__A2 _02917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10489_ _00233_ clknet_leaf_46_clk rf_ram.memory\[193\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_250_clk_I clknet_5_20__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_166_3476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05748__B1 _01646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_166_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06051__B _01629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_16_Left_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05212__A2 _01411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_183_3790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_159_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_leaf_265_clk_I clknet_5_17__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_127_2748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_127_2759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06720_ _02797_ _02867_ _02868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_56_1223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08162__A1 net237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06651_ rf_ram.memory\[346\]\[1\] _02816_ _02818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_95_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06173__B1 _01654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06712__A2 _02846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_188_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05602_ rf_ram.memory\[308\]\[0\] _01709_ _01715_ rf_ram.memory\[309\]\[0\] _01713_
+ rf_ram.memory\[311\]\[0\] _01798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_149_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09370_ net207 _04549_ _04552_ net208 _04557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06582_ cpu.immdec.imm11_7\[2\] _02730_ _02763_ _02764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_8_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05533_ _01349_ _01718_ _01728_ _01729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_08321_ _03884_ _03885_ _03886_ _00628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_157_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08465__A2 net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_25_Left_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08252_ rf_ram.memory\[527\]\[0\] _03843_ _03844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_89_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05464_ _01599_ _01660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_12
XFILLER_0_156_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_203_clk_I clknet_5_24__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_670 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07203_ _03161_ _03187_ _03189_ _00207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_172_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_160_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_31_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08183_ _03790_ _03799_ _03801_ _00575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05395_ _01587_ _01588_ _01589_ _01590_ _01564_ _01591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__09414__A1 _04463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_31_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07134_ rf_ram.memory\[486\]\[1\] _03145_ _03147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_125_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_160_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_43_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07065_ rf_ram.memory\[375\]\[1\] _03102_ _03104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_101_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_218_clk_I clknet_5_22__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput220 net220 o_ibus_adr[26] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_100_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput231 net231 o_ibus_adr[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_64_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06016_ _01351_ _02199_ _02210_ _01569_ _02211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_54_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05451__A2 _01644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_54_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_34_Left_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_26_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05356__I _01551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input36_I i_ibus_rdt[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_1313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07967_ _02921_ _02954_ _03665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06951__A2 _02829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09706_ _04739_ _04781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_06918_ _02975_ _03004_ _03006_ _00105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07898_ rf_ram.memory\[461\]\[1\] _03620_ _03623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08153__A1 _03754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09637_ _04524_ net61 _04727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_97_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06849_ _02958_ _02960_ _02961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_35_1318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07900__A1 _02839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09568_ _03992_ cpu.immdec.imm30_25\[3\] _04684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_139_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_43_Left_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_93_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08519_ _02838_ _03949_ _04020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_176_970 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09499_ _04633_ _01059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_37_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_851 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_92_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_102_2291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11530_ _01262_ clknet_leaf_205_clk rf_ram.memory\[30\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_147_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05959__C rf_ram.i_raddr\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_137_Right_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_11461_ _01193_ clknet_leaf_137_clk rf_ram.memory\[292\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_18_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10412_ _00156_ clknet_leaf_182_clk rf_ram.memory\[494\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_116_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11392_ _01124_ clknet_leaf_225_clk net106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__07967__A1 _02921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10343_ _00087_ clknet_leaf_178_clk rf_ram.memory\[283\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_131_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05978__B1 _01655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_21_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_52_Left_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_104_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_1063 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10274_ _00018_ clknet_leaf_276_clk rf_ram.memory\[235\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07719__A1 _03491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_148_3140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_1171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_148_3151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_1223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08392__A1 _03919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_109_2423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_1289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_161_3384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06155__B1 _01678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_17_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_61_Left_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_17_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_122_2656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_122_2667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_173_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_145_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09644__A1 cpu.mem_bytecnt\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_1164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_138_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10254__A2 _03035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_104_Right_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_71_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11659_ net110 net182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_114_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10006__A2 _03072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05180_ cpu.decode.opcode\[2\] _01380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_25_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_168_3505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_168_3516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05885__B _01928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06630__A1 _02795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_3_1_0_clk clknet_0_clk clknet_3_1_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_185_3830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_1244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_1255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08870_ rf_ram.memory\[130\]\[1\] _04239_ _04241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_32_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_181_3749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07821_ _02761_ _03234_ _03575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_19_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_84_clk_I clknet_5_10__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07752_ _02781_ _03481_ _03532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08135__A1 _03757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06703_ rf_ram.memory\[522\]\[0\] _02856_ _02857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06146__B1 _01725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07683_ _02908_ _03390_ _03489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09883__A1 _04884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09422_ _04586_ _01029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_17_1026 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06697__A1 _02781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06634_ _02748_ _02802_ _02804_ _00023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_leaf_99_clk_I clknet_5_14__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09353_ _04547_ _00999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09635__A1 _04524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_47_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06565_ _02739_ _02748_ _02749_ _00009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_19_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_47_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11641__I net120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_142_clk_I clknet_5_27__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08304_ rf_ram.memory\[221\]\[0\] _03875_ _03876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06449__A1 _01903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05516_ rf_ram.memory\[320\]\[0\] _01711_ _01602_ _01712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_63_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09284_ _01485_ _04504_ _04505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06496_ _01376_ _02690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_0_117_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_22_clk_I clknet_5_3__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08235_ _03823_ _03831_ _03833_ _00595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_74_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05447_ _01508_ _01643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_90_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_144_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05672__A2 _01709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_1100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08166_ rf_ram.memory\[544\]\[1\] _03788_ _03791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05378_ rf_ram.memory\[554\]\[0\] _01532_ _01521_ rf_ram.memory\[555\]\[0\] _01517_
+ rf_ram.memory\[553\]\[0\] _01574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XANTENNA_clkbuf_leaf_157_clk_I clknet_5_26__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_120_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07117_ rf_ram.memory\[500\]\[0\] _03136_ _03137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08097_ _03724_ _03745_ _03747_ _00543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08610__A2 _04078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_37_clk_I clknet_5_7__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07048_ rf_ram.memory\[391\]\[1\] _03090_ _03093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_63_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08374__A1 net245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10181__A1 _05049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08999_ _04298_ _04319_ _04320_ _00872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_177_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08126__A1 _02829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_3_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06137__B1 _01778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_97_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10961_ _00698_ clknet_leaf_65_clk rf_ram.memory\[69\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08677__A2 _03765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_104_2331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_151_1310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_67_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_168_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_168_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10892_ _00636_ clknet_leaf_303_clk rf_ram.memory\[214\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_66_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_156_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_84_1961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_183_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09626__A1 _04643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06645__I _02812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_182_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09021__I _04061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11513_ _01245_ clknet_leaf_197_clk rf_ram.memory\[506\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_110_1073 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05663__A2 _01856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09929__A2 _03072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_1200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08860__I _04057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11444_ _01176_ clknet_leaf_293_clk rf_ram.memory\[5\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_124_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_149_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_33_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_0_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11375_ _01107_ clknet_leaf_233_clk net98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_150_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_132_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05415__A2 _01606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10326_ _00070_ clknet_leaf_122_clk rf_ram.memory\[290\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_163_3413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10257_ rf_ram.memory\[9\]\[1\] _05122_ _05124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_163_3424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08365__A1 _03884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10188_ _05081_ _05079_ _05082_ _01300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06376__B1 _01793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_124_2707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08117__A1 _03754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09865__A1 _04840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_88_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_1160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_186_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05351__A1 _01495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09617__A1 _04637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_186_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_158_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06350_ _02541_ _02542_ _02543_ _02544_ _01717_ _02545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_139_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05301_ rf_ram.i_raddr\[1\] _01497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_139_2972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_139_2983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06281_ _01951_ _02474_ _02475_ _02476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
Xclkbuf_leaf_150_clk clknet_5_26__leaf_clk clknet_leaf_150_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_142_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08840__A2 _04195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08020_ _02822_ _03693_ _03700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05232_ cpu.immdec.imm24_20\[0\] _01432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_71_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06851__A1 _02927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_42_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_130_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_987 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05163_ _01364_ _01365_ _01366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_25_1317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06603__A1 _01496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09971_ _04918_ _04947_ _04948_ _01217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_126_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08922_ rf_ram.memory\[389\]\[1\] _04271_ _04273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_23_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07159__A2 _02946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08853_ rf_ram.memory\[132\]\[1\] _04228_ _04230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_97_1142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07804_ rf_ram.memory\[435\]\[1\] _03563_ _03565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_174_1321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08784_ _04167_ _04186_ _04187_ _00790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_98_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05996_ rf_ram.memory\[520\]\[1\] _01524_ _01528_ _02191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_27_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_0_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07735_ _03355_ _03521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_0_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_49_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06119__B1 _01668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09856__A1 cpu.state.genblk1.misalign_trap_sync_r vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07666_ _02866_ _03089_ _03478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_95_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_177_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09405_ _04575_ _01023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06617_ _02743_ _02789_ _02790_ _00020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_48_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09608__A1 net249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07597_ _03425_ _03433_ _03435_ _00355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_133_1073 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09459__I1 net80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_9_Left_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_137_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09336_ rf_ram.memory\[99\]\[1\] _04536_ _04538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06548_ _01353_ _01358_ _02733_ _01341_ _02734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XTAP_TAPCELL_ROW_62_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_164_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_146_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_146_984 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09267_ cpu.genblk3.csr.mcause31 _04492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xclkbuf_leaf_141_clk clknet_5_27__leaf_clk clknet_leaf_141_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_06479_ rf_ram.memory\[14\]\[1\] _01640_ _01503_ _02674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_173_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08218_ _03689_ _03823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__05645__A2 _01644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09198_ _04434_ _04442_ _04444_ _00947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_161_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08149_ rf_ram.memory\[547\]\[1\] _03778_ _03780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_43_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09631__I1 net58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08595__A1 _04058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11160_ _00896_ clknet_leaf_66_clk rf_ram.memory\[100\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_105_1142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10111_ rf_ram.memory\[392\]\[0\] _05034_ _05035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11091_ _00828_ clknet_leaf_98_clk rf_ram.memory\[419\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06070__A2 _01677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_8_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_max_cap236_I _02922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10042_ _04985_ _04990_ _04992_ _01244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_output67_I net67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10154__A1 _05046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06358__B1 _01959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08898__A2 _04257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_141_3007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_141_3018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_188_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_wire239_I _02893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09847__A1 _01382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_1070 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10944_ _00682_ clknet_leaf_103_clk rf_ram.memory\[379\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_39_1092 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_129_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05869__C1 _01702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10875_ _00619_ clknet_leaf_35_clk rf_ram.memory\[203\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_168_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_151_1184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_155_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10209__A2 _03547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05884__A2 _01808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_156_3283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07086__A1 _03092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_171_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_164_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_156_3294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_132_clk clknet_5_24__leaf_clk clknet_leaf_132_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_152_921 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09686__I _04766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06833__A1 _02930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_117_2566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_117_2577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_5 _01804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11427_ _01159_ clknet_leaf_212_clk rf_ram.memory\[249\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_151_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_134_2880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05719__I _01536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_134_2891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08586__A1 _04062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_50_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11358_ _01090_ clknet_leaf_22_clk rf_ram.memory\[72\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_162_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10309_ _00053_ clknet_leaf_271_clk rf_ram.memory\[516\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11289_ _01024_ clknet_leaf_249_clk net226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__08338__A1 _03884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06349__B1 _01811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_199_clk clknet_5_25__leaf_clk clknet_leaf_199_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_20_1247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_174_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05850_ _01674_ _02033_ _02045_ _01362_ _02046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__05454__I _01601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07561__A2 _02917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_156_1051 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_178_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05781_ rf_ram.memory\[130\]\[0\] _01606_ _01608_ rf_ram.memory\[131\]\[0\] _01610_
+ rf_ram.memory\[129\]\[0\] _01977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_156_1073 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07520_ _03356_ _03386_ _03387_ _00326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_77_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_1023 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_1165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_174_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07451_ _03323_ _03343_ _03344_ _00300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_176_3659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_146_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06402_ rf_ram.memory\[86\]\[1\] _01785_ _01707_ _02597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_45_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07382_ _03289_ _03300_ _03301_ _00274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_128_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09121_ _04367_ _04393_ _04395_ _00919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07077__A1 _02788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06333_ rf_ram.memory\[217\]\[1\] _01515_ _02528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
Xclkbuf_leaf_123_clk clknet_5_13__leaf_clk clknet_leaf_123_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_155_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_72_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_40_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06824__A1 _02927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06264_ _01674_ _02447_ _02458_ _01569_ _02459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_60_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09052_ _04331_ _04352_ _04353_ _00892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05627__A2 _01687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_1120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05215_ cpu.immdec.imm11_7\[0\] cpu.immdec.imm24_20\[0\] _01414_ _01415_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_53_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08003_ _03686_ _03687_ _03688_ _00508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_13_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06195_ _01769_ _02388_ _02389_ _02390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_142_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xmax_cap241 _02882_ net241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_64_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08577__A1 _04026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05146_ _01348_ _01349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_29_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_1147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06052__A2 _01631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09954_ _04911_ _02946_ _04938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_5_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08329__A1 _03887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08905_ rf_ram.memory\[126\]\[1\] _04260_ _04262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10136__A1 _05049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09264__C _02713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09885_ _04887_ _04893_ _04895_ _01184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_57_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07001__A1 _03053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08836_ rf_ram.memory\[469\]\[0\] _04219_ _04220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_174_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08767_ _02945_ _04152_ _04177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09829__A1 _04837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05979_ rf_ram.memory\[10\]\[0\] _01686_ _01525_ _02175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_169_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07718_ rf_ram.memory\[380\]\[1\] _03509_ _03511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09280__B cpu.genblk3.csr.o_new_irq vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_1243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08698_ _04129_ _04131_ _04133_ _00758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_71_1134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07649_ rf_ram.memory\[405\]\[1\] _03466_ _03468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_output105_I net105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_24_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05866__A2 _01989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10660_ _00404_ clknet_leaf_129_clk rf_ram.memory\[37\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_94_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_165_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09319_ _04526_ net35 _04521_ cpu.immdec.imm11_7\[4\] _04522_ cpu.immdec.imm11_7\[3\]
+ _04528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_106_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10591_ _00335_ clknet_leaf_165_clk rf_ram.memory\[320\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_114_clk clknet_5_15__leaf_clk clknet_leaf_114_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_106_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_90_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_181_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_79_1860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_161_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_151_3191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_79_1871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05539__I _01536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08568__A1 net247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_146_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09765__B1 _04760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11212_ _00948_ clknet_leaf_65_clk rf_ram.memory\[70\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_102_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07240__A1 _03193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_1258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11143_ _00879_ clknet_leaf_35_clk rf_ram.memory\[10\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_112_2474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_112_2485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput75 net75 o_dbus_adr[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput86 net86 o_dbus_adr[29] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput97 net97 o_dbus_cyc vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__10127__A1 _05014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11074_ _00811_ clknet_leaf_54_clk rf_ram.memory\[469\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10025_ _04953_ _04979_ _04981_ _01238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08740__A1 _04157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06200__C1 _01726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05554__A1 _01603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_1078 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_188_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_187_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_158_3323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_158_3334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10927_ _00671_ clknet_leaf_8_clk rf_ram.memory\[174\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06319__B _01923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10858_ _00602_ clknet_leaf_315_clk rf_ram.memory\[527\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_128_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_186_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_119_2606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07059__A1 _03092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_105_clk clknet_5_15__leaf_clk clknet_leaf_105_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_136_2920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10789_ _00533_ clknet_leaf_323_clk rf_ram.memory\[562\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_81_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_136_2931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_171_3567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_171_3578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_147_1039 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_5_17__f_clk clknet_3_4_0_clk clknet_5_17__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_48_1114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05877__C _01569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_132_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05449__I _01609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_10_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09756__B1 _04760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_5_8__f_clk_I clknet_3_2_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_495 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07231__A1 _02829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06034__A2 _01538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06951_ _02766_ _02829_ _03029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_94_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05902_ rf_ram.memory\[80\]\[0\] _01863_ _01602_ _02098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_158_1146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09670_ net124 _04737_ _04753_ _04739_ _04754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_158_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_59_1232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06882_ _02975_ _02980_ _02982_ _00093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_94_1123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08621_ rf_ram.memory\[529\]\[0\] _04085_ _04086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_27_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_20_1099 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05833_ _02026_ _02028_ _01928_ _02029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_179_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08552_ _04026_ _04039_ _04041_ _00704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05764_ rf_ram.memory\[153\]\[0\] _01515_ _01960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_76_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07503_ _02781_ _03101_ _03377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_175_810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08483_ net244 _03496_ _03995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_175_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05695_ rf_ram.memory\[388\]\[0\] _01846_ _01891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_119_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07434_ _02788_ _02815_ _03334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_147_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_1065 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_21_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_57_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_175_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_130_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07365_ rf_ram.memory\[251\]\[0\] _03290_ _03291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_128_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08798__A1 _02787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09104_ _04364_ _04384_ _04385_ _00912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06316_ _02507_ _02508_ _02509_ _02510_ _01860_ _02511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XPHY_EDGE_ROW_99_Left_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_33_738 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07296_ rf_ram.memory\[25\]\[0\] _03247_ _03248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_26_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_1247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09035_ net249 _04339_ _04343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_116_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06273__A2 _01958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_1209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_1258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_96_2182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06247_ rf_ram.memory\[442\]\[1\] _01719_ _01925_ rf_ram.memory\[443\]\[1\] _02441_
+ _02442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_170_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_946 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05359__I _01516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input66_I i_timer_irq vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06178_ rf_ram.memory\[498\]\[1\] _01500_ _01763_ rf_ram.memory\[499\]\[1\] _01668_
+ rf_ram.memory\[497\]\[1\] _02373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_13_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_57_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_57_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06025__A2 _01544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05129_ cpu.decode.op21 _01331_ _01332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__05295__S _01491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08970__A1 _04301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06430__C1 _01696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09937_ rf_ram.memory\[340\]\[1\] _04926_ _04928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10109__A1 _05017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09868_ rf_ram.memory\[60\]\[0\] _04885_ _04886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07525__A2 _03390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_70_1698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08819_ _04205_ _04207_ _04209_ _00803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_29_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09799_ _04837_ _04842_ _04843_ _01149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_29_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_185_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_185_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07289__A1 _03225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_178_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05839__A2 _01649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10712_ _00456_ clknet_leaf_134_clk rf_ram.memory\[42\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_165_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_82_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10643_ _00387_ clknet_leaf_96_clk rf_ram.memory\[402\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_153_3231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_153_3242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08789__A1 _04167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06653__I _02742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_181_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10574_ _00318_ clknet_leaf_169_clk rf_ram.memory\[324\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_106_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_114_2514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07461__A1 _03323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07213__A1 _03190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08961__A1 _04266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06421__C1 _01786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11126_ _00862_ clknet_leaf_72_clk rf_ram.memory\[117\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_1320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06321__C _01978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11057_ _00794_ clknet_leaf_10_clk rf_ram.memory\[139\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08713__A1 _04129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_129_2790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10008_ _04950_ _04970_ _04971_ _01231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06828__I _02945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05732__I _01563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_188_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_8_1247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_1271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_326_clk clknet_5_4__leaf_clk clknet_leaf_326_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_47_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_173_3607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_157_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05480_ rf_ram.memory\[350\]\[0\] _01543_ _01676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_74_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_15_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_144_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_156_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06563__I _02747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07150_ _03126_ _03154_ _03156_ _00187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_54_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06101_ rf_ram.memory\[273\]\[1\] _01626_ _02296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__06255__A2 _01808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07081_ _03092_ _03111_ _03113_ _00161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_125_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_180_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_152_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06032_ _02223_ _02224_ _02225_ _02226_ _01494_ _02227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_23_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_61_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_188_3883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_188_3894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06007__A2 _01511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_1275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_1128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_91_2090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_35_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_35_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07983_ _03654_ _03673_ _03675_ _00501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09722_ net105 _04790_ _04791_ net106 _04792_ _04793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XTAP_TAPCELL_ROW_52_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06934_ rf_ram.memory\[297\]\[1\] _03015_ _03019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_52_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08704__A1 _02991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09653_ _04739_ _04740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_06865_ _02773_ _02786_ _02971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_08604_ rf_ram.memory\[164\]\[0\] _04074_ _04075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_59_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05816_ rf_ram.memory\[176\]\[0\] _01922_ _01923_ _02012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_96_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_145_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09584_ _04477_ cpu.immdec.imm24_20\[1\] _04696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06796_ _02921_ _02923_ _02924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_78_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_179_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_78_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_167_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_132_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_118_Right_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_78_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08535_ _04026_ _04028_ _04030_ _00698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05747_ rf_ram.memory\[416\]\[0\] _01755_ _01756_ _01943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xclkbuf_leaf_317_clk clknet_5_5__leaf_clk clknet_leaf_317_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_132_1149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08466_ cpu.state.init_done _01364_ _02709_ _03983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_64_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05678_ rf_ram.memory\[448\]\[0\] _01649_ _01756_ _01874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_147_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_98_2211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07417_ _03013_ _03323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__07691__A1 _03488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_98_2222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_162_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08397_ _03919_ _03933_ _03934_ _00656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_46_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07348_ _02813_ _02997_ _03280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_33_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_59_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06406__C _01670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06246__A2 _01918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07443__A1 _03326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07279_ _03225_ _03235_ _03237_ _00235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_103_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_60_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_1077 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09018_ _02787_ _04303_ _04332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07994__A2 _02923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output172_I net172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10290_ _00034_ clknet_leaf_314_clk rf_ram.memory\[525\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_143_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09196__A1 _04431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_1217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08943__A1 _04269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06403__C1 _01763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_87_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_1037 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_107_2384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_150_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_308_clk clknet_5_5__leaf_clk clknet_leaf_308_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_84_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06485__A2 _01643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_181_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_154_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_153_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05693__B1 _01786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_64_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10626_ _00370_ clknet_leaf_114_clk rf_ram.memory\[406\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_107_740 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06316__C _01860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07434__A1 _02788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10557_ _00301_ clknet_leaf_148_clk rf_ram.memory\[368\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_10_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_52_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_1286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10488_ _00232_ clknet_leaf_45_clk rf_ram.memory\[193\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06332__B _01551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05727__I _01550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08934__A1 _02953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_166_3477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_1053 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11109_ _00845_ clknet_leaf_85_clk rf_ram.memory\[124\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_75_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_183_3791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_127_2749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_1183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08162__A2 _03765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_182_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06650_ _02743_ _02816_ _02817_ _00026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_177_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_1208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_177_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05462__I _01563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05601_ rf_ram.memory\[310\]\[0\] _01719_ _01707_ _01797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05381__C1 _01540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06581_ _02732_ _02762_ _02763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__05920__A1 _01909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09111__A1 _04367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08320_ rf_ram.memory\[242\]\[0\] _03885_ _03886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05532_ _01720_ _01722_ _01723_ _01727_ _01658_ _01728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_129_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_1099 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_185_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_131_1160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08251_ _02845_ _02954_ _03843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_46_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06476__A2 _01633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05463_ _01651_ _01657_ _01658_ _01659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_43_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07202_ rf_ram.memory\[273\]\[1\] _03187_ _03189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08182_ rf_ram.memory\[541\]\[1\] _03799_ _03801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_171_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_31_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05394_ rf_ram.memory\[570\]\[0\] _01544_ _01540_ rf_ram.memory\[571\]\[0\] _01539_
+ rf_ram.memory\[569\]\[0\] _01590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_172_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_31_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06228__A2 _01755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07133_ _03123_ _03145_ _03146_ _00180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_15_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_1229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_93_2130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07064_ _03087_ _03102_ _03103_ _00154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_30_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput210 net210 o_ibus_adr[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XPHY_EDGE_ROW_12_Right_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_63_1239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05987__A1 _01348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput221 net221 o_ibus_adr[27] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_2_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11639__I net98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09178__A1 _03134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput232 net232 o_ibus_adr[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_06015_ _02204_ _02209_ _01351_ _02210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_54_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_54_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_103_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06400__A2 _01801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07966_ _03654_ _03662_ _03664_ _00495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09705_ _04780_ _01118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input29_I i_dbus_rdt[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06917_ rf_ram.memory\[298\]\[1\] _03004_ _03006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07897_ _03359_ _03622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xclkbuf_leaf_94_clk clknet_5_14__leaf_clk clknet_leaf_94_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09636_ _04524_ _01433_ _04726_ _01103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06848_ _02959_ _02960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XPHY_EDGE_ROW_21_Right_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_69_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_78_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07900__A2 _03547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09567_ _04683_ _01077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06779_ _02910_ _02911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_38_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09102__A1 _02908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08518_ _03956_ _04017_ _04019_ _00692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_72_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09498_ cpu.alu.cmp_r _04632_ _01491_ _04633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_72_1092 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_310_clk_I clknet_5_5__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_102_2292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_167_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08449_ net34 _03967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__06467__A2 _01682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_163_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11460_ _01192_ clknet_leaf_167_clk rf_ram.memory\[345\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_92_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07416__A1 _03292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06219__A2 _01785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10411_ _00155_ clknet_leaf_111_clk rf_ram.memory\[375\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_61_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_1318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11391_ _01123_ clknet_leaf_228_clk net105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XPHY_EDGE_ROW_30_Right_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_clkbuf_leaf_325_clk_I clknet_5_4__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_1306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07967__A2 _02954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10342_ _00086_ clknet_leaf_178_clk rf_ram.memory\[283\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_33_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05978__B2 rf_ram.memory\[13\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09169__A1 _04397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10273_ _00017_ clknet_leaf_261_clk rf_ram.memory\[234\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_148_3141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_148_3152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05991__B _02186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_109_2424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_1268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_161_3385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_85_clk clknet_5_10__leaf_clk clknet_leaf_85_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_69_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_17_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_122_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_185_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05363__C1 _01554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_122_2668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_1241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_1170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_56_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_167_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_1188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09644__A2 _01376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_166_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07655__A1 _03458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06458__A2 _01508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_154_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_153_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11658_ net108 net180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_154_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_181_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10609_ _00353_ clknet_leaf_156_clk rf_ram.memory\[355\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_153_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11589_ _01321_ clknet_leaf_302_clk rf_ram.memory\[213\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_52_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_168_3506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_168_3517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08080__A1 _03721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_185_3820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_185_3831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06630__A2 _02801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06062__B _01504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_1212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05457__I _01518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08907__A1 _02959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_1159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_32_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07820_ _03557_ _03572_ _03574_ _00439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09580__A1 _01391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06394__A1 _01972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07751_ _03524_ _03529_ _03531_ _00413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_leaf_76_clk clknet_5_10__leaf_clk clknet_leaf_76_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09332__A1 _04466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06702_ _02775_ _02846_ _02856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_56_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07682_ _03355_ _03488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_79_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09421_ net91 net92 _02707_ _04586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06633_ rf_ram.memory\[293\]\[1\] _02802_ _02804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07894__A1 _02836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06697__A2 _02846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_165_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09352_ net230 _03991_ _04540_ net231 _04547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06564_ rf_ram.memory\[200\]\[1\] _02739_ _02749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09635__A2 net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_47_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_158_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_47_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08303_ _03230_ _02960_ _03875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__07646__A1 _03071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05515_ _01613_ _01711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_117_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09283_ _01393_ _01340_ _04504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06495_ _01371_ _02235_ _02462_ _02689_ _00001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_75_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06237__B _02431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05657__B1 _01778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08234_ rf_ram.memory\[531\]\[1\] _03831_ _03833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05141__B cpu.state.genblk1.misalign_trap_sync_r vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05446_ rf_ram.memory\[382\]\[0\] _01641_ _01642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_145_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_173_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_160_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08165_ _03689_ _03790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_172_495 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05377_ rf_ram.memory\[552\]\[0\] _01524_ _01528_ _01573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_160_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_160_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07116_ _02915_ _03135_ _03136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_42_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08096_ rf_ram.memory\[557\]\[1\] _03745_ _03747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_63_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_1313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07047_ _03017_ _03092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_113_595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05367__I _01562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08374__A2 _03903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08998_ rf_ram.memory\[112\]\[0\] _04319_ _04320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_103_1092 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_138_1111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output135_I net135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07949_ _03359_ _03654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_143_3060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_67_clk clknet_5_8__leaf_clk clknet_leaf_67_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08126__A2 _03765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_3_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09323__A1 net243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_173_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_170_Right_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_3_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10960_ _00697_ clknet_leaf_65_clk rf_ram.memory\[69\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09874__A2 _01418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_67_1637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_104_2321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_168_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_67_1648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_104_2332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_151_1322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_1296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09619_ _04643_ _01333_ _04705_ _01093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07885__A1 _03587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05345__C1 _01540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10891_ _00635_ clknet_leaf_215_clk rf_ram.memory\[240\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_70_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_168_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_84_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_84_1962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05360__A2 _01501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_65_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_530 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_167_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06147__B _01650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11512_ _01244_ clknet_leaf_144_clk rf_ram.memory\[305\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_135_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_leaf_264_clk_I clknet_5_17__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11443_ _01175_ clknet_leaf_293_clk rf_ram.memory\[5\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_150_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_180_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_34_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_85_1272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08062__A1 net242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06661__I _02825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11374_ _01106_ clknet_leaf_61_clk rf_ram.memory\[78\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10325_ _00069_ clknet_leaf_123_clk rf_ram.memory\[291\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_104_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_1289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_279_clk_I clknet_5_17__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10256_ _02819_ _05122_ _05123_ _01327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_163_3414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_163_3425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_1170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10187_ rf_ram.memory\[190\]\[1\] _05079_ _05082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10172__A2 _03134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_202_clk_I clknet_5_25__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_124_2708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_58_clk clknet_5_9__leaf_clk clknet_leaf_58_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09314__A1 _04524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09314__B2 cpu.immdec.imm11_7\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_186_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_217_clk_I clknet_5_22__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_158_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_178_3690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07628__A1 _03425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_139_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_127_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05300_ rf_ram.i_raddr\[0\] _01496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_16_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_154_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_139_2973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06280_ rf_ram.memory\[150\]\[1\] _01940_ _01959_ rf_ram.memory\[151\]\[1\] _01968_
+ rf_ram.memory\[149\]\[1\] _02475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_0_127_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_139_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_182_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05231_ cpu.bufreg.i_sh_signed net134 _01405_ cpu.branch_op _01431_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_170_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_42_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_188_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_13_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05162_ cpu.genblk3.csr.o_new_irq _01340_ _01365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_110_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07800__A1 _03557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09970_ rf_ram.memory\[464\]\[0\] _04947_ _04948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_110_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08921_ _04266_ _04271_ _04272_ _00842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_62_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08852_ _04202_ _04228_ _04229_ _00816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07803_ _03554_ _03563_ _03564_ _00432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_88_2040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08783_ rf_ram.memory\[141\]\[0\] _04186_ _04187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05995_ rf_ram.memory\[524\]\[1\] _01511_ _01517_ rf_ram.memory\[525\]\[1\] _01521_
+ rf_ram.memory\[527\]\[1\] _02190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
Xclkbuf_leaf_49_clk clknet_5_12__leaf_clk clknet_leaf_49_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_58_1149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09305__A1 _04463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07734_ _03491_ _03518_ _03520_ _00407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_0_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_49_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09856__A2 _01413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07665_ _03458_ _03475_ _03477_ _00381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07867__A1 _03590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09404_ net225 _03990_ _04539_ net226 _04575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06616_ rf_ram.memory\[236\]\[0\] _02789_ _02790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_153_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07596_ rf_ram.memory\[315\]\[1\] _03433_ _03435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_149_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05650__I _01536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_530 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09608__A2 _04507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09122__I _02742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07619__A1 _02904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09335_ _04463_ _04536_ _04537_ _00991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06547_ _01352_ cpu.immdec.imm11_7\[1\] _02733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_118_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_80_Left_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09266_ _04480_ _04481_ _04491_ _00968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08292__A1 _03855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06478_ _02661_ _02665_ _02669_ _02672_ _02673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_16_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08217_ _03820_ _03821_ _03822_ _00588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_161_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05429_ _01624_ _01625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_12
XFILLER_0_16_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09197_ rf_ram.memory\[82\]\[1\] _04442_ _04444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_50_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_160_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08148_ _03754_ _03778_ _03779_ _00562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08044__A1 _03690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08079_ rf_ram.memory\[560\]\[0\] _03736_ _03737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_140_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10110_ net250 _03088_ _05034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05802__B1 _01520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11090_ _00827_ clknet_leaf_26_clk rf_ram.memory\[128\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_8_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_1180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_1142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09544__A1 _04478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10041_ rf_ram.memory\[305\]\[1\] _04990_ _04992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_41_1175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_141_3008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_141_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10943_ _00681_ clknet_leaf_255_clk cpu.state.ibus_cyc vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07858__A1 _02728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05869__B1 _01625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_565 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06656__I _02821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_3_0_0_clk clknet_0_clk clknet_3_0_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_10874_ _00618_ clknet_leaf_35_clk rf_ram.memory\[203\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05333__A2 _01524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05560__I _01601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_27_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_1200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_1209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_1282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_156_3284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08283__A1 _03230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_156_3295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10090__A1 _03445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_83_clk_I clknet_5_11__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_117_2567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08035__A1 _02991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11426_ _01158_ clknet_leaf_201_clk rf_ram.memory\[259\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_117_2578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_134_2881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06046__B1 _01608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_134_2892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11357_ _01089_ clknet_leaf_22_clk rf_ram.memory\[73\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_22_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_46_1075 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10308_ _00052_ clknet_leaf_271_clk rf_ram.memory\[516\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_98_clk_I clknet_5_14__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11288_ _01023_ clknet_leaf_248_clk net225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_141_clk_I clknet_5_27__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10239_ _02737_ _03071_ _05113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05735__I _01626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_21_clk_I clknet_5_3__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05557__C1 _01636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05780_ rf_ram.memory\[128\]\[0\] _01915_ _01923_ _01976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_156_1063 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_156_clk_I clknet_5_26__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_1144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07450_ rf_ram.memory\[368\]\[0\] _03343_ _03344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_53_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_36_clk_I clknet_5_6__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05470__I _01643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06401_ _02594_ _02595_ _01746_ _02596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_44_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07381_ rf_ram.memory\[266\]\[0\] _03300_ _03301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_17_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_146_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09120_ rf_ram.memory\[575\]\[1\] _04393_ _04395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_17_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06332_ rf_ram.memory\[216\]\[1\] _01537_ _01551_ _02527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_29_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07077__A2 _02911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10081__A1 _05014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_40_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09051_ rf_ram.memory\[102\]\[0\] _04352_ _04353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06263_ _01350_ _02452_ _02457_ _02458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_114_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_6_Right_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_13_600 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_143_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08002_ rf_ram.memory\[465\]\[0\] _03687_ _03688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_115_668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05214_ net134 _01395_ _01414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_130_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_170_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06194_ rf_ram.memory\[476\]\[1\] _01863_ _01848_ rf_ram.memory\[477\]\[1\] _01696_
+ rf_ram.memory\[479\]\[1\] _02389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_130_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_128_1165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_4_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09774__A1 _04637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xmax_cap242 _02865_ net242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_05145_ cpu.csr_imm _01346_ _01347_ _01348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_141_1310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xmax_cap253 _01568_ net253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_60_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_1137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09953_ _04921_ _04935_ _04937_ _01210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05260__A1 _01436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11647__I net128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_109_clk_I clknet_5_15__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09526__A1 _03967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08904_ _04234_ _04260_ _04261_ _00836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_110_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09884_ rf_ram.memory\[229\]\[1\] _04893_ _04895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08835_ _03672_ _03072_ _04219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08766_ _04170_ _04174_ _04176_ _00783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05978_ rf_ram.memory\[12\]\[0\] _01643_ _01655_ rf_ram.memory\[13\]\[0\] _01653_
+ rf_ram.memory\[15\]\[0\] _02174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XANTENNA_input11_I i_dbus_rdt[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_5_25__f_clk_I clknet_3_6_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07717_ _03488_ _03509_ _03510_ _00400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_36_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09280__C _01391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08697_ rf_ram.memory\[153\]\[1\] _04131_ _04133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_73_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_178_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_95_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07648_ _03455_ _03466_ _03467_ _00374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_32_1108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_81_1910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07579_ _03422_ _03423_ _03424_ _00348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_24_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_24_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09318_ _04527_ _00984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08265__A1 _03823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08691__I _04061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10590_ _00334_ clknet_leaf_165_clk rf_ram.memory\[320\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_63_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_1253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10072__A1 _04985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09249_ _04477_ _04478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_106_635 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05618__A3 _01813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08017__A1 _03686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_79_1861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_79_1872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_151_3192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_142_1107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_133_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06144__C _01717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11211_ _00947_ clknet_leaf_47_clk rf_ram.memory\[82\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08568__A2 _03949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_1264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_118_Left_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_11142_ _00878_ clknet_leaf_35_clk rf_ram.memory\[10\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_112_2475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_112_2486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput76 net76 o_dbus_adr[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__09517__A1 _04643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput87 net87 o_dbus_adr[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_11073_ _00810_ clknet_leaf_54_clk rf_ram.memory\[469\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_179_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput98 net98 o_dbus_dat[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__06160__B _01746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10024_ rf_ram.memory\[246\]\[1\] _04979_ _04981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_99_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06200__B1 _01725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_127_Left_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_158_3324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05504__B _01620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_158_3335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10926_ _00670_ clknet_leaf_8_clk rf_ram.memory\[174\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_168_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10857_ _00601_ clknet_leaf_309_clk rf_ram.memory\[528\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_119_2607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08256__A1 _02845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10788_ _00532_ clknet_leaf_323_clk rf_ram.memory\[562\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_26_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_136_2921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10063__A1 _03445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_59_Right_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_171_3568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_1321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06335__B _01928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08008__A1 _02730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_1039 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_136_Left_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_112_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09756__B2 net118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11409_ _01141_ clknet_leaf_20_clk rf_ram.memory\[77\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_1_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07945__I _03355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07231__A2 _03040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05778__C1 _01925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06950_ _03018_ _03026_ _03028_ _00115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_182_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_input3_I i_dbus_rdt[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_37_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06990__A1 _03053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05465__I _01499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_68_Right_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05901_ rf_ram.memory\[84\]\[0\] _01709_ _01656_ rf_ram.memory\[85\]\[0\] _01763_
+ rf_ram.memory\[87\]\[0\] _02097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_06881_ rf_ram.memory\[301\]\[1\] _02980_ _02982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08620_ _02760_ _02881_ _04085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05832_ rf_ram.memory\[218\]\[0\] _01940_ _01959_ rf_ram.memory\[219\]\[0\] _02027_
+ _02028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__06742__A1 _02881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05545__A2 _01623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_145_Left_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_55_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08551_ rf_ram.memory\[119\]\[1\] _04039_ _04041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05763_ _01695_ _01959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_77_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05950__C1 _01635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07502_ _03360_ _03374_ _03376_ _00319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_89_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08495__A1 _03953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08482_ _03991_ _03993_ _03994_ _00681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05694_ _01887_ _01889_ _01790_ _01890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_49_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_1180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_130_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07433_ _03326_ _03331_ _03333_ _00293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_43_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_76_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_175_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_77_Right_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07364_ _03055_ _02822_ _03290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_73_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09103_ rf_ram.memory\[95\]\[0\] _04384_ _04385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_174_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06315_ rf_ram.memory\[184\]\[1\] _01711_ _01848_ rf_ram.memory\[185\]\[1\] _01773_
+ rf_ram.memory\[187\]\[1\] _02510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XANTENNA__09995__A1 _04953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08798__A2 _04195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07295_ _02984_ _02997_ _03247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_154_Left_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06245__B _01923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09034_ _04334_ _04340_ _04342_ _00885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06246_ rf_ram.memory\[441\]\[1\] _01918_ _02441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_131_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_142_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_96_2183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_170_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09747__A1 net114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09747__B2 net115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06177_ rf_ram.memory\[496\]\[1\] _01644_ _01526_ _02372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_7_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_57_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05128_ cpu.decode.op26 _01331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input59_I i_ibus_rdt[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_57_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_86_Right_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_leaf_280_clk clknet_5_19__leaf_clk clknet_leaf_280_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_74_1780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06430__B1 _01848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09936_ _04918_ _04926_ _04927_ _01203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06981__A1 _03014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05784__A2 _01770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09867_ _02838_ _02921_ _04885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_163_Left_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_70_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08818_ rf_ram.memory\[137\]\[1\] _04207_ _04209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06194__C1 _01696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06733__A1 _02876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09798_ rf_ram.memory\[58\]\[0\] _04842_ _04843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_29_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_29_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08749_ _04126_ _04164_ _04165_ _00777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_5_23__f_clk clknet_3_5_0_clk clknet_5_23__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_95_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_184_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_36_1063 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_1074 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_95_Right_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10711_ _00455_ clknet_leaf_134_clk rf_ram.memory\[40\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_152_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_1310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_181_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10642_ _00386_ clknet_leaf_96_clk rf_ram.memory\[402\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_138_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08238__A1 _03820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_153_3232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_172_Left_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_165_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_153_3243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10045__A1 _04982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09986__A1 _02915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_181_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10573_ _00317_ clknet_leaf_162_clk rf_ram.memory\[364\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_64_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_114_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_1062 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_122_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_958 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_146_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05994__B _01506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08410__A1 _02761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06421__B1 _01772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11125_ _00861_ clknet_leaf_73_clk rf_ram.memory\[118\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_271_clk clknet_5_16__leaf_clk clknet_leaf_271_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_120_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_181_Left_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_11056_ _00793_ clknet_leaf_1_clk rf_ram.memory\[149\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09910__A1 _04887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10007_ rf_ram.memory\[277\]\[0\] _04970_ _04971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_129_2791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05527__A2 _01706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06724__A1 _02820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_99_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_1142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08477__A1 _01491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_1114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_169_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_129_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_173_3608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_1196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10909_ _00653_ clknet_leaf_26_clk rf_ram.memory\[189\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_7_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_184_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_15_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_1248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_15_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_184_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_156_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_144_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09977__A1 _04950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06100_ rf_ram.memory\[272\]\[1\] _01614_ _01615_ _02295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_125_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07080_ rf_ram.memory\[492\]\[1\] _03111_ _03113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_152_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_164_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06031_ rf_ram.memory\[562\]\[1\] _01544_ _01554_ rf_ram.memory\[563\]\[1\] _01555_
+ rf_ram.memory\[561\]\[1\] _02226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_11_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_160_1026 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_39_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_140_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_125_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_188_3884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_188_3895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_262_clk clknet_5_17__leaf_clk clknet_leaf_262_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_10_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_91_2091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07982_ rf_ram.memory\[478\]\[1\] _03673_ _03675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_35_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06933_ _03017_ _03018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_09721_ _04781_ net9 _04792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_52_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09901__A1 _03319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08704__A2 _04078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06864_ _02819_ _02970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_09652_ net1 _04739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_3
XANTENNA__06176__C1 _01519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08603_ net241 _04067_ _04074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_78_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05815_ rf_ram.memory\[180\]\[0\] _01799_ _01772_ rf_ram.memory\[181\]\[0\] _01786_
+ rf_ram.memory\[183\]\[0\] _02011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_171_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09583_ _04695_ _01081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06795_ _02922_ _02923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__05923__C1 _01625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06191__A2 _01856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08534_ rf_ram.memory\[69\]\[1\] _04028_ _04030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05746_ rf_ram.memory\[420\]\[0\] _01666_ _01810_ rf_ram.memory\[421\]\[0\] _01646_
+ rf_ram.memory\[423\]\[0\] _01942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_166_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_148_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_1263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08465_ _01381_ net1 _03982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_77_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05677_ rf_ram.memory\[452\]\[0\] _01666_ _01810_ rf_ram.memory\[453\]\[0\] _01811_
+ rf_ram.memory\[455\]\[0\] _01873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_77_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07140__A1 _03126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07416_ _03292_ _03320_ _03322_ _00287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_161_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_98_2212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08396_ rf_ram.memory\[17\]\[0\] _03933_ _03934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_98_2223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10027__A1 _04911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09968__A1 _04921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07347_ _03260_ _03277_ _03279_ _00261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_33_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_59_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07278_ rf_ram.memory\[417\]\[1\] _03235_ _03237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_60_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_76_1820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09017_ _04057_ _04331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_06229_ rf_ram.memory\[410\]\[1\] _01801_ _01726_ rf_ram.memory\[411\]\[1\] _01721_
+ rf_ram.memory\[409\]\[1\] _02424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_130_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09440__I0 net70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_991 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_72_1739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_253_clk clknet_5_20__leaf_clk clknet_leaf_253_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__06403__B1 _01656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09919_ _04884_ _04915_ _04916_ _01197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06706__A1 _02826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06182__A2 _01846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_107_2385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_945 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_185_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08459__A1 net120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_185_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07131__A1 _02806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_458 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_166_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_153_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10018__A1 _04950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09959__A1 _04911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_12_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10186__I _02747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10625_ _00369_ clknet_leaf_95_clk rf_ram.memory\[388\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_153_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_1210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_148_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07434__A2 _02815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10556_ _00300_ clknet_leaf_148_clk rf_ram.memory\[368\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_49_1254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10487_ _00231_ clknet_leaf_42_clk rf_ram.memory\[196\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05996__A2 _01524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07198__A1 _03161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_184_Right_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_20_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_244_clk clknet_5_21__leaf_clk clknet_leaf_244_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08934__A2 _03559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_166_3478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05748__A2 _01662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06945__A1 _03018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11108_ _00844_ clknet_leaf_85_clk rf_ram.memory\[124\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_183_3792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11039_ _00776_ clknet_leaf_275_clk rf_ram.i_raddr\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_4
XANTENNA__08698__A1 _04129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07370__A1 _02781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_1258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06173__A2 _01652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05600_ _01775_ _01781_ _01791_ _01795_ _01796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_177_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_148_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06580_ _02734_ _02762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__05381__B1 _01539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_19_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05531_ rf_ram.memory\[328\]\[0\] _01724_ _01725_ rf_ram.memory\[329\]\[0\] _01726_
+ rf_ram.memory\[331\]\[0\] _01727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_59_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05899__B _01746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_157_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08250_ _03823_ _03840_ _03842_ _00601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_117_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_89_1034 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05462_ _01563_ _01658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_129_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07201_ _03157_ _03187_ _03188_ _00206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_55_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08181_ _03787_ _03799_ _03800_ _00574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_55_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05393_ rf_ram.memory\[568\]\[0\] _01524_ _01528_ _01589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_15_525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_31_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_144_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_31_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07132_ rf_ram.memory\[486\]\[0\] _03145_ _03146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_43_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08622__A1 _04058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_93_2120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_1207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_93_2131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07063_ rf_ram.memory\[375\]\[0\] _03102_ _03103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_113_744 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput200 net200 o_ext_rs2[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput211 net211 o_ibus_adr[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_06014_ _02205_ _02206_ _02207_ _02208_ _01564_ _02209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
Xoutput222 net222 o_ibus_adr[28] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_11_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput233 net233 o_ibus_adr[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__09178__A2 _04418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_1040 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_54_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07189__A1 _02836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_151_Right_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_leaf_235_clk clknet_5_22__leaf_clk clknet_leaf_235_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_26_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06397__C1 _01773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05739__A2 _01804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06936__A1 _02766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07965_ rf_ram.memory\[470\]\[1\] _03662_ _03664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11655__I net105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_1296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09704_ net100 _04767_ _04768_ net101 _04779_ _04780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__06749__I _02888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06916_ _02970_ _03004_ _03005_ _00104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07896_ _03619_ _03620_ _03621_ _00468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09350__A2 _03991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09635_ _04524_ net60 _04726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_69_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06847_ _02750_ _02837_ _02959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_179_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_139_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_1072 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09566_ cpu.immdec.imm30_25\[1\] _04682_ _04678_ _04683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08964__I _04057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06778_ _02764_ _02830_ _02910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_69_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05911__A2 _01787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10248__A1 _02825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09102__A2 _04005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08517_ rf_ram.memory\[172\]\[1\] _04017_ _04019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05729_ _01695_ _01925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_09497_ _04628_ _04629_ _04630_ _04631_ _01440_ _04632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XANTENNA__07113__A1 _03126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08861__A1 _02983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08448_ _03956_ _03964_ _03966_ _00675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_102_2293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_1320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_184_1313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_136_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_981 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08379_ _03922_ _03920_ _03923_ _00649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_151_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10410_ _00154_ clknet_leaf_111_clk rf_ram.memory\[375\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_18_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11390_ _01122_ clknet_leaf_228_clk net104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_116_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10341_ _00085_ clknet_leaf_173_clk rf_ram.memory\[284\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_60_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_182_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_1032 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05978__A2 _01643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10272_ _00016_ clknet_leaf_261_clk rf_ram.memory\[234\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_103_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_226_clk clknet_5_23__leaf_clk clknet_leaf_226_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_148_3142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_148_3153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05991__C _01373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_109_2414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_109_2425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_161_3386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07352__A1 _03260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06155__A2 _01677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_17_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_186_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_158_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05363__B1 _01555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_17_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_122_2658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_100_Left_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05902__A2 _01863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_122_2669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10239__A1 _02737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07104__A1 _02915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_1069 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_948 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05512__B _01707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_1177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08852__A1 _04202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_1229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11657_ net107 net179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_36_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_154_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10608_ _00352_ clknet_leaf_156_clk rf_ram.memory\[355\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_36_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_181_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11588_ _01320_ clknet_leaf_32_clk rf_ram.memory\[208\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_101_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_168_3507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10539_ _00283_ clknet_leaf_213_clk rf_ram.memory\[247\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_122_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_168_3518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06343__B _01916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05969__A2 _01682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_185_3821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_150_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_185_3832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_217_clk clknet_5_22__leaf_clk clknet_leaf_217_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08907__A2 _04038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06918__A1 _02975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_1314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07750_ rf_ram.memory\[377\]\[1\] _03529_ _03531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_56_1000 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06701_ _02826_ _02853_ _02855_ _00039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07681_ _03458_ _03485_ _03487_ _00387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06146__A2 _01724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07343__A1 _03055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06632_ _02743_ _02802_ _02803_ _00022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09420_ _04585_ _01028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_17_1028 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07894__A2 _02844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_1099 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06563_ _02747_ _02748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_09351_ _04546_ _00998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_59_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09096__A1 _04367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_47_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05514_ rf_ram.memory\[324\]\[0\] _01709_ _01656_ rf_ram.memory\[325\]\[0\] _01654_
+ rf_ram.memory\[327\]\[0\] _01710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_08302_ _03855_ _03872_ _03874_ _00621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09282_ _04497_ _04502_ _04503_ _00972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_47_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_173_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07646__A2 _03089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06494_ _01371_ _02688_ _02689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_63_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_173_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06237__C net254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08233_ _03820_ _03831_ _03832_ _00594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_51_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_970 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05445_ _01640_ _01641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__05141__C cpu.genblk3.csr.o_new_irq vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_173_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08164_ _03787_ _03788_ _03789_ _00568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05376_ rf_ram.memory\[556\]\[0\] _01511_ _01517_ rf_ram.memory\[557\]\[0\] _01521_
+ rf_ram.memory\[559\]\[0\] _01572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_126_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_1102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_166_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07115_ _03134_ _03135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_30_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_995 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08095_ _03721_ _03745_ _03746_ _00542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06253__B _01805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06082__A1 _01603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_140_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07046_ _03087_ _03090_ _03091_ _00148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_140_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_208_clk clknet_5_19__leaf_clk clknet_leaf_208_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09020__A1 _04331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06909__A1 _02822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input41_I i_ibus_rdt[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08997_ _02945_ _04303_ _04319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06385__A2 _01918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07582__A1 _03425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05593__B1 _01786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07948_ _03651_ _03652_ _03653_ _00488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_143_3050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09323__A2 _04037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06137__A2 _01777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07879_ rf_ram.memory\[446\]\[0\] _03610_ _03611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_output128_I net128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_1106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_104_2322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09618_ _04643_ _01460_ _04707_ _01092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_67_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_104_2333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05345__B1 _01539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_67_1649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10890_ _00634_ clknet_leaf_214_clk rf_ram.memory\[240\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_70_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_1139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05896__A1 _01769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_84_1952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09087__A1 _02983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09549_ _01447_ _01339_ _04669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_84_1963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_155_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08834__A1 _04205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_175_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11511_ _01243_ clknet_leaf_150_clk rf_ram.memory\[305\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_53_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_163_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11442_ _01174_ clknet_leaf_239_clk cpu.state.genblk1.misalign_trap_sync_r vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__05986__C _01493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11373_ _01105_ clknet_leaf_60_clk rf_ram.memory\[78\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_150_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08062__A2 _03693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10324_ _00068_ clknet_leaf_135_clk rf_ram.memory\[291\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_131_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05820__A1 _01768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10255_ rf_ram.memory\[9\]\[0\] _05122_ _05123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09011__A1 _04301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_163_3415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_1000 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_163_3426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10186_ _02747_ _05081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__07573__A1 _03389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06376__A2 _01863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_180_3740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05584__B1 _01778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1088 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_124_2709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09314__A2 net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07325__A1 _03257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06128__A2 _01692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_178_3691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_155_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07628__A2 _03452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08825__A1 _02828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05639__A1 _01527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_139_2974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06300__A2 _01846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_139_2985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_127_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05230_ _01429_ _01430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_127_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_154_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_42_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_181_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_42_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_108_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_25_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05161_ cpu.state.genblk1.misalign_trap_sync_r _01364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__09250__A1 _04478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05468__I _01514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08920_ rf_ram.memory\[389\]\[0\] _04271_ _04272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09002__A1 _02953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_1032 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_62_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08851_ rf_ram.memory\[132\]\[0\] _04228_ _04229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07802_ rf_ram.memory\[435\]\[0\] _03563_ _03564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_88_2030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05994_ rf_ram.memory\[526\]\[1\] _01502_ _01506_ _02189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08782_ net243 _04152_ _04186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_88_2041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07733_ rf_ram.memory\[397\]\[1\] _03518_ _03520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_5_4__f_clk clknet_3_1_0_clk clknet_5_4__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_0_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06119__A2 _01509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_49_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07664_ rf_ram.memory\[385\]\[1\] _03475_ _03477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_324_clk_I clknet_5_5__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_79_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_172_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09403_ _04574_ _01022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__05878__A1 _01368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06615_ _02766_ _02788_ _02789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_94_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07595_ _03422_ _03433_ _03434_ _00354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09069__A1 _04334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_149_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_1150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06248__B _01928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06546_ rf_ram_if.rtrig1 rf_ram_if.wen0_r rf_ram_if.wen1_r _01347_ _02732_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_09334_ rf_ram.memory\[99\]\[0\] _04536_ _04537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07619__A2 _03390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_1003 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_339_clk_I clknet_5_0__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_146_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09265_ cpu.genblk3.csr.mstatus_mpie _04481_ _04491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06477_ _01903_ _02670_ _02671_ _02672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_173_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_161_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_69_1246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08216_ rf_ram.memory\[534\]\[0\] _03821_ _03822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_16_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05428_ _01518_ _01624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_173_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09196_ _04431_ _04442_ _04443_ _00946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_105_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05359_ _01516_ _01555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_08147_ rf_ram.memory\[547\]\[0\] _03778_ _03779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09241__A1 _01418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08078_ _02945_ _03729_ _03736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_30_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07029_ _02738_ _02992_ _03079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_101_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_8_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10040_ _04982_ _04990_ _04991_ _01243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_105_1188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09544__A2 net42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06358__A2 _01940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07555__A1 _03393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_141_3009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_168_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10942_ _00680_ clknet_leaf_280_clk rf_ram_if.rdata1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_98_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07858__A2 _02869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09313__I _03992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10873_ _00617_ clknet_leaf_46_clk rf_ram.memory\[192\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_27_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_149_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08807__A1 _04170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_186_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_54_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_1313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_156_3285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08283__A2 _02788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_156_3296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10090__A2 _03009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_117_2568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11425_ _01157_ clknet_leaf_201_clk rf_ram.memory\[259\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_117_2579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09232__A1 _04463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_989 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08035__A2 _03693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_954 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_134_2882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_134_2893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_22_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11356_ _01088_ clknet_leaf_20_clk rf_ram.memory\[73\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_104_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07794__A1 _03557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10307_ _00051_ clknet_leaf_273_clk rf_ram.memory\[517\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11287_ _01022_ clknet_leaf_243_clk net223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10238_ _02825_ _05110_ _05112_ _01320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06349__A2 _01801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07546__A1 _02921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10169_ _05046_ _05069_ _05070_ _01293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05557__B1 _01645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_1101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_1172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_88_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_1074 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_159_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_1204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06400_ rf_ram.memory\[90\]\[1\] _01801_ _01646_ rf_ram.memory\[91\]\[1\] _01810_
+ rf_ram.memory\[89\]\[1\] _02595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_07380_ _02775_ _03253_ _03300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_44_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06331_ _02523_ _02525_ _01978_ _02526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_128_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06285__A1 _01972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09050_ _02805_ _04339_ _04352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_06262_ _02453_ _02454_ _02455_ _02456_ _01717_ _02457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_154_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_115_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_170_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05213_ cpu.state.cnt_r\[3\] cpu.mem_bytecnt\[1\] _01385_ cpu.state.o_cnt\[2\] _01413_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_08001_ _02761_ _02832_ _03687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_128_1133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09223__A1 _04434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06193_ rf_ram.memory\[478\]\[1\] _01543_ _02388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_142_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_1252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05144_ rf_ram_if.rtrig0 _01347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_64_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07785__A1 _03521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_1127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_141_1322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09952_ rf_ram.memory\[337\]\[1\] _04935_ _04937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_60_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08903_ rf_ram.memory\[126\]\[0\] _04260_ _04261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05260__A2 _01437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09883_ _04884_ _04893_ _04894_ _01183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08834_ _04205_ _04216_ _04218_ _00809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_32_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_139_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_leaf_263_clk_I clknet_5_17__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08765_ rf_ram.memory\[145\]\[1\] _04174_ _04176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05977_ rf_ram.memory\[14\]\[0\] _01640_ _01503_ _02173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_100_1096 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11663__I net114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07716_ rf_ram.memory\[380\]\[0\] _03509_ _03510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_68_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_170_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08696_ _04126_ _04131_ _04132_ _00757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05661__I _01695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_1114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_1136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07647_ rf_ram.memory\[405\]\[0\] _03466_ _03467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_177_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_81_1900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06512__A2 cpu.decode.opcode\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_81_1911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_1289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11368__CLK clknet_5_20__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_278_clk_I clknet_5_17__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07578_ rf_ram.memory\[356\]\[0\] _03423_ _03424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_24_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_24_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09317_ _04526_ net64 _04521_ cpu.immdec.imm11_7\[3\] _04522_ cpu.immdec.imm11_7\[2\]
+ _04527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_06529_ _02714_ _02715_ net234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_36_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05610__B _01805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_69_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_173_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09248_ net34 _04477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_0_63_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output195_I net195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_201_clk_I clknet_5_25__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05484__C1 _01679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_161_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09214__A1 net240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09179_ rf_ram.memory\[84\]\[0\] _04432_ _04433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_79_1862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_151_3193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_79_1873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11210_ _00946_ clknet_leaf_47_clk rf_ram.memory\[82\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_32_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09765__A2 _04766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07776__A1 _03524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_max_cap241_I _02882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11141_ _00877_ clknet_leaf_69_clk rf_ram.memory\[110\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_216_clk_I clknet_5_22__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_112_2476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output72_I net72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_112_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput77 net77 o_dbus_adr[20] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_11072_ _00809_ clknet_leaf_52_clk rf_ram.memory\[459\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xoutput88 net88 o_dbus_adr[30] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput99 net99 o_dbus_dat[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_10023_ _04950_ _04979_ _04980_ _01237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_76_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_169_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10925_ _00669_ clknet_leaf_296_clk rf_ram.memory\[59\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_85_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_158_3325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_158_3336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07700__A1 _02945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06503__A2 cpu.genblk3.csr.o_new_irq vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_1070 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_168_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10856_ _00600_ clknet_leaf_309_clk rf_ram.memory\[528\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_6_1165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_175_3650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_184_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_119_2608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08256__A2 _02972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10787_ _00531_ clknet_leaf_332_clk rf_ram.memory\[563\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_125_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_137_783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_136_2922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06267__A1 _01373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10063__A2 _02866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_1143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_171_3569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_152_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09756__A2 _04766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11408_ _01140_ clknet_5_28__leaf_clk rf_ram.memory\[269\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_10_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07767__A1 _02752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11339_ _01071_ clknet_leaf_215_clk cpu.immdec.imm19_12_20\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05778__B1 _01912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06351__B _01350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_37_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05900_ rf_ram.memory\[86\]\[0\] _01785_ _01707_ _02096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_06880_ _02970_ _02980_ _02981_ _00092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_94_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_1114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_175_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_59_1245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_1079 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05831_ rf_ram.memory\[217\]\[0\] _01515_ _02027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_179_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06742__A2 _02883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05762_ _01640_ _01958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_08550_ _04023_ _04039_ _04040_ _00703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_89_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05950__B1 _01609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05481__I _01633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07501_ rf_ram.memory\[324\]\[1\] _03374_ _03376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05693_ rf_ram.memory\[386\]\[0\] _01856_ _01786_ rf_ram.memory\[387\]\[0\] _01888_
+ _01889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_08481_ cpu.state.ibus_cyc _03993_ _03994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_159_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_840 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09692__B2 net128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07432_ rf_ram.memory\[370\]\[1\] _03331_ _03333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_186_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_174_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_147_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07363_ _03013_ _03289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_72_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09102_ _02908_ _04005_ _04384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06314_ rf_ram.memory\[186\]\[1\] _01989_ _01916_ _02509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07294_ _03225_ _03244_ _03246_ _00241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_66_1205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_115_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_127_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_26_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09033_ rf_ram.memory\[106\]\[1\] _04340_ _04342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06245_ rf_ram.memory\[440\]\[1\] _01922_ _01923_ _02440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_142_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_96_2173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_96_2184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06176_ rf_ram.memory\[500\]\[1\] _01509_ _01668_ rf_ram.memory\[501\]\[1\] _01519_
+ rf_ram.memory\[503\]\[1\] _02371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_13_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_1093 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_57_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_159_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05769__B1 _01953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_57_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_74_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09935_ rf_ram.memory\[340\]\[0\] _04926_ _04927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_141_1174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_74_1781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_1125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_1147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_1282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09866_ _04396_ _04884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__08183__A1 _03790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08817_ _04202_ _04207_ _04208_ _00802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06194__B1 _01848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09797_ net245 _02921_ _04842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07930__A1 _02991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_82_clk_I clknet_5_11__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08748_ rf_ram.memory\[147\]\[0\] _04164_ _04165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_96_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_913 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_36_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08679_ _04094_ _04120_ _04121_ _00751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09683__A1 net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10710_ _00454_ clknet_leaf_134_clk rf_ram.memory\[40\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_67_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_97_clk_I clknet_5_14__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_187_1322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10641_ _00385_ clknet_leaf_92_clk rf_ram.memory\[384\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_48_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_140_clk_I clknet_5_27__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_153_3233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_153_3244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10572_ _00316_ clknet_leaf_162_clk rf_ram.memory\[364\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09986__A2 _03083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_945 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_165_Right_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_134_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_20_clk_I clknet_5_3__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_114_2516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_131_2830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_155_clk_I clknet_5_26__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_913 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07749__A1 _03521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08410__A2 _03903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_35_clk_I clknet_5_6__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11124_ _00860_ clknet_leaf_76_clk rf_ram.memory\[118\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_43_1079 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11055_ _00792_ clknet_leaf_1_clk rf_ram.memory\[149\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10006_ _02940_ _03072_ _04970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_129_2792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_1121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_157_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_118_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_1078 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08477__A2 _03989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_156_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10908_ _00652_ clknet_leaf_13_clk rf_ram.memory\[189\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_173_3609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_670 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05696__C1 _01848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_184_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_108_clk_I clknet_5_15__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10839_ _00583_ clknet_leaf_314_clk rf_ram.memory\[537\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_156_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_15_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06346__B _01805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_171_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09977__A2 _04951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_132_Right_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07988__A1 _03654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06030_ rf_ram.memory\[560\]\[1\] _01511_ _01552_ _02225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_124_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_948 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_39_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_39_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_188_3885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_188_3896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_1146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_91_2081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_91_2092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07981_ _03651_ _03673_ _03674_ _00500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09720_ _04760_ _04791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_06932_ _02747_ _03017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_52_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09901__A2 _02984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09651_ net98 _04737_ _04738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06863_ _02930_ _02967_ _02969_ _00087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06176__B1 _01668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07912__A1 _03619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08602_ _04062_ _04071_ _04073_ _00722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05425__B _01620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05814_ rf_ram.memory\[182\]\[0\] _01631_ _01505_ _02010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09582_ cpu.immdec.imm30_25\[5\] _04678_ _04694_ _04695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06794_ _02773_ _02759_ _02922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_78_913 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05923__B1 _01702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_1231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_89_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08533_ _04023_ _04028_ _04029_ _00697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05745_ rf_ram.memory\[422\]\[0\] _01940_ _01805_ _01941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_49_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08464_ _01442_ _01447_ _03980_ _01399_ _03981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_05676_ rf_ram.memory\[454\]\[0\] _01804_ _01805_ _01872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_175_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07415_ rf_ram.memory\[334\]\[1\] _03320_ _03322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_147_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08395_ _02761_ _02997_ _03933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_98_2213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_98_2224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_169_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_162_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10027__A2 _02829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07346_ rf_ram.memory\[253\]\[1\] _03277_ _03279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_116_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07979__A1 _03672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_61_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07277_ _03222_ _03235_ _03236_ _00234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_115_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_33_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_115_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_76_1810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09016_ _04301_ _04328_ _04330_ _00879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06228_ rf_ram.memory\[408\]\[1\] _01755_ _01615_ _02423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06770__I _02903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_76_1821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06159_ rf_ram.memory\[490\]\[1\] _01687_ _01688_ rf_ram.memory\[491\]\[1\] _02353_
+ _02354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__09440__I1 net71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_1729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output158_I net158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05611__C1 _01726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09918_ rf_ram.memory\[343\]\[0\] _04915_ _04916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08156__A1 net238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09849_ _02713_ _04873_ _01169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_137_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_154_1321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_1137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_87_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_1039 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_107_2386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_150_1218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_139_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_178_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07131__A2 _02911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_7_1293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_12_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10624_ _00368_ clknet_leaf_94_clk rf_ram.memory\[388\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09959__A2 _02954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05693__A2 _01856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06890__A1 _02788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_12_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_153_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_1200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_1136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_107_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_1109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10555_ _00299_ clknet_leaf_151_clk rf_ram.memory\[331\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_134_561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09477__B _03989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_24_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06642__A1 _02756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_1168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10486_ _00230_ clknet_leaf_43_clk rf_ram.memory\[196\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_32_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_121_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09431__I1 net67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08395__A1 _02761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_166_3468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_166_3479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05602__C1 _01713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11107_ _00843_ clknet_leaf_116_clk rf_ram.memory\[389\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_120_1055 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_183_3793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11038_ _00775_ clknet_leaf_285_clk rf_ram.i_raddr\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__09895__A1 _04887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07370__A2 _03253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05530_ _01635_ _01726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_75_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05461_ rf_ram.memory\[378\]\[0\] _01652_ _01654_ rf_ram.memory\[379\]\[0\] _01656_
+ rf_ram.memory\[377\]\[0\] _01657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_138_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_leaf_180_clk clknet_5_31__leaf_clk clknet_leaf_180_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__06330__B1 _02019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06076__B _01684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_144_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07200_ rf_ram.memory\[273\]\[0\] _03187_ _03188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05684__A2 _01770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08180_ rf_ram.memory\[541\]\[0\] _03799_ _03800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05392_ rf_ram.memory\[572\]\[0\] _01538_ _01555_ rf_ram.memory\[573\]\[0\] _01554_
+ rf_ram.memory\[575\]\[0\] _01588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_89_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_43_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_31_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07131_ _02806_ _02911_ _03145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_15_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07686__I _03359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_93_2121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05436__A2 _01631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07062_ _03082_ _03101_ _03102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_93_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput201 net201 o_ext_rs2[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_06013_ rf_ram.memory\[538\]\[1\] _01544_ _01540_ rf_ram.memory\[539\]\[1\] _01539_
+ rf_ram.memory\[537\]\[1\] _02208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
Xoutput212 net212 o_ibus_adr[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput223 net223 o_ibus_adr[29] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput234 net234 o_ibus_cyc vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_140_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_54_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_140_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07189__A2 _02984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10193__A1 _05081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06397__B1 _01772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06936__A2 _02883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_1310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_1253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07964_ _03651_ _03662_ _03663_ _00494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08138__A1 _03754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09703_ _04740_ net4 _04779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_06915_ rf_ram.memory\[298\]\[0\] _03004_ _03005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07895_ rf_ram.memory\[461\]\[0\] _03620_ _03621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09886__A1 _03892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09634_ _04524_ _01380_ _04725_ _01102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06846_ _02940_ _02958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_09565_ _03992_ _04680_ _04681_ _04682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05372__A1 _01347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06777_ _02908_ _02909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__09638__A1 _04524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_69_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11671__I cpu.ctrl.pc vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_69_1691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_167_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08516_ _03953_ _04017_ _04018_ _00691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_93_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05728_ rf_ram.memory\[440\]\[0\] _01922_ _01923_ _01924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_33_1023 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09496_ cpu.alu.cmp_r _01388_ _04630_ _04631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_77_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08310__A1 _03852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08447_ rf_ram.memory\[176\]\[1\] _03964_ _03966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_171_clk clknet_5_30__leaf_clk clknet_leaf_171_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_93_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_102_2294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05659_ rf_ram.memory\[472\]\[0\] _01782_ _01783_ _01855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_175_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08861__A2 _03559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06872__A1 _02975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08378_ rf_ram.memory\[186\]\[1\] _03920_ _03923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_135_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_12_Left_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_61_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07329_ rf_ram.memory\[271\]\[0\] _03268_ _03269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_162_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_150_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06085__C1 _01654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06624__A1 cpu.immdec.imm11_7\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10340_ _00084_ clknet_leaf_173_clk rf_ram.memory\[284\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_116_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06433__C _01978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10271_ _00015_ clknet_leaf_277_clk rf_ram.memory\[233\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_44_1141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_148_3143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_21_Left_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_109_2415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09316__I _03992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_109_2426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_126_2740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_161_3376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_161_3387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_159_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_1322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_154_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_17_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09629__A1 _04524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_1135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_122_2659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_1270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_1150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10239__A2 _03071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_1168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07104__A2 _03072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_162_clk clknet_5_30__leaf_clk clknet_leaf_162_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_167_995 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_166_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06863__A1 _02930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05666__A2 _01543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11656_ net106 net178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_181_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10607_ _00351_ clknet_leaf_154_clk rf_ram.memory\[316\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_153_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_153_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11587_ _01319_ clknet_leaf_300_clk rf_ram.memory\[208\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09801__A1 _04840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06615__A1 _02766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10538_ _00282_ clknet_leaf_208_clk rf_ram.memory\[247\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_101_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_168_3508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_168_3519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_161_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06091__A2 _01706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_185_3822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10469_ _00213_ clknet_leaf_195_clk rf_ram.memory\[260\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_185_3833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_946 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08368__A1 _02983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_1214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09654__C _04740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07040__A1 _03053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09317__C2 cpu.immdec.imm11_7\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06700_ rf_ram.memory\[523\]\[1\] _02853_ _02855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07680_ rf_ram.memory\[402\]\[1\] _03485_ _03487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08540__A1 _04026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07343__A2 _02960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06000__C1 _01540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06631_ rf_ram.memory\[293\]\[0\] _02802_ _02803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_149_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09350_ net229 _03991_ _04540_ net230 _04546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_48_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_177_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06562_ _02746_ _02747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_176_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_59_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08301_ rf_ram.memory\[244\]\[1\] _03872_ _03874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_47_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05513_ _01508_ _01709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_09281_ cpu.genblk3.csr.mcause3_0\[2\] _04497_ _04503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_47_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_153_clk clknet_5_26__leaf_clk clknet_leaf_153_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_142_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06493_ _02519_ _02575_ _02687_ _01373_ _02688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_117_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06854__A1 _02839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08232_ rf_ram.memory\[531\]\[0\] _03831_ _03832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05657__A2 _01785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05444_ _01499_ _01640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_142_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_173_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_172_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_1022 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08163_ rf_ram.memory\[544\]\[0\] _03788_ _03789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_43_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05375_ rf_ram.memory\[558\]\[0\] _01502_ _01506_ _01571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_172_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06534__B _01347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07114_ _02716_ _03007_ _03134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__06606__A1 _02766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08094_ rf_ram.memory\[557\]\[0\] _03745_ _03746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_42_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_1185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_1027 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07045_ rf_ram.memory\[391\]\[0\] _03090_ _03091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_63_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_11_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_5_19__f_clk_I clknet_3_4_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10166__A1 _05049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06909__A2 _02997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07031__A1 _03050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08996_ _04301_ _04316_ _04318_ _00871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05664__I _01563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input34_I i_ibus_ack vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07947_ rf_ram.memory\[456\]\[0\] _03652_ _03653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_143_3051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07878_ _02916_ _03234_ _03610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_3_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08531__A1 _02794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09617_ _04637_ _04717_ _04719_ _01091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06829_ _02935_ _02946_ _02947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_67_1639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_104_2323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_104_2334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_168_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05613__B _01650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09548_ _04667_ _04654_ _04668_ _01073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_66_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_84_1953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_84_1964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09087__A2 _03765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07098__A1 _02921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06428__C _01860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_144_clk clknet_5_27__leaf_clk clknet_leaf_144_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09479_ cpu.bufreg.i_sh_signed net89 _03989_ _04617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_164_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11510_ _01242_ clknet_leaf_143_clk rf_ram.memory\[326\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_108_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06845__A1 _02930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_163_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_993 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_136_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_1065 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11441_ _01173_ clknet_leaf_233_clk cpu.mem_if.signbit vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_80_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_151_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08598__A1 _02794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11372_ _01104_ clknet_leaf_235_clk cpu.branch_op vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_33_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05805__C1 _01953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06073__A2 _01626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10323_ _00067_ clknet_leaf_288_clk rf_ram.memory\[50\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_81_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10254_ net249 _03035_ _05122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10157__A1 _02787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_163_3416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_163_3427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10185_ _05078_ _05079_ _05080_ _01299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05574__I _01530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_180_3730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_180_3741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05887__A2 _01918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_186_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_1196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_178_3692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07089__A1 _03087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_173_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_135_clk clknet_5_24__leaf_clk clknet_leaf_135_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_16_1073 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08825__A2 _04195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06836__A1 _02927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_166_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_139_2975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_139_2986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_126_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11639_ net98 net170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_71_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_108_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_42_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08589__A1 _04058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05160_ _01334_ _01337_ _01363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__08125__I _03692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09250__A2 cpu.bufreg.i_sh_signed vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06064__A2 _01666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05811__A2 _01641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09002__A2 _04303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08850_ net241 _04195_ _04228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_100_1201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07801_ _02866_ _03234_ _03563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_08781_ _04170_ _04183_ _04185_ _00789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_88_2031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_174_1313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05993_ _01371_ _01594_ _01950_ _02188_ _00000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_TAPCELL_ROW_88_2042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07732_ _03488_ _03518_ _03519_ _00406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_0_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09561__I0 cpu.immdec.imm30_25\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_49_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07663_ _03455_ _03475_ _03476_ _00380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_79_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09402_ net223 _03990_ _04564_ net225 _04574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_149_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06614_ _02787_ _02788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__05878__A2 _02046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07594_ rf_ram.memory\[315\]\[0\] _03433_ _03434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_62_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07204__I _03013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09333_ net240 _04037_ _04536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_146_910 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06545_ cpu.immdec.imm11_7\[3\] _02729_ _02730_ _02731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
Xclkbuf_leaf_126_clk clknet_5_13__leaf_clk clknet_leaf_126_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_47_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_62_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06827__A1 _02716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_62_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09264_ _04486_ _04489_ _04490_ _02713_ _00967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_30_1037 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06476_ rf_ram.memory\[28\]\[1\] _01633_ _01609_ rf_ram.memory\[29\]\[1\] _01607_
+ rf_ram.memory\[31\]\[1\] _02671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_0_28_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_173_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08215_ _03798_ _03009_ _03821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_117_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05427_ _01605_ _01623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_09195_ rf_ram.memory\[82\]\[0\] _04442_ _04443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_161_946 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06264__B _02458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08146_ _02888_ _03765_ _03778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_05358_ _01520_ _01554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_30_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09241__A2 _03989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08077_ _03724_ _03733_ _03735_ _00535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_144_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05289_ _01431_ _01486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_140_1003 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_1172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_12_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05802__A2 _01989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07028_ _03053_ _03076_ _03078_ _00143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06460__C1 _01655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10139__A1 _05046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_1171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_8_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07004__A1 _03050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_1144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08979_ _04298_ _04307_ _04308_ _00864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08504__A1 _03956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10941_ _00679_ clknet_leaf_280_clk rf_ram_if.rdata0\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_168_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06439__B _01601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05869__A2 _01606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10872_ _00616_ clknet_leaf_46_clk rf_ram.memory\[192\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_38_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_1176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_155_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_117_clk clknet_5_14__leaf_clk clknet_leaf_117_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_27_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_1284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06818__A1 _02930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_156_3286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_156_3297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06174__B _01629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_911 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09768__B1 _04760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11424_ _01156_ clknet_leaf_293_clk rf_ram.memory\[7\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_124_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_149_1094 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_117_2569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_151_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07243__A1 _03190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06046__A2 _01606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_134_2883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11355_ _01087_ clknet_leaf_259_clk cpu.decode.op26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_134_2894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08991__A1 _04301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10306_ _00050_ clknet_leaf_270_clk rf_ram.memory\[517\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11286_ _01021_ clknet_leaf_242_clk net222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_123_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10237_ rf_ram.memory\[208\]\[1\] _05110_ _05112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_120_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_5_Left_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07546__A2 _02889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06203__C1 _01811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10168_ rf_ram.memory\[447\]\[0\] _05069_ _05070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_156_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10099_ _05017_ _05025_ _05027_ _01266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_107_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_159_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_107_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05253__B cpu.mem_bytecnt\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_179_Right_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_18_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_159_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06068__C net253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09440__S _04593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_130_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_29_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_108_clk clknet_5_15__leaf_clk clknet_leaf_108_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_44_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06330_ rf_ram.memory\[210\]\[1\] _01804_ _02019_ rf_ram.memory\[211\]\[1\] _02524_
+ _02525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_123_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_84_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07482__A1 _03360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06261_ rf_ram.memory\[418\]\[1\] _01801_ _01646_ rf_ram.memory\[419\]\[1\] _01645_
+ rf_ram.memory\[417\]\[1\] _02456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_143_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06084__B _01707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_128_1112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08000_ _03685_ _03686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__05479__I _01602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_985 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05212_ _01375_ _01411_ _01412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__09759__B1 _04760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06192_ _02384_ _02386_ _01860_ _02387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_25_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05143_ _01332_ _01338_ _01341_ _01345_ _01346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_124_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_151_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_1106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07694__I _03100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08982__A1 net242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09951_ _04918_ _04935_ _04936_ _01209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_40_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08902_ _02916_ _04038_ _04260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_5_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09882_ rf_ram.memory\[229\]\[0\] _04893_ _04894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08734__A1 _04129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08833_ rf_ram.memory\[459\]\[1\] _04216_ _04218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08764_ _04167_ _04174_ _04175_ _00782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05976_ _02160_ _02164_ _02168_ _02171_ _02172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_25_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07715_ _02839_ _03496_ _03509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_135_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_170_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_1202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08695_ rf_ram.memory\[153\]\[0\] _04131_ _04132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_75_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07646_ _03071_ _03089_ _03466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_71_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_146_Right_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_81_1901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_841 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_81_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07577_ _02882_ _03390_ _03423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_76_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_24_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_24_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09316_ _03992_ _04526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_06528_ cpu.state.ibus_cyc _02715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_119_954 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_987 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07473__A1 _03356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09247_ _03967_ net56 _04476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06276__A2 _01664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06459_ rf_ram.memory\[48\]\[1\] _01643_ _01525_ _02654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_90_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05484__B1 _01678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_1288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_1200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09178_ _03134_ _04418_ _04432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_185_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_160_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output188_I net188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09214__A2 _04418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_79_1863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_160_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_79_1874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07225__A1 _03193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_151_3194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06028__A2 _01532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08129_ rf_ram.memory\[551\]\[1\] _03766_ _03768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11140_ _00876_ clknet_leaf_69_clk rf_ram.memory\[110\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_31_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_112_2477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput67 net67 o_dbus_adr[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput78 net78 o_dbus_adr[21] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_11071_ _00808_ clknet_leaf_52_clk rf_ram.memory\[459\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_179_1032 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput89 net89 o_dbus_adr[31] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_10022_ rf_ram.memory\[246\]\[0\] _04979_ _04980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_99_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06200__A2 _01724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_338_clk clknet_5_0__leaf_clk clknet_leaf_338_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_98_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09150__A1 _04401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10924_ _00668_ clknet_leaf_296_clk rf_ram.memory\[59\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_85_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_158_3326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_158_3337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_113_Right_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_85_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10855_ _00599_ clknet_leaf_297_clk rf_ram.memory\[52\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_116_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_175_3640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_175_3651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_119_2609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10786_ _00530_ clknet_leaf_329_clk rf_ram.memory\[563\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_9_clk_I clknet_5_0__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_136_2923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07464__A1 _02921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05299__I _01494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06019__A2 _01524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07216__A1 _02883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11407_ _01139_ clknet_leaf_191_clk rf_ram.memory\[269\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_10_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_323_clk_I clknet_5_4__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11338_ _01070_ clknet_leaf_216_clk cpu.csr_imm vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_123_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06351__C _02545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11269_ _01004_ clknet_leaf_246_clk net204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08716__A1 _04126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_37_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_338_clk_I clknet_5_0__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05830_ rf_ram.memory\[216\]\[0\] _01537_ _01551_ _02026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_59_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05762__I _01640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_89_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05761_ rf_ram.memory\[152\]\[0\] _01735_ _01956_ _01957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xclkbuf_leaf_329_clk clknet_5_4__leaf_clk clknet_leaf_329_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__06079__B _01620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07500_ _03356_ _03374_ _03375_ _00318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09141__A1 net245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08480_ _02713_ _03992_ _01418_ _03993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_77_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05692_ rf_ram.memory\[385\]\[0\] _01787_ _01888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_134_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_59_Left_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07431_ _03323_ _03331_ _03332_ _00292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_3_7_0_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05711__B _01660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07362_ _03260_ _03286_ _03288_ _00267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_169_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_1079 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09101_ _04367_ _04381_ _04383_ _00911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06313_ rf_ram.memory\[188\]\[1\] _01677_ _01793_ rf_ram.memory\[189\]\[1\] _01679_
+ rf_ram.memory\[191\]\[1\] _02508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XANTENNA__06258__A2 _01940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07293_ rf_ram.memory\[468\]\[1\] _03244_ _03246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_143_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09032_ _04331_ _04340_ _04341_ _00884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06244_ _02436_ _02438_ _01790_ _02439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_32_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_60_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_1239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_96_2174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_96_2185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07207__A1 _03190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06175_ rf_ram.memory\[502\]\[1\] _01662_ _01504_ _02370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_29_1061 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_40_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_68_Left_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_57_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_57_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_141_1142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09934_ _04911_ _03135_ _04926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_74_1771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06430__A2 _01863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_111_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_74_1782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09865_ _04840_ _04881_ _04883_ _01176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_176_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_175_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08816_ rf_ram.memory\[137\]\[0\] _04207_ _04208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09796_ _04840_ _04838_ _04841_ _01148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_139_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07930__A2 _03547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08747_ net242 _04152_ _04164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_139_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05959_ _02151_ _02152_ _02153_ _02154_ rf_ram.i_raddr\[3\] _02155_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_68_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_77_Left_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_95_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08678_ rf_ram.memory\[559\]\[0\] _04120_ _04121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_96_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_178_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_165_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07629_ _03355_ _03455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__06497__A2 _01375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output103_I net103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10640_ _00384_ clknet_leaf_92_clk rf_ram.memory\[384\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_119_740 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_165_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_181_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07446__A1 _03323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_153_3234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06249__A2 _01531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10571_ _00315_ clknet_leaf_171_clk rf_ram.memory\[325\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_153_3245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_888 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_107_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_134_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_106_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_114_2506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_114_2517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09199__A1 _02805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_86_Left_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_131_2831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08946__A1 _04266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_1172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_1058 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11123_ _00859_ clknet_leaf_37_clk rf_ram.memory\[11\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06421__A2 _01799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11054_ _00791_ clknet_leaf_9_clk rf_ram.memory\[141\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10005_ _04953_ _04967_ _04969_ _01230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05582__I _01695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_129_2793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_95_Left_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_87_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05932__A1 _01350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_1110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_98_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_969 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07685__A1 _03488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10907_ _00651_ clknet_leaf_19_clk rf_ram.memory\[180\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_86_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_184_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05696__B1 _01773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10838_ _00582_ clknet_leaf_312_clk rf_ram.memory\[537\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_183_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_73_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_15_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_15_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10769_ _00513_ clknet_leaf_304_clk rf_ram.memory\[572\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_70_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_120_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_35_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_262_clk_I clknet_5_17__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_39_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05757__I _01695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_39_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_1148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_188_3875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_188_3886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_188_3897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06412__A2 _01915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_91_2082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07980_ rf_ram.memory\[478\]\[0\] _03673_ _03674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_91_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_277_clk_I clknet_5_16__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06931_ _03014_ _03015_ _03016_ _00108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_129_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_52_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09650_ _03972_ _04737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_06862_ rf_ram.memory\[283\]\[1\] _02967_ _02969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_101_1181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05492__I _01624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08601_ rf_ram.memory\[165\]\[1\] _04071_ _04073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05813_ _02005_ _02006_ _02007_ _02008_ _01860_ _02009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA_clkbuf_leaf_200_clk_I clknet_5_25__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09581_ _03992_ _04693_ _04678_ _04476_ _04694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_59_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06793_ _02868_ _02921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__09114__A1 _04364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08532_ rf_ram.memory\[69\]\[0\] _04028_ _04029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05744_ _01640_ _01940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_78_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_1243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_1254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07676__A1 _03458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08463_ _03971_ _03979_ _03980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06479__A2 _01640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05675_ _01867_ _01868_ _01869_ _01870_ _01658_ _01871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_187_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_175_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_215_clk_I clknet_5_19__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07414_ _03289_ _03320_ _03321_ _00286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_64_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08394_ _03922_ _03930_ _03932_ _00655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_98_2214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_162_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_98_2225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07428__A1 _03326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07345_ _03257_ _03277_ _03278_ _00260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_46_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_30_clk clknet_5_6__leaf_clk clknet_leaf_30_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_92_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_115_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07979__A2 _02917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07276_ rf_ram.memory\[417\]\[0\] _03235_ _03236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_6_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_143_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09015_ rf_ram.memory\[10\]\[1\] _04328_ _04330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06227_ _01603_ _02420_ _02421_ _02422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XTAP_TAPCELL_ROW_76_1811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_1301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05667__I _01633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08928__A1 _04269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input64_I i_ibus_rdt[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_182_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06158_ rf_ram.memory\[489\]\[1\] _01626_ _02353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_112_993 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07600__A1 _03422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06403__A2 _01509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06089_ rf_ram.memory\[334\]\[1\] _01719_ _01707_ _02284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_111_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05611__B1 _01725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_1092 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09917_ _04911_ _03083_ _04915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_97_clk clknet_5_14__leaf_clk clknet_leaf_97_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08156__A2 _03765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09848_ cpu.ctrl.i_jump _01413_ _04870_ _04872_ _04873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06167__A1 _01603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_1127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09779_ _04637_ _04828_ _04830_ _01142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_73_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_107_2387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_969 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_178_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_139_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_165_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_181_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10623_ _00367_ clknet_leaf_102_clk rf_ram.memory\[407\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_10_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06890__A2 _02801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_12_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_load_slew254_I _01361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_21_clk clknet_5_3__leaf_clk clknet_leaf_21_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_187_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_148_1148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10554_ _00298_ clknet_leaf_152_clk rf_ram.memory\[331\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08092__A1 _03724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_1234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_1278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_121_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10485_ _00229_ clknet_leaf_98_clk rf_ram.memory\[418\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_49_1289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08919__A1 _02794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05577__I _01695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08395__A2 _02997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07792__I _03359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_166_3469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05602__B1 _01715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11106_ _00842_ clknet_leaf_118_clk rf_ram.memory\[389\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_34_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_183_3783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_88_clk clknet_5_11__leaf_clk clknet_leaf_88_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_60_1191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_183_3794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09344__A1 net224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09344__B2 net227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11037_ _00774_ clknet_leaf_275_clk rf_ram.i_raddr\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_1175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_155_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05381__A2 _01538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07658__A1 _03455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05460_ _01655_ _01656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_12
XFILLER_0_74_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_89_1036 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_157_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05391_ rf_ram.memory\[574\]\[0\] _01502_ _01506_ _01587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_144_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_12_clk clknet_5_2__leaf_clk clknet_leaf_12_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07130_ _03126_ _03142_ _03144_ _00179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_131_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_31_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08083__A1 _03668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07061_ _03100_ _03101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_93_2122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07830__A1 _03557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_81_clk_I clknet_5_11__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_93_2133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_140_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05487__I _01682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06012_ rf_ram.memory\[536\]\[1\] _01511_ _01552_ _02207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xoutput202 net202 o_ibus_adr[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_70_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput213 net213 o_ibus_adr[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_11_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput224 net224 o_ibus_adr[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_26_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_54_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_96_clk_I clknet_5_14__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07963_ rf_ram.memory\[470\]\[0\] _03662_ _03663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_177_1322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_79_clk clknet_5_11__leaf_clk clknet_leaf_79_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09335__A1 _04463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09702_ _04778_ _01117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06914_ _02775_ _02801_ _03004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07894_ _02836_ _02844_ _03620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09886__A2 _02822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06845_ _02930_ _02955_ _02957_ _00081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09633_ _04524_ net59 _04725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_179_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_78_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09564_ _03992_ net51 _04681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06776_ _02779_ _02837_ _02908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__09638__A2 _01391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_5_1__f_clk_I clknet_3_0_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_69_1681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_154_clk_I clknet_5_26__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08515_ rf_ram.memory\[172\]\[0\] _04017_ _04018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_33_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05727_ _01550_ _01923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_09495_ _01442_ _01342_ _04630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_33_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_175_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08446_ _03953_ _03964_ _03965_ _00674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_77_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_34_clk_I clknet_5_6__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05658_ _01851_ _01853_ _01790_ _01854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_148_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_102_2284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_102_2295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_175_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_162_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_849 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_1322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08377_ _03689_ _03922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_68_1109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05589_ _01686_ _01785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA_clkbuf_leaf_169_clk_I clknet_5_30__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07328_ _02958_ _02954_ _03268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_144_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06085__B1 _01656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_49_clk_I clknet_5_12__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07259_ _03222_ _03223_ _03224_ _00228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07821__A1 _02761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06624__A2 _02730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05832__B1 _01959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10270_ _00014_ clknet_leaf_277_clk rf_ram.memory\[233\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_output170_I net170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_131_598 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_148_3144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_107_clk_I clknet_5_15__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_109_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05346__B _01528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_109_2427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_126_2730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_126_2741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_161_3377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07888__A1 _02959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_161_3388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06560__A1 _01369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05363__A2 _01538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_17_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09629__A2 net55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_17_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06177__B _01526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_154_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11655_ net105 net177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_65_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05520__C1 _01715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10606_ _00350_ clknet_leaf_154_clk rf_ram.memory\[316\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11586_ _01318_ clknet_leaf_284_clk rf_ram.memory\[237\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_49_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_181_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06615__A2 _02788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10537_ _00281_ clknet_leaf_212_clk rf_ram.memory\[248\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_10_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_168_3509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10468_ _00212_ clknet_leaf_195_clk rf_ram.memory\[260\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_185_3823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_185_3834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09565__A1 _03992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08368__A2 _03903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10399_ _00143_ clknet_leaf_302_clk rf_ram.memory\[218\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06379__A1 _01768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09317__A1 _04526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09317__B2 cpu.immdec.imm11_7\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_1_clk clknet_5_1__leaf_clk clknet_leaf_1_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__06000__B1 _01539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06630_ _02795_ _02801_ _02802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06866__I _02971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_1057 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06551__A1 _02731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_1079 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_177_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06561_ _01353_ rf_ram_if.wdata1_r\[1\] _02745_ _02746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08300_ _03852_ _03872_ _03873_ _00620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_158_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05512_ rf_ram.memory\[326\]\[0\] _01706_ _01707_ _01708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09280_ cpu.genblk3.csr.mcause3_0\[3\] _01341_ cpu.genblk3.csr.o_new_irq _01391_
+ _04502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_129_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_47_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06492_ _02603_ _02630_ _01372_ _02686_ _02687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_145_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_185_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08231_ _03798_ _02866_ _03831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05443_ _01612_ _01621_ _01630_ _01638_ _01639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_144_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06854__A2 _02941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_28_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08056__A1 _03134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08162_ net237 _03765_ _03788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05374_ _01351_ _01547_ _01566_ _01569_ _01570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_173_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_1131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_160_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07113_ _03126_ _03131_ _03133_ _00173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_67_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07803__A1 _03554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08093_ _02843_ _03729_ _03745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06606__A2 _02781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_1321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07044_ _02829_ _03089_ _03090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_113_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05290__A1 _01434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05578__C1 _01773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08995_ rf_ram.memory\[113\]\[1\] _04316_ _04318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07946_ _02728_ _02832_ _03652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05593__A2 _01785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06790__A1 _02873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_143_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input27_I i_dbus_rdt[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07877_ _03590_ _03607_ _03609_ _00461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_3_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08477__B net65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_3_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_1255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08531__A2 _04005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09616_ rf_ram.memory\[72\]\[1\] _04717_ _04719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_183_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06828_ _02945_ _02946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_104_2324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05345__A2 _01538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_104_2335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_168_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06759_ _02873_ _02895_ _02896_ _00056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09547_ _04478_ net43 _04650_ cpu.immdec.imm19_12_20\[7\] _04668_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_149_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_84_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_84_1965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07098__A2 _02946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08295__A1 _03852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09478_ _02703_ _02705_ _04615_ _04616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_4_1231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_110_1022 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08429_ rf_ram.memory\[59\]\[0\] _03954_ _03955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_53_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11440_ _01172_ clknet_leaf_241_clk cpu.mem_bytecnt\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_4
XANTENNA__08047__A1 _03686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_110_1077 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_117_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08598__A2 _04067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_1196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11371_ _01103_ clknet_leaf_236_clk net134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_85_1253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_841 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05805__B1 _01516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10322_ _00066_ clknet_leaf_288_clk rf_ram.memory\[50\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_104_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09547__A1 _04478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10253_ _02825_ _05119_ _05121_ _01326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_5_29__f_clk clknet_3_7_0_clk clknet_5_29__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__10157__A2 _02921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_163_3417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10184_ rf_ram.memory\[190\]\[0\] _05079_ _05080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_163_3428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_180_3731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_180_3742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05584__A2 _01777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_89_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06686__I _02845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05590__I _01695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_186_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_97_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_178_3693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_1310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_139_2976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_154_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11638_ net89 net162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_182_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_42_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_170_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11569_ _01301_ clknet_leaf_285_clk rf_ram.memory\[238\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09438__S _04593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09665__C _04740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05272__A1 cpu.ctrl.pc vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09538__A1 _04526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_1170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_1181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_1061 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06370__B _01684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07800_ _03557_ _03560_ _03562_ _00431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08780_ rf_ram.memory\[142\]\[1\] _04183_ _04185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05992_ _01371_ _02187_ _02188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_127_Right_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05575__A2 _01770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_88_2032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_88_2043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07731_ rf_ram.memory\[397\]\[0\] _03518_ _03519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05980__C1 _01653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_49_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09710__A1 _04781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07662_ rf_ram.memory\[385\]\[0\] _03475_ _03476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_0_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_49_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_40_Left_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_137_1180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09401_ _04573_ _01021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06613_ _02716_ _02786_ _02787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_88_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_177_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07593_ _02935_ _02822_ _03433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_177_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09332_ _04466_ _04533_ _04535_ _00990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06544_ _01347_ _01366_ _02730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__08277__A1 _03855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_1077 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_158_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10084__A1 _05017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09263_ _01484_ _04489_ _04490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_62_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_1196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_62_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06475_ rf_ram.memory\[30\]\[1\] _01530_ _02670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_47_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_161_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08214_ _03685_ _03820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_05426_ rf_ram.memory\[360\]\[0\] _01614_ _01615_ _01622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_8_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08029__A1 _03690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09194_ net236 _04418_ _04442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_16_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_161_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06264__C _01569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08145_ _03757_ _03775_ _03777_ _00561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09777__A1 _04634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_181_1318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_172_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05357_ rf_ram.memory\[528\]\[0\] _01511_ _01552_ _01553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_16_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08076_ rf_ram.memory\[561\]\[1\] _03733_ _03735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05288_ _01389_ _01341_ _01485_ cpu.o_wdata1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_70_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07027_ rf_ram.memory\[218\]\[1\] _03076_ _03078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06460__B1 _01518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_1270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_101_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_1146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_8_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08201__A1 _03787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_1134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_1178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08978_ rf_ram.memory\[116\]\[0\] _04307_ _04308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05566__A2 _01644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output133_I net133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07929_ _03622_ _03639_ _03641_ _00481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09701__A1 net99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10940_ _00678_ clknet_leaf_256_clk rf_ram_if.rgnt vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_39_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06515__A1 cpu.alu.i_rs1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_1074 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_79_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10871_ _00615_ clknet_leaf_34_clk rf_ram.memory\[204\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_168_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_94_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_94_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_39_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_1188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_155_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10075__A1 _04982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_93_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_156_3287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_156_3298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_152_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_151_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11423_ _01155_ clknet_leaf_294_clk rf_ram.memory\[7\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_46_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11354_ _01086_ clknet_leaf_280_clk cpu.immdec.imm24_20\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_104_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_134_2884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10305_ _00049_ clknet_leaf_268_clk rf_ram.memory\[518\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_46_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11285_ _01020_ clknet_leaf_242_clk net221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10236_ _02819_ _05110_ _05111_ _01319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_20_1207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06203__B1 _01725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10167_ _02908_ _03547_ _05069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06754__A1 _02876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05557__A2 _01644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10098_ rf_ram.memory\[351\]\[1\] _05025_ _05027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_88_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_156_1055 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_156_1066 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_1077 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_107_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_1039 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_1174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_1054 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_1027 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_1169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_128_911 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_44_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_44_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_174_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_106_Left_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_44_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06260_ rf_ram.memory\[416\]\[1\] _01755_ _01756_ _02455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_26_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_127_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05211_ _01401_ _01403_ _01404_ _01410_ _01411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_4
XANTENNA__09759__A1 net118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_1124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09759__B2 net119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06191_ rf_ram.memory\[474\]\[1\] _01856_ _01786_ rf_ram.memory\[475\]\[1\] _02385_
+ _02386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_170_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_170_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_68_1281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_163_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05142_ _01334_ _01337_ _01344_ cpu.immdec.imm24_20\[0\] _01345_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_64_1123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_292_clk clknet_5_24__leaf_clk clknet_leaf_292_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09950_ rf_ram.memory\[337\]\[0\] _04935_ _04936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08982__A2 _04303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_3_3_0_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05796__A2 _01846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08901_ _04237_ _04257_ _04259_ _00835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09881_ _03309_ _02795_ _04893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_110_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_5_12__f_clk clknet_3_3_0_clk clknet_5_12__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_5_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09931__A1 _04918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08832_ _04202_ _04216_ _04217_ _00808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05548__A2 _01697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_178_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_139_1242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08763_ rf_ram.memory\[145\]\[0\] _04174_ _04175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05975_ _01903_ _02169_ _02170_ _02171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_140_3000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05953__C1 _01655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_1098 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07714_ _03491_ _03506_ _03508_ _00399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08498__A1 _02736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08694_ _02983_ _04078_ _04131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_36_1214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09631__S _04526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07645_ _03458_ _03463_ _03465_ _00373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_79_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_81_1902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_81_1913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07576_ _03355_ _03422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_137_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10057__A1 _04985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06527_ _02713_ _02714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_24_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09315_ _04525_ _00983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_75_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09998__A1 _04950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_24_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06275__B _01956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_180_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09246_ _02714_ _04475_ _00964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06458_ rf_ram.memory\[52\]\[1\] _01508_ _01655_ rf_ram.memory\[53\]\[1\] _01518_
+ rf_ram.memory\[55\]\[1\] _02653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_63_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_1172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_1280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_185_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_17_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05409_ _01499_ _01605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_146_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09177_ _04396_ _04431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_06389_ rf_ram.memory\[65\]\[1\] _01918_ _02584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_161_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08128_ _03754_ _03766_ _03767_ _00554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_43_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_79_1864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08422__A1 net243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_79_1875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_151_3195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_120_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_283_clk clknet_5_18__leaf_clk clknet_leaf_283_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08059_ _03689_ _03724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__05787__A2 _01922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_179_1000 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_112_2478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11070_ _00807_ clknet_leaf_15_clk rf_ram.memory\[135\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_101_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput68 net68 o_dbus_adr[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput79 net79 o_dbus_adr[22] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_10021_ _03309_ _03009_ _04979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06736__A1 _02873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_98_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10923_ _00667_ clknet_leaf_4_clk rf_ram.memory\[173\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_19_Right_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07161__A1 _03157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_158_3327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_158_3338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10854_ _00598_ clknet_leaf_297_clk rf_ram.memory\[52\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_184_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_156_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_175_3641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10048__A1 _03445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_175_3652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_183_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10785_ _00529_ clknet_leaf_326_clk rf_ram.memory\[564\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_82_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06185__B _01693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_136_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_137_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_136_2924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08661__A1 _04097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07464__A2 _02904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06121__C1 _01668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_1107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_164_1313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07795__I _03088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11406_ _01138_ clknet_leaf_233_clk net122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__07216__A2 _02941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09461__I0 net80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_10_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_151_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_28_Right_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_10_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_775 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_274_clk clknet_5_16__leaf_clk clknet_leaf_274_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_11337_ _01069_ clknet_leaf_217_clk cpu.immdec.imm19_12_20\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_22_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05778__A2 _01649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11268_ _01003_ clknet_leaf_248_clk net203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_123_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_37_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_37_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10219_ _02996_ _03082_ _05101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_11199_ _00935_ clknet_leaf_49_clk rf_ram.memory\[87\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_118_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_1236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_1127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05935__C1 _01607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_89_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05760_ _01526_ _01956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_178_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_37_Right_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07035__I net235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05950__A2 _01633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09141__A2 _04005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05691_ rf_ram.memory\[384\]\[0\] _01782_ _01783_ _01887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07430_ rf_ram.memory\[370\]\[0\] _03331_ _03332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_76_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_1172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_1003 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_119_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05702__A2 _01614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_114_Left_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_187_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07361_ rf_ram.memory\[268\]\[1\] _03286_ _03288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_73_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06312_ rf_ram.memory\[190\]\[1\] _01641_ _02004_ _02507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09100_ rf_ram.memory\[96\]\[1\] _04381_ _04383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_72_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07292_ _03222_ _03244_ _03245_ _00240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08652__A1 net237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09031_ rf_ram.memory\[106\]\[0\] _04340_ _04341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06243_ rf_ram.memory\[434\]\[1\] _01856_ _01857_ rf_ram.memory\[435\]\[1\] _02437_
+ _02438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_115_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_969 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_46_Right_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_60_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_96_2175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_1040 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08404__A1 _03922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_96_2186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06174_ _02367_ _02368_ _01629_ _02369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__09452__I0 net76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_980 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_130_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_265_clk clknet_5_17__leaf_clk clknet_leaf_265_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__10211__A1 _05078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05769__A2 _01958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_57_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06966__A1 _03018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_123_Left_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_57_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09933_ _04921_ _04923_ _04925_ _01202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_99_1016 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_74_1772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_74_1783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09864_ rf_ram.memory\[5\]\[1\] _04881_ _04883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08815_ net249 _04195_ _04207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_99_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09795_ rf_ram.memory\[80\]\[1\] _04838_ _04841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06194__A2 _01863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_55_Right_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08746_ _04157_ _04163_ _00776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05958_ rf_ram.memory\[50\]\[0\] _01499_ _01653_ rf_ram.memory\[51\]\[0\] _01655_
+ rf_ram.memory\[49\]\[0\] _02154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XANTENNA__05941__A2 _01682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_132_Left_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08677_ _02953_ _03765_ _04120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_68_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07143__A1 _03123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05889_ _02082_ _02084_ _01978_ _02085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_178_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_1055 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07628_ _03425_ _03452_ _03454_ _00367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_49_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05902__B _01602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08891__A1 _04237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07559_ rf_ram.memory\[358\]\[1\] _03410_ _03412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_119_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10570_ _00314_ clknet_leaf_163_clk rf_ram.memory\[325\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_153_3235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_64_Right_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_17_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09229_ _04396_ _04463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_170_3560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_114_2507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_114_2518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09199__A2 _04418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_141_Left_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_133_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_131_2821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_131_2832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_256_clk clknet_5_20__leaf_clk clknet_leaf_256_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_102_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_31_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11122_ _00858_ clknet_leaf_37_clk rf_ram.memory\[11\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_7_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_120_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11053_ _00790_ clknet_leaf_9_clk rf_ram.memory\[141\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06709__A1 _02820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_73_Right_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10004_ rf_ram.memory\[504\]\[1\] _04967_ _04969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07382__A1 _03289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06185__A2 _01782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_129_2794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_639 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_1264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10906_ _00650_ clknet_leaf_19_clk rf_ram.memory\[180\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08882__A1 net240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09070__I _04057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10837_ _00581_ clknet_leaf_314_clk rf_ram.memory\[538\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_144_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_82_Right_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_15_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_184_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_880 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08634__A1 _04062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10768_ _00512_ clknet_leaf_327_clk rf_ram.memory\[572\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_137_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10699_ _00443_ clknet_leaf_91_clk rf_ram.memory\[412\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_23_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05999__A2 _01502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_563 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_140_703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_39_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_247_clk clknet_5_21__leaf_clk clknet_leaf_247_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_140_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_39_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_188_3876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06948__A1 _03014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_188_3887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_188_3898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09446__S _04593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_1279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_91_2083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_91_2094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05620__A1 net252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_91_Right_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06930_ rf_ram.memory\[297\]\[0\] _03015_ _03016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_129_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_180_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_input1_I i_dbus_ack vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_52_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06861_ _02927_ _02967_ _02968_ _00086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05908__C1 _01931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06176__A2 _01509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08600_ _04058_ _04071_ _04072_ _00721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05812_ rf_ram.memory\[184\]\[0\] _01711_ _01848_ rf_ram.memory\[185\]\[0\] _01773_
+ rf_ram.memory\[187\]\[0\] _02008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_179_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09580_ _01391_ _01469_ cpu.immdec.imm7 _04691_ _04692_ _04693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_06792_ _02876_ _02918_ _02920_ _00065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05923__A2 _01677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_175_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_59_1099 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05743_ _01935_ _01936_ _01937_ _01938_ _01658_ _01939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_08531_ _02794_ _04005_ _04028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_72_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07125__A1 _03126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08462_ _03972_ _03978_ _03979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05674_ rf_ram.memory\[456\]\[0\] _01724_ _01725_ rf_ram.memory\[457\]\[0\] _01726_
+ rf_ram.memory\[459\]\[0\] _01870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_07413_ rf_ram.memory\[334\]\[0\] _03320_ _03321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08393_ rf_ram.memory\[199\]\[1\] _03930_ _03932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_163_806 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_98_2215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07344_ rf_ram.memory\[253\]\[0\] _03277_ _03278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_98_2226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08625__A1 _02821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_128_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07275_ _02899_ _03234_ _03235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_182_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06100__A2 _01614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06226_ rf_ram.memory\[412\]\[1\] _01634_ _01702_ rf_ram.memory\[413\]\[1\] _01608_
+ rf_ram.memory\[415\]\[1\] _02421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_143_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09014_ _04298_ _04328_ _04329_ _00878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_103_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_76_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_238_clk clknet_5_21__leaf_clk clknet_leaf_238_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_131_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06157_ rf_ram.memory\[488\]\[1\] _01683_ _01684_ _02352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09050__A1 _02805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input57_I i_ibus_rdt[31] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_983 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06088_ _02279_ _02280_ _02281_ _02282_ _01717_ _02283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_106_1071 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09916_ _04887_ _04912_ _04914_ _01196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_leaf_8_clk_I clknet_5_0__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09847_ _01382_ _04871_ _01391_ _04872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07364__A1 _03055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09778_ rf_ram.memory\[77\]\[1\] _04828_ _04830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05914__A2 _01915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output213_I net213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08729_ _04077_ _04152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_107_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07116__A1 _02915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_107_2388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_179_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_95_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_322_clk_I clknet_5_4__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05632__B _01620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_124_2691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11671_ cpu.ctrl.pc net202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_48_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_181_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10622_ _00366_ clknet_leaf_102_clk rf_ram.memory\[407\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_37_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_12_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_337_clk_I clknet_5_0__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_984 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_744 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_1273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10553_ _00297_ clknet_leaf_130_clk rf_ram.memory\[36\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_91_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_1148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10484_ _00228_ clknet_leaf_98_clk rf_ram.memory\[418\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_229_clk clknet_5_23__leaf_clk clknet_leaf_229_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_121_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08919__A2 _03559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05850__A1 _01674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11105_ _00841_ clknet_leaf_79_clk rf_ram.memory\[439\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_34_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_34_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_183_3784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09344__A2 _03991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_183_3795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_159_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11036_ _00773_ clknet_leaf_278_clk rf_ram_if.rtrig0 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07355__A1 _03257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06158__A2 _01626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08855__A1 net240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06315__C1 _01773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05669__A1 _01769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06330__A2 _01804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_1026 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_845 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05390_ _01582_ _01583_ _01584_ _01585_ _01495_ _01586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__08607__A1 _04062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_172_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_166_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_82_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_153_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_31_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08083__A2 _03083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06373__B _02004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06094__A1 _01349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07060_ _02764_ _02799_ _03100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_125_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_93_2123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_152_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_93_2134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06011_ rf_ram.memory\[540\]\[1\] _01538_ _01555_ rf_ram.memory\[541\]\[1\] _01554_
+ rf_ram.memory\[543\]\[1\] _02206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
Xoutput203 net203 o_ibus_adr[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_113_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09032__A1 _04331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput214 net214 o_ibus_adr[20] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput225 net225 o_ibus_adr[30] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_140_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_54_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06397__A2 _01711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_71_1720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07962_ _02836_ _03009_ _03662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09701_ net99 _04767_ _04768_ net100 _04777_ _04778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_06913_ _02975_ _03001_ _03003_ _00103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07893_ _03355_ _03619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_09632_ _04724_ _01101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06844_ rf_ram.memory\[303\]\[1\] _02955_ _02957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_78_701 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09563_ cpu.immdec.imm30_25\[2\] _04680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09099__A1 _04364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06775_ _02876_ _02905_ _02907_ _00061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_78_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08514_ _02787_ _03949_ _04017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_69_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05726_ _01536_ _01922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_09494_ _01439_ _04625_ _04627_ _04629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_147_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_1074 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08445_ rf_ram.memory\[176\]\[0\] _03964_ _03965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_72_1096 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_92_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05657_ rf_ram.memory\[466\]\[0\] _01785_ _01778_ rf_ram.memory\[467\]\[0\] _01852_
+ _01853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_18_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_102_2285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_102_2296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05588_ rf_ram.memory\[288\]\[0\] _01782_ _01783_ _01784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08376_ _03919_ _03920_ _03921_ _00648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_147_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07327_ _03260_ _03265_ _03267_ _00253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09271__A1 _01364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_116_563 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_150_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07258_ rf_ram.memory\[418\]\[0\] _03223_ _03224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07821__A2 _03234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_103_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06209_ _01368_ _02376_ _02403_ _02404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_07189_ _02836_ _02984_ _03181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09023__A1 _04334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_1121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07893__I _03355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_1177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07585__A1 _03422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_148_3145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06388__A2 _01922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_109_2417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_109_2428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07337__A1 _03260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_126_2731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_126_2742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07888__A2 _03234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_161_3378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_161_3389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_159_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_261_clk_I clknet_5_17__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_17_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_115_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05362__B _01505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08837__A1 _04202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_1245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_1158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06312__A2 _01641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_1289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_139_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_276_clk_I clknet_5_16__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05520__B1 _01713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11654_ net104 net176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_181_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_83_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_984 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_181_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10605_ _00349_ clknet_leaf_157_clk rf_ram.memory\[356\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_36_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_921 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09262__A1 _01461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11585_ _01317_ clknet_leaf_284_clk rf_ram.memory\[237\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_107_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10536_ _00280_ clknet_leaf_212_clk rf_ram.memory\[248\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_122_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09014__A1 _04298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_108_Right_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_110_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10467_ _00211_ clknet_leaf_195_clk rf_ram.memory\[261\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_185_3824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_185_3835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10398_ _00142_ clknet_leaf_302_clk rf_ram.memory\[218\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_20_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_214_clk_I clknet_5_19__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09317__A2 net64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07328__A1 _02958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11019_ _00756_ clknet_leaf_330_clk rf_ram.memory\[154\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_126_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_229_clk_I clknet_5_23__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06551__A2 _02736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06368__B _02004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06560_ _01369_ rf_ram_if.wdata0_r\[1\] _02745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_59_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_172_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07043__I _03088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_157_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05511_ _01503_ _01707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_06491_ net252 _02658_ _02685_ _02686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XTAP_TAPCELL_ROW_47_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_173_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07500__A1 _03356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05442_ _01527_ _01632_ _01637_ _01638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_08230_ _03823_ _03828_ _03830_ _00593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_145_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_64_1590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08161_ _03685_ _03787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_05373_ _01568_ _01569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__08056__A2 _03693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09253__A1 _01366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_126_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07112_ rf_ram.memory\[488\]\[1\] _03131_ _03133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08092_ _03724_ _03742_ _03744_ _00541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_127_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07043_ _03088_ _03089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_30_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_67_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05578__B1 _01772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08994_ _04298_ _04316_ _04317_ _00870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_48_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07945_ _03355_ _03651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_138_1115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_177_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_143_3053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_1212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07876_ rf_ram.memory\[463\]\[1\] _03607_ _03609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_3_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09615_ _04634_ _04717_ _04718_ _01090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06827_ _02716_ _02759_ _02945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_74_1136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_104_2325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06278__B _01494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_104_2336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09546_ cpu.immdec.imm19_12_20\[8\] _04667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_92_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_5_28__f_clk_I clknet_3_7_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06758_ rf_ram.memory\[514\]\[0\] _02895_ _02896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08819__A1 _04205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_84_1955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_121_2650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_84_1966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05709_ rf_ram.memory\[402\]\[0\] _01500_ _01763_ rf_ram.memory\[403\]\[0\] _01656_
+ rf_ram.memory\[401\]\[0\] _01905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_65_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09477_ _02703_ _02705_ _03989_ _04615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_78_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06689_ _02820_ _02847_ _02848_ _00034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_65_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_176_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_163_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05910__B _01916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08428_ _02822_ _02869_ _03954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_109_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_188_1260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_175_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_163_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_93_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_164_956 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08359_ rf_ram.memory\[183\]\[0\] _03910_ _03911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_62_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_184_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06058__A1 _01527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11370_ _01102_ clknet_leaf_235_clk cpu.decode.opcode\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_150_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10321_ _00065_ clknet_leaf_221_clk rf_ram.memory\[510\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_131_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output88_I net88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09547__A2 net43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05281__A2 _01478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10252_ rf_ram.memory\[28\]\[1\] _05119_ _05121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07558__A1 _03389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05357__B _01552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10183_ _02916_ _03902_ _05079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_163_3418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_163_3429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_1174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_180_3732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_180_3743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_1110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07730__A1 _02844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_80_clk_I clknet_5_11__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06188__B _01790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_9_1198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_178_3694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_155_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_95_clk_I clknet_5_14__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_1322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_155_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_139_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09235__A1 _04466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11637_ net88 net161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_53_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_182_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11568_ _01300_ clknet_leaf_25_clk rf_ram.memory\[190\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_53_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_122_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10519_ _00263_ clknet_leaf_209_clk rf_ram.memory\[26\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11499_ _01231_ clknet_leaf_178_clk rf_ram.memory\[277\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09538__A2 net39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_153_clk_I clknet_5_26__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_33_clk_I clknet_5_6__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09454__S _04593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05991_ _02017_ _02074_ _02186_ _01373_ _02187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XPHY_EDGE_ROW_179_Left_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_88_2033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07730_ _02844_ _03481_ _03518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_168_clk_I clknet_5_30__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05980__B1 _01714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07661_ net238 _03089_ _03475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_49_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09710__A2 net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_48_clk_I clknet_5_12__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06524__A2 _02709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_1170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09400_ net222 _03990_ _04564_ net223 _04573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06612_ _02785_ _02725_ _02786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_07592_ _03425_ _03430_ _03432_ _00353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_172_1072 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_137_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_66_1630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09331_ rf_ram.memory\[309\]\[1\] _04533_ _04535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06543_ cpu.immdec.imm11_7\[4\] _02729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_87_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_1089 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_1164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09262_ _01461_ _04487_ _04488_ _04489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_62_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_173_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06474_ _02666_ _02668_ _01563_ _02669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_28_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_188_Left_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_44_921 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08213_ _03790_ _03817_ _03819_ _00587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05425_ _01616_ _01619_ _01620_ _01621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_172_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_106_clk_I clknet_5_15__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09226__A1 _04431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09193_ _04434_ _04439_ _04441_ _00945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_28_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_173_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08144_ rf_ram.memory\[548\]\[1\] _03775_ _03777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_44_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05356_ _01551_ _01552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_71_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05287_ _01341_ _01484_ _01485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08075_ _03721_ _03733_ _03734_ _00534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_144_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05263__A2 _01460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07026_ _03050_ _03076_ _03077_ _00142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_140_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_8_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_1184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08201__A2 _03811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06212__A1 _01769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08977_ _03134_ _04303_ _04307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06787__I _02916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05905__B _01660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07928_ rf_ram.memory\[458\]\[1\] _03639_ _03641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05971__B1 _01624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output126_I net126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07859_ rf_ram.memory\[40\]\[0\] _03598_ _03599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07712__A1 _03488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_1112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10870_ _00614_ clknet_leaf_34_clk rf_ram.memory\[204\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_97_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_149_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09529_ cpu.immdec.imm19_12_20\[2\] _04654_ _04656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_13_1204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05640__B _01756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_1248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07411__I _02814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_1073 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_156_3288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_156_3299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_188_1090 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_164_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11422_ _01154_ clknet_leaf_35_clk rf_ram.memory\[74\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_123_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09768__A2 _04766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11353_ _01085_ clknet_leaf_216_clk cpu.immdec.imm24_20\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_105_875 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_134_2885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06471__B _01550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10304_ _00048_ clknet_leaf_269_clk rf_ram.memory\[518\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11284_ _01019_ clknet_leaf_243_clk net220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10235_ rf_ram.memory\[208\]\[0\] _05110_ _05111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_20_1219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10166_ _05049_ _05066_ _05068_ _01292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07951__A1 _03654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10097_ _05014_ _05025_ _05026_ _01265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_89_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05534__C _01361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_1022 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_1164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_186_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10999_ _00736_ clknet_leaf_334_clk rf_ram.memory\[162\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_44_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_139_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_155_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_910 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09208__A1 _04434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05210_ _01408_ _01409_ _01410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_170_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05493__A2 _01626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09759__A2 _04766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06190_ rf_ram.memory\[473\]\[1\] _01787_ _02385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XPHY_EDGE_ROW_160_Right_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_154_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_130_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05141_ _01343_ _01336_ cpu.state.genblk1.misalign_trap_sync_r cpu.genblk3.csr.o_new_irq
+ _01344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_128_1169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xmax_cap235 _03082_ net235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__09248__I net34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05776__I _01615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xmax_cap246 _02780_ net246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_64_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08900_ rf_ram.memory\[429\]\[1\] _04257_ _04259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09880_ _04887_ _04890_ _04892_ _01182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09392__B1 _04564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08831_ rf_ram.memory\[459\]\[0\] _04216_ _04217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_100_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07942__A1 _03619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05725__B _01790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08762_ _02760_ _04152_ _04174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05953__B1 _01653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05974_ rf_ram.memory\[28\]\[0\] _01633_ _01617_ rf_ram.memory\[29\]\[0\] _01607_
+ rf_ram.memory\[31\]\[0\] _02170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XTAP_TAPCELL_ROW_140_3001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07713_ rf_ram.memory\[3\]\[1\] _03506_ _03508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08693_ _04129_ _04127_ _04130_ _00756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09695__A1 net128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08498__A2 _02867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_1204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09695__B2 net129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_1106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07644_ rf_ram.memory\[387\]\[1\] _03463_ _03465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_73_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_81_1903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07575_ _03393_ _03419_ _03421_ _00347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_119_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09314_ _04524_ net63 _04521_ cpu.immdec.imm11_7\[2\] _04522_ cpu.immdec.imm11_7\[1\]
+ _04525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_06526_ net65 _02713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XTAP_TAPCELL_ROW_24_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05469__C1 _01519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_921 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09245_ cpu.genblk3.csr.o_new_irq _01413_ _04473_ _04474_ _04475_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06457_ rf_ram.memory\[54\]\[1\] _01661_ _01503_ _02652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_119_989 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06130__B1 _01778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_173_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_146_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05408_ rf_ram.memory\[356\]\[0\] _01537_ _01604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05484__A2 _01677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_1292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09176_ _04401_ _04428_ _04430_ _00939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_32_913 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06388_ rf_ram.memory\[64\]\[1\] _01922_ _01551_ _02583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_105_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_160_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_160_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08127_ rf_ram.memory\[551\]\[0\] _03766_ _03767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_82_1213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05339_ rf_ram.memory\[518\]\[0\] _01502_ _01506_ _01535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_79_1865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_116_2560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_151_3196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08422__A2 _03949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_79_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08058_ _03721_ _03722_ _03723_ _00528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05619__C net253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07009_ _03050_ _03065_ _03066_ _00136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05641__C1 _01715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_112_2479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput69 net69 o_dbus_adr[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__08186__A1 _03787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10020_ _04953_ _04976_ _04978_ _01236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_122_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_1310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_99_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_169_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10922_ _00666_ clknet_leaf_5_clk rf_ram.memory\[173\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_58_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_158_3328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10853_ _00597_ clknet_leaf_309_clk rf_ram.memory\[530\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05172__A1 _01351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_175_3642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10048__A2 _02923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05370__B _01351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10784_ _00528_ clknet_leaf_325_clk rf_ram.memory\[564\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_52_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_136_2914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_136_2925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_1135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06121__B1 _01519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_109_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_425 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_164_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11405_ _01137_ clknet_leaf_230_clk net121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05880__C1 _02019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_946 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09610__A1 _04634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09461__I1 net81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_10_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11336_ _01068_ clknet_leaf_218_clk cpu.immdec.imm19_12_20\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_50_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_162_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11267_ _01002_ clknet_leaf_248_clk net233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_123_1066 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08177__A1 _03790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_1077 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10218_ _05081_ _05098_ _05100_ _01312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_37_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_37_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11198_ _00934_ clknet_leaf_49_clk rf_ram.memory\[87\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_59_1204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07924__A1 _03622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10149_ _05046_ _05057_ _05058_ _01285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05935__B1 _01609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_1139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_171_1318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05690_ _01883_ _01885_ _01746_ _01886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_89_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_159_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05163__A1 _01364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_174_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_174_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_1101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_1112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07360_ _03257_ _03286_ _03287_ _00266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_128_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06095__C _01361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06311_ _02494_ _02498_ _02502_ _02505_ _02506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_72_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07291_ rf_ram.memory\[468\]\[0\] _03244_ _03245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08652__A2 _04067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09030_ net247 _04339_ _04340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06242_ rf_ram.memory\[433\]\[1\] _01787_ _02437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__06663__A1 _02826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_96_2176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_130_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_96_2187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06173_ rf_ram.memory\[506\]\[1\] _01652_ _01654_ rf_ram.memory\[507\]\[1\] _01715_
+ rf_ram.memory\[505\]\[1\] _02368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_13_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09452__I1 net77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_170_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_141_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_57_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05623__C1 _01679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09932_ rf_ram.memory\[341\]\[1\] _04923_ _04925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_110_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_1144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08168__A1 _02881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_74_1773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_1028 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_74_1784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_110_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_1139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09863_ _04837_ _04881_ _04882_ _01175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07915__A1 _02844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08814_ _04205_ _04203_ _04206_ _00801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05455__B _01650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09794_ _04400_ _04840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_30_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08745_ _01495_ _04160_ _04163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__09668__A1 net120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05957_ rf_ram.memory\[48\]\[0\] _01633_ _01525_ _02153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08676_ _04097_ _04117_ _04119_ _00750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_68_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_1072 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05888_ rf_ram.memory\[66\]\[0\] _01804_ _02019_ rf_ram.memory\[67\]\[0\] _02083_
+ _02084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__08340__A1 _03887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07627_ rf_ram.memory\[407\]\[1\] _03452_ _03454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_36_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05154__A1 _01347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06286__B _01923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07558_ _03389_ _03410_ _03411_ _00340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_165_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06509_ _02697_ _02698_ _02696_ _00006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_181_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_701 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_180_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07489_ rf_ram.memory\[325\]\[0\] _03368_ _03369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_153_3236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09228_ _04434_ _04460_ _04462_ _00959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_107_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_170_3550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output193_I net193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_114_2508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_114_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_146_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09159_ _04397_ _04419_ _04420_ _00932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_115_970 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_131_2822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_131_2833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_82_1054 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11121_ _00857_ clknet_leaf_85_clk rf_ram.memory\[120\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_82_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_43_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output70_I net70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11052_ _00789_ clknet_leaf_6_clk rf_ram.memory\[142\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_101_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10003_ _04950_ _04967_ _04968_ _01229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_129_2784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_129_2795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09659__A1 net120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_1124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_99_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_1146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_28_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_1243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_153_1059 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08331__A1 _03892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10905_ _00649_ clknet_leaf_19_clk rf_ram.memory\[186\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_129_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_192_clk clknet_5_30__leaf_clk clknet_leaf_192_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_15_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_1167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_156_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08882__A2 _03547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05696__A2 _01777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10836_ _00580_ clknet_leaf_270_clk rf_ram.memory\[538\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_95_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_184_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_184_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_184_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_15_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10767_ _00511_ clknet_leaf_327_clk rf_ram.memory\[573\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09831__A1 _04840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10698_ _00442_ clknet_leaf_91_clk rf_ram.memory\[412\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_152_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_1242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_125_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_50_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_1252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_39_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_39_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_188_3877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_188_3888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_188_3899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11319_ _01052_ clknet_leaf_263_clk net84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_121_984 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_91_2084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_91_2095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09898__A1 _04884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06860_ rf_ram.memory\[283\]\[0\] _02967_ _02968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_52_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05908__B1 _01911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_173_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08570__A1 _04023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05811_ rf_ram.memory\[186\]\[0\] _01641_ _01916_ _02007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_175_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06791_ rf_ram.memory\[510\]\[1\] _02918_ _02920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_136_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08530_ _04026_ _04024_ _04027_ _00696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05742_ rf_ram.memory\[424\]\[0\] _01666_ _01810_ rf_ram.memory\[425\]\[0\] _01811_
+ rf_ram.memory\[427\]\[0\] _01938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_145_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_148_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08461_ cpu.bufreg2.o_sh_done_r _03977_ _03978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_72_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05673_ rf_ram.memory\[458\]\[0\] _01719_ _01650_ _01869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_148_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_183_clk clknet_5_29__leaf_clk clknet_leaf_183_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_159_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07412_ _03319_ _02972_ _03320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05687__A2 _01782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08392_ _03919_ _03930_ _03931_ _00654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_169_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07343_ _03055_ _02960_ _03277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_73_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_98_2216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_98_2227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_174_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_162_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08625__A2 _02881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09822__A1 _03309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07274_ _03039_ _03234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_33_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_851 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09013_ rf_ram.memory\[10\]\[0\] _04328_ _04329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06225_ rf_ram.memory\[414\]\[1\] _01631_ _02420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_60_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09425__I1 net94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08389__A1 _03922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_76_1813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_170_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_79_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06156_ _01675_ _02349_ _02350_ _02351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_130_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10196__A1 _05078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09050__A2 _04339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_106_1050 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06087_ rf_ram.memory\[322\]\[1\] _01652_ _01654_ rf_ram.memory\[323\]\[1\] _01715_
+ rf_ram.memory\[321\]\[1\] _02282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XANTENNA__05611__A2 _01724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09915_ rf_ram.memory\[344\]\[1\] _04912_ _04914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09846_ _01452_ _04632_ _04871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__07364__A2 _02822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09777_ _04634_ _04828_ _04829_ _01141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_154_1313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06989_ rf_ram.memory\[227\]\[1\] _03051_ _03054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_38_1129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05913__B _01790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06795__I _02922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08728_ _04129_ _04149_ _04151_ _00770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_107_2378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08313__A1 _03230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07116__A2 _03135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_107_2389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08659_ _04094_ _04108_ _04109_ _00743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_124_2692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_174_clk clknet_5_31__leaf_clk clknet_leaf_174_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__10120__A1 _03008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05678__A2 _01649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06875__A1 _02970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11670_ net122 net194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_83_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_187_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_36_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10621_ _00365_ clknet_leaf_157_clk rf_ram.memory\[352\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_37_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_148_1106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_12_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_153_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10552_ _00296_ clknet_leaf_205_clk rf_ram.memory\[36\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_106_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_36_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_134_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06463__C _01568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05835__C1 _02019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_1258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10483_ _00227_ clknet_leaf_132_clk rf_ram.memory\[41\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_122_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07052__A1 _03087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11104_ _00840_ clknet_leaf_79_clk rf_ram.memory\[439\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_120_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05602__A2 _01709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_34_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_34_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_1182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_183_3785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11035_ _00772_ clknet_leaf_0_clk rf_ram.memory\[148\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_183_3796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08552__A1 _04026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_1207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_95_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_165_clk clknet_5_27__leaf_clk clknet_leaf_165_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_24_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06315__B1 _01848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08855__A2 _04195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_157_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_185_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_157_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_1251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10819_ _00563_ clknet_leaf_317_clk rf_ram.memory\[547\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_156_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09804__A1 _04837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_171_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_137_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09280__A2 _01341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_495 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_93_2124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_93_2135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06010_ rf_ram.memory\[542\]\[1\] _01532_ _01505_ _02205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09457__S _04604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05841__A2 _01915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput204 net204 o_ibus_adr[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_3_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput215 net215 o_ibus_adr[21] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_112_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput226 net226 o_ibus_adr[31] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_140_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_54_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09256__I _01356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08791__A1 _04170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_71_1721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07961_ _03654_ _03659_ _03661_ _00493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_160_Left_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09700_ _04740_ net3 _04777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_06912_ rf_ram.memory\[27\]\[1\] _03001_ _03003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07892_ _03590_ _03616_ _03618_ _00467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08543__A1 _04023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09631_ cpu.decode.opcode\[1\] net58 _04526_ _04724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06843_ _02927_ _02955_ _02956_ _00080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_136_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09562_ _04679_ _01076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05733__B _01928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06774_ rf_ram.memory\[512\]\[1\] _02905_ _02907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08513_ _04009_ _04015_ _04016_ _00690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06548__C _01341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05725_ _01917_ _01920_ _01790_ _01921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_19_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_69_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10102__A1 _05014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_1162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06306__B1 _01520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09493_ _01439_ _04625_ _04627_ _04628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_81_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_156_clk clknet_5_26__leaf_clk clknet_leaf_156_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_37_1184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08444_ _02945_ _03949_ _03964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05656_ rf_ram.memory\[465\]\[0\] _01787_ _01852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_136_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_102_2286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_102_2297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08375_ rf_ram.memory\[186\]\[0\] _03920_ _03921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_110_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05587_ _01550_ _01783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_45_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_985 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07326_ rf_ram.memory\[255\]\[1\] _03265_ _03267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_128_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05817__C1 _01931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06085__A2 _01709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07282__A1 _03222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07257_ _02894_ _03040_ _03223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_104_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_1003 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06208_ _01674_ _02391_ _02402_ net254 _02403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__05832__A2 _01940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10169__A1 _05046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07188_ _03161_ _03178_ _03180_ _00201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_143_1036 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07034__A1 _02779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06139_ _02322_ _02326_ _02330_ _02333_ _02334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_112_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_148_3135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_148_3146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08782__A1 net243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output156_I net156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_1199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_165_3460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_109_2418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_109_2429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09829_ _04837_ _04860_ _04861_ _01161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_126_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_126_2743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_161_3379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05643__B _01504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_1314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_185_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_147_clk clknet_5_26__leaf_clk clknet_leaf_147_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_55_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_1137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11653_ net103 net175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_126_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06474__B _01563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10604_ _00348_ clknet_leaf_152_clk rf_ram.memory\[356\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_119_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11584_ _01316_ clknet_leaf_30_clk rf_ram.memory\[212\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_91_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10535_ _00279_ clknet_leaf_140_clk rf_ram.memory\[265\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06076__A2 _01692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07273__A1 _03225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_843 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10466_ _00210_ clknet_leaf_138_clk rf_ram.memory\[261\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_165_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_0_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_185_3825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_185_3836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10397_ _00141_ clknet_leaf_214_clk rf_ram.memory\[245\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_20_565 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08525__A1 net248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07328__A2 _02954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11018_ _00755_ clknet_leaf_329_clk rf_ram.memory\[154\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06000__A2 _01538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_172_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_158_910 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_138_clk clknet_5_25__leaf_clk clknet_leaf_138_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__06839__A1 _02779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05510_ _01686_ _01706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_129_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06490_ _01349_ _02673_ _02684_ net254 _02685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_142_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_47_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_173_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05441_ rf_ram.memory\[364\]\[0\] _01634_ _01610_ rf_ram.memory\[365\]\[0\] _01636_
+ rf_ram.memory\[367\]\[0\] _01637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_0_142_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_64_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06384__B _01551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_173_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08160_ _03757_ _03784_ _03786_ _00567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_43_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05372_ _01347_ cpu.immdec.imm19_12_20\[5\] _01567_ _01568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XANTENNA__09253__A2 _01418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_7_clk_I clknet_5_0__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07111_ _03123_ _03131_ _03132_ _00172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_126_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08091_ rf_ram.memory\[558\]\[1\] _03742_ _03744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_310_clk clknet_5_5__leaf_clk clknet_leaf_310_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_125_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07042_ _02830_ _02939_ _03088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_30_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05814__A2 _01631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_1199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_113_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07016__A1 _03053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05728__B _01923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_321_clk_I clknet_5_5__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08764__A1 _04167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08993_ rf_ram.memory\[113\]\[0\] _04316_ _04317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07944_ _03622_ _03648_ _03650_ _00487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08516__A1 _03953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_143_3043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_173_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07875_ _03587_ _03607_ _03608_ _00460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_143_3054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_336_clk_I clknet_5_0__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_3_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05463__B _01658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06826_ _02930_ _02942_ _02944_ _00075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_3_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09614_ rf_ram.memory\[72\]\[0\] _04717_ _04718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_97_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_104_2326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_167_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09545_ _01595_ _04654_ _04666_ _01072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_78_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_104_2337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06757_ _02881_ _02894_ _02895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
Xclkbuf_leaf_129_clk clknet_5_13__leaf_clk clknet_leaf_129_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__05750__A1 _01350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_921 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_167_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_121_2640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_84_1956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_174_Right_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05708_ rf_ram.memory\[400\]\[0\] _01634_ _01903_ _01904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_84_1967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_121_2651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09476_ _04614_ _01055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_148_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06688_ rf_ram.memory\[525\]\[0\] _02847_ _02848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_148_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_149_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08427_ _03685_ _03953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_176_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05639_ _01527_ _01833_ _01834_ _01835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_108_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06294__B _01928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_175_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08358_ net235 _03903_ _03910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_188_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_163_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_61_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_149_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07255__A1 _03193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07309_ rf_ram.memory\[257\]\[1\] _03254_ _03256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_301_clk clknet_5_6__leaf_clk clknet_leaf_301_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08289_ rf_ram.memory\[192\]\[0\] _03866_ _03867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_34_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_1266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10320_ _00064_ clknet_leaf_211_clk rf_ram.memory\[510\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05805__A2 _01692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_1239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_167_3500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07007__A1 _02738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10251_ _02819_ _05119_ _05120_ _01325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08755__A1 _04167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10182_ _02742_ _05078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_121_1131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_163_3419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_1015 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_180_3733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_180_3744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_156_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09180__A1 _04431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_97_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_141_Right_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_69_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_178_3695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_166_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06297__A2 _01523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05820__C _01569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11636_ net86 net159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_108_840 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_139_2978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_142_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_42_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06049__A2 _01617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07246__A1 _02882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_154_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_42_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11567_ _01299_ clknet_leaf_24_clk rf_ram.memory\[190\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_52_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08994__A1 _04298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10518_ _00262_ clknet_leaf_211_clk rf_ram.memory\[26\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11498_ _01230_ clknet_leaf_185_clk rf_ram.memory\[504\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_150_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10449_ _00193_ clknet_leaf_186_clk rf_ram.memory\[483\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08746__A1 _04157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_1194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06221__A2 _01846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_1069 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05990_ _02102_ _02129_ _01372_ _02185_ _02186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XTAP_TAPCELL_ROW_88_2034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06379__B _02573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09171__A1 _04401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07660_ _03458_ _03472_ _03474_ _00379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_0_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_49_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_49_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_172_1040 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06611_ _02717_ _02718_ _02785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_07591_ rf_ram.memory\[355\]\[1\] _03430_ _03432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_149_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_66_1620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_177_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_66_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_172_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09330_ _04463_ _04533_ _04534_ _00989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_73_1170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06542_ _02727_ _02728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_62_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07485__A1 _03356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09261_ cpu.mem_bytecnt\[1\] _01385_ cpu.decode.co_ebreak _01460_ _04488_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_06473_ rf_ram.memory\[26\]\[1\] _01686_ _01624_ rf_ram.memory\[27\]\[1\] _02667_
+ _02668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_29_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08212_ rf_ram.memory\[535\]\[1\] _03817_ _03819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_146_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05424_ _01493_ _01620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_90_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09192_ rf_ram.memory\[83\]\[1\] _04439_ _04441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_56_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08143_ _03754_ _03775_ _03776_ _00560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_44_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05355_ _01550_ _01551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_70_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08074_ rf_ram.memory\[561\]\[0\] _03733_ _03734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05286_ _01468_ _01481_ _01483_ _01480_ _01484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_0_114_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_260_clk_I clknet_5_17__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_109_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07025_ rf_ram.memory\[218\]\[0\] _03076_ _03077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_140_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06460__A2 _01499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08737__A1 _01369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_1147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_1196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08976_ _04301_ _04304_ _04306_ _00863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_leaf_275_clk_I clknet_5_16__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input32_I i_dbus_rdt[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07927_ _03619_ _03639_ _03640_ _00480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_39_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09162__A1 net235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07858_ _02728_ _02869_ _03598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_168_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06809_ rf_ram.memory\[290\]\[0\] _02932_ _02933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_116_1211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07789_ _03039_ _03135_ _03555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA_output119_I net119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09528_ _04646_ _04650_ _04651_ _04655_ _01066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_112_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09459_ net79 net80 _04604_ _04606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06279__A2 _01523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_213_clk_I clknet_5_19__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_156_3289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07228__A1 _03190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11421_ _01153_ clknet_leaf_24_clk rf_ram.memory\[74\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_123_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_145_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08976__A1 _04301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11352_ _01084_ clknet_leaf_280_clk cpu.immdec.imm24_20\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_61_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_228_clk_I clknet_5_23__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_134_2886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_958 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10303_ _00047_ clknet_leaf_286_clk rf_ram.memory\[51\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_104_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11283_ _01018_ clknet_leaf_243_clk net219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06451__A2 _01530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08728__A1 _04129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10234_ _02737_ _02946_ _05110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06203__A2 _01724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07400__A1 _03292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10165_ rf_ram.memory\[448\]\[1\] _05066_ _05068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_22_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10096_ rf_ram.memory\[351\]\[0\] _05025_ _05026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_22_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09153__A1 _04397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06199__B _01650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_1105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_1198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10998_ _00735_ clknet_leaf_334_clk rf_ram.memory\[162\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_44_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_26_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_154_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11619_ net69 net141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_170_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_167_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_64_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08967__A1 _04298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05140_ cpu.decode.co_mem_word cpu.bne_or_bge _01342_ _01343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XANTENNA__06427__C1 _01679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_1148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_1125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xmax_cap236 _02922_ net236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_40_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xmax_cap247 _02774_ net247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_110_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08719__A1 _02983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09465__S _04604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_59_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08830_ net246 _02832_ _04216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08761_ _04172_ _04009_ _04173_ _00781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05973_ rf_ram.memory\[30\]\[0\] _01530_ _02169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_140_3002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07712_ _03488_ _03506_ _03507_ _00398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08692_ rf_ram.memory\[154\]\[1\] _04127_ _04130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_174_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_79_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07643_ _03455_ _03463_ _03464_ _00372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_36_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_71_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05741__B _01756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07574_ rf_ram.memory\[317\]\[1\] _03419_ _03421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_81_1904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09313_ _03992_ _04524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__07458__A1 _03326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06525_ _02712_ net97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_119_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05469__B1 _01664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_60_clk clknet_5_9__leaf_clk clknet_leaf_60_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09244_ cpu.genblk3.csr.timer_irq_r _04474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06456_ _02649_ _02650_ _01562_ _02651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_1_Left_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_7_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_134_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05407_ _01602_ _01603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_16_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09175_ rf_ram.memory\[85\]\[1\] _04428_ _04430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06387_ _02579_ _02581_ _01928_ _02582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_133_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_1301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_161_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08958__A1 _04269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08126_ _02829_ _03765_ _03766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05338_ _01507_ _01522_ _01529_ _01533_ _01534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_43_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_116_2550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_79_1866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_116_2561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_151_3197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_1_Right_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07630__A1 _02882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08057_ rf_ram.memory\[564\]\[0\] _03722_ _03723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_82_1258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05269_ _01363_ _01459_ _01463_ cpu.genblk3.csr.mstatus_mie _01467_ _01468_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_141_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07008_ rf_ram.memory\[223\]\[0\] _03065_ _03066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_101_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05641__B1 _01654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_112_2469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_991 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_94_clk_I clknet_5_14__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_157_1322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08959_ net246 _03945_ _04295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09135__A1 _04401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07697__A1 _03488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10921_ _00665_ clknet_leaf_206_clk rf_ram.memory\[29\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_98_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_158_3329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10852_ _00596_ clknet_leaf_308_clk rf_ram.memory\[530\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_6_1114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_5_12__f_clk_I clknet_3_3_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05172__A2 _01362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_152_clk_I clknet_5_26__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_175_3643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07449__A1 _02946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10783_ _00527_ clknet_leaf_326_clk rf_ram.memory\[565\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_17_1182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_1169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_51_clk clknet_5_12__leaf_clk clknet_leaf_51_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_186_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_81_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_66_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_32_clk_I clknet_5_6__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_136_2915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_136_2926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_151_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_167_clk_I clknet_5_30__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08949__A1 _02983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11404_ _01136_ clknet_leaf_231_clk net119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__05880__B1 _01912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_958 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_10_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_47_clk_I clknet_5_12__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07621__A1 _03422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_10_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11335_ _01067_ clknet_leaf_217_clk cpu.immdec.imm19_12_20\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_104_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06424__A2 _01641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11266_ _01001_ clknet_leaf_247_clk net232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_10217_ rf_ram.memory\[207\]\[1\] _05098_ _05100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05826__B _01551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_37_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11197_ _00933_ clknet_leaf_58_clk rf_ram.memory\[88\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_20_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_37_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10148_ rf_ram.memory\[451\]\[0\] _05057_ _05058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_59_1216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_19_Left_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_59_1238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_105_clk_I clknet_5_15__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09126__A1 _04397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10079_ _02814_ _02917_ _05015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07688__A1 _03491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_159_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_1141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05561__B _01756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_130_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_42_clk clknet_5_13__leaf_clk clknet_leaf_42_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_128_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06310_ _01552_ _02503_ _02504_ _02505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_127_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07290_ _02836_ _03135_ _03244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_183_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_155_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_28_Left_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_84_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06241_ rf_ram.memory\[432\]\[1\] _01782_ _01916_ _02436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_4_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07860__A1 _03587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_182_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06172_ rf_ram.memory\[504\]\[1\] _01755_ _01756_ _02367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_14_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_96_2177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_958 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_96_2188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07612__A1 _03425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05623__B1 _01793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09931_ _04918_ _04923_ _04924_ _01201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_1_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_111_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08168__A2 _02909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_74_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_1129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09862_ rf_ram.memory\[5\]\[0\] _04881_ _04882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_37_Left_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07915__A2 _02869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08813_ rf_ram.memory\[138\]\[1\] _04203_ _04206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05387__C1 _01554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09793_ _04837_ _04838_ _04839_ _01147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09117__A1 _02908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08744_ _04157_ _04162_ _00775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05956_ rf_ram.memory\[52\]\[0\] _01508_ _01655_ rf_ram.memory\[53\]\[0\] _01518_
+ rf_ram.memory\[55\]\[0\] _02152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_23_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07679__A1 _03455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08675_ rf_ram.memory\[156\]\[1\] _04117_ _04119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_68_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05887_ rf_ram.memory\[65\]\[0\] _01918_ _02083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_36_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05471__B _01526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07626_ _03422_ _03452_ _03453_ _00366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_177_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_138_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05154__A2 _01356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07557_ rf_ram.memory\[358\]\[0\] _03410_ _03411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_76_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_46_Left_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_leaf_33_clk clknet_5_6__leaf_clk clknet_leaf_33_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_06508_ _01412_ _01383_ _01423_ _01398_ _02698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_36_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_48_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07488_ _02795_ _02815_ _03368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_146_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_153_3237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09227_ rf_ram.memory\[339\]\[1\] _04460_ _04462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06439_ rf_ram.memory\[40\]\[1\] _01613_ _01601_ _02634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_173_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_170_3551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09158_ rf_ram.memory\[88\]\[0\] _04419_ _04420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_114_2509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_1000 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output186_I net186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_131_2823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08109_ net247 _03729_ _03755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_82_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_1018 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07603__A1 _02935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_146_1078 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_131_2834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09089_ _04364_ _04375_ _04376_ _00906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_82_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11120_ _00856_ clknet_leaf_86_clk rf_ram.memory\[120\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_31_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_55_Left_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_120_1218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11051_ _00788_ clknet_leaf_7_clk rf_ram.memory\[142\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_101_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07417__I _03013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10002_ rf_ram.memory\[504\]\[0\] _04967_ _04968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05378__C1 _01517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_129_2785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_129_2796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06590__A1 _02752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05393__A2 _01524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_28_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_1271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_153_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_1173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_58_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08331__A2 _02984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10904_ _00648_ clknet_leaf_20_clk rf_ram.memory\[186\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_39_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06342__A1 _01972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_64_Left_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_169_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_1179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10835_ _00579_ clknet_leaf_285_clk rf_ram.memory\[53\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_66_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_27_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_24_clk clknet_5_3__leaf_clk clknet_leaf_24_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_109_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08095__A1 _03721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10766_ _00510_ clknet_leaf_327_clk rf_ram.memory\[573\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_125_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_171_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_137_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07842__A1 _02953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10697_ _00441_ clknet_leaf_82_clk rf_ram.memory\[433\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_120_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_124_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_1129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_39_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_563 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_39_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_61_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_73_Left_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_188_3878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_188_3889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11318_ _01051_ clknet_leaf_263_clk net83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_91_2085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_91_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11249_ _00985_ clknet_leaf_279_clk cpu.immdec.imm11_7\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_4
XTAP_TAPCELL_ROW_52_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05810_ rf_ram.memory\[188\]\[0\] _01677_ _01793_ rf_ram.memory\[189\]\[0\] _01679_
+ rf_ram.memory\[191\]\[0\] _02006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_59_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06790_ _02873_ _02918_ _02919_ _00064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_89_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_166_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05741_ rf_ram.memory\[426\]\[0\] _01808_ _01756_ _01937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_171_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06387__B _01928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_82_Left_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_89_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08460_ net124 _03976_ _03977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_89_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_159_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_72_1246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05672_ rf_ram.memory\[460\]\[0\] _01709_ _01721_ rf_ram.memory\[461\]\[0\] _01713_
+ rf_ram.memory\[463\]\[0\] _01868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_07411_ _02814_ _03319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_187_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_174_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08391_ rf_ram.memory\[199\]\[0\] _03930_ _03931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_175_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05541__C1 _01678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_15_clk clknet_5_2__leaf_clk clknet_leaf_15_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_163_808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_161_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07342_ _03260_ _03274_ _03276_ _00259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_98_2217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_169_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_98_2228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09822__A2 _02984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07833__A1 _03554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07273_ _03225_ _03231_ _03233_ _00233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_112_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_147_1310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_115_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09012_ _02774_ _03945_ _04328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06224_ _02407_ _02411_ _02415_ _02418_ _02419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__05310__I _01505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_76_1803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_171_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_530 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_76_1814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09586__A1 net134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_91_Left_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_79_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06155_ rf_ram.memory\[492\]\[1\] _01677_ _01678_ rf_ram.memory\[493\]\[1\] _01679_
+ rf_ram.memory\[495\]\[1\] _02350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_112_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06086_ rf_ram.memory\[320\]\[1\] _01711_ _01602_ _02281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09338__A1 net65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09914_ _04884_ _04912_ _04913_ _01195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_42_1061 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08010__A1 _02959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09845_ _01413_ _03989_ _04870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_77_1102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_1108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09776_ rf_ram.memory\[77\]\[0\] _04828_ _04829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05375__A2 _01502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06988_ _03017_ _03053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_08727_ rf_ram.memory\[14\]\[1\] _04149_ _04151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05939_ rf_ram.memory\[42\]\[0\] _01605_ _01607_ rf_ram.memory\[43\]\[0\] _02134_
+ _02135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_68_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_107_2379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08313__A2 _02839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06324__A1 net251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08658_ rf_ram.memory\[15\]\[0\] _04108_ _04109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_178_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10120__A2 _03547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_124_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_1242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_178_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07609_ rf_ram.memory\[353\]\[0\] _03442_ _03443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_152_1071 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output101_I net101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08589_ _04058_ _04064_ _04065_ _00717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_95_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10620_ _00364_ clknet_leaf_158_clk rf_ram.memory\[352\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08077__A1 _03724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10551_ _00295_ clknet_leaf_165_clk rf_ram.memory\[332\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06627__A2 cpu.immdec.imm11_7\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_162_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_1226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05835__B1 _01968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_565 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10482_ _00226_ clknet_leaf_132_clk rf_ram.memory\[41\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_161_1318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_161_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11103_ _00839_ clknet_leaf_83_clk rf_ram.memory\[125\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_124_1173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_1270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11034_ _00771_ clknet_leaf_0_clk rf_ram.memory\[148\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_34_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08001__A1 _02761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_183_3786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_183_3797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_188_Right_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_21_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_1219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09501__A1 _03445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_157_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_1144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_184_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08068__A1 net236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_184_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10818_ _00562_ clknet_leaf_317_clk rf_ram.memory\[547\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_32_1263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_1039 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07815__A1 _03557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10749_ _00493_ clknet_leaf_186_clk rf_ram.memory\[480\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_54_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_530 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_93_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_152_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09568__A1 _03992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput205 net205 o_ibus_adr[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_26_1023 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput216 net216 o_ibus_adr[22] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput227 net227 o_ibus_adr[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_26_1034 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08240__A1 _03823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_54_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_1078 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_71_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_71_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07960_ rf_ram.memory\[480\]\[1\] _03659_ _03661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_4_clk clknet_5_1__leaf_clk clknet_leaf_4_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_103_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09473__S _04604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06911_ _02970_ _03001_ _03002_ _00102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_4_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07891_ rf_ram.memory\[445\]\[1\] _03616_ _03618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_155_Right_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09630_ _04643_ _01382_ _04723_ _01100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06842_ rf_ram.memory\[303\]\[0\] _02955_ _02956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06896__I _02991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05357__A2 _01511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06554__A1 _01369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09561_ cpu.immdec.imm30_25\[0\] _04675_ _04678_ _04679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06773_ _02873_ _02905_ _02906_ _00060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_136_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05724_ rf_ram.memory\[434\]\[0\] _01856_ _01911_ rf_ram.memory\[435\]\[0\] _01919_
+ _01920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_08512_ _01353_ rf_ram_if.wen0_r _04016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_19_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_19_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09492_ _01490_ _04626_ _04627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_69_1684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05305__I _01500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_1027 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08443_ _03956_ _03961_ _03963_ _00673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05655_ rf_ram.memory\[464\]\[0\] _01782_ _01693_ _01851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05514__C1 _01654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08374_ net245 _03903_ _03920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_102_2287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_175_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_493 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_102_2298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05586_ _01682_ _01782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_73_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07325_ _03257_ _03265_ _03266_ _00252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07806__A1 _02916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_5_18__f_clk clknet_3_4_0_clk clknet_5_18__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_46_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05817__B1 _01911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07256_ _03013_ _03222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_147_1140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09559__A1 _01491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06207_ _01350_ _02396_ _02401_ _02402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_42_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_143_1015 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07187_ rf_ram.memory\[198\]\[1\] _03178_ _03180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_41_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input62_I i_ibus_rdt[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06138_ _01675_ _02331_ _02332_ _02333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_41_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08231__A1 _03798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_148_3136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08782__A2 _04152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_148_3147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06069_ rf_ram.memory\[350\]\[1\] _01543_ _02264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_100_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05596__A2 _01735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_165_3450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_165_3461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_109_2419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09828_ rf_ram.memory\[62\]\[0\] _04860_ _04861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05924__B _01783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_122_Right_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06545__A1 cpu.immdec.imm11_7\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_126_2733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_126_2744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_158_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09759_ net118 _04766_ _04760_ net119 _04817_ _04818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_0_119_1242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08298__A1 _03309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_1252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_1128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_167_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_167_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11652_ net102 net174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05520__A2 _01652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_182_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_166_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10603_ _00347_ clknet_leaf_154_clk rf_ram.memory\[317\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_36_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11583_ _01315_ clknet_leaf_30_clk rf_ram.memory\[212\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_107_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10534_ _00278_ clknet_leaf_140_clk rf_ram.memory\[265\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_122_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_1202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_10_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_165_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_134_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10465_ _00209_ clknet_leaf_196_clk rf_ram.memory\[262\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_122_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_185_3826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10396_ _00140_ clknet_leaf_214_clk rf_ram.memory\[245\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_185_3837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05818__C _01978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06784__A1 _02876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08525__A2 _02869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09722__A1 net105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11017_ _00754_ clknet_leaf_332_clk rf_ram.memory\[155\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05339__A2 _01502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_59_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_47_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_157_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_47_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05440_ _01635_ _01636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_74_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_185_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_145_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_64_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_64_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_172_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09789__A1 _04637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_51_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05371_ _01355_ _01360_ _01567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_71_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_166_1026 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_923 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07110_ rf_ram.memory\[488\]\[0\] _03131_ _03132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_55_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08090_ _03721_ _03742_ _03743_ _00540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_126_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_1313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07041_ _03013_ _03087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_140_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08213__A1 _03790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10020__A1 _04953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09961__A1 _04918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08992_ net248 _04303_ _04316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05578__A2 _01711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06775__A1 _02876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_177_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07943_ rf_ram.memory\[43\]\[1\] _03648_ _03650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_10_Left_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_76_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05983__C1 _01635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09713__A1 _04781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_143_3044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07874_ rf_ram.memory\[463\]\[0\] _03607_ _03608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_143_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09613_ net250 _04507_ _04717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06825_ rf_ram.memory\[287\]\[1\] _02942_ _02944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_39_1247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_104_2327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09544_ _04478_ net42 _04650_ cpu.immdec.imm19_12_20\[6\] _04666_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_TAPCELL_ROW_104_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06756_ _02893_ _02894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_66_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10087__A1 _05014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_121_2641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_84_1957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05707_ _01525_ _01903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_121_2652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09475_ net88 net89 _04604_ _04614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06687_ _02844_ _02846_ _02847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_66_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_84_1968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08426_ _03922_ _03950_ _03952_ _00667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_136_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05638_ rf_ram.memory\[508\]\[0\] _01644_ _01610_ rf_ram.memory\[509\]\[0\] _01636_
+ rf_ram.memory\[511\]\[0\] _01834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XANTENNA__05502__A2 _01697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_136_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08357_ _03887_ _03907_ _03909_ _00641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05569_ _01760_ _01761_ _01762_ _01764_ _01670_ _01765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_135_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_1069 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_1212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07308_ _03222_ _03254_ _03255_ _00246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_150_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08452__A1 _01369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08288_ _03230_ _02904_ _03866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_22_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_1199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_132_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05266__A1 _01409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07239_ rf_ram.memory\[422\]\[1\] _03210_ _03212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_116_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_167_3501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10250_ rf_ram.memory\[28\]\[0\] _05119_ _05120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_132_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08204__A1 _03798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07007__A2 _02909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06215__B1 _01778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10011__A1 _04911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10181_ _05049_ _05075_ _05077_ _01298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06766__A1 _02873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05974__C1 _01607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_180_3734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_180_3745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09704__B2 net101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07191__A1 _03157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05741__A2 _01808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_1156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_178_3696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_167_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_1077 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11635_ net85 net158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_53_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_139_2979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_154_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07246__A2 _03040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_42_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08443__A1 _03956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_181_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_42_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11566_ _01298_ clknet_leaf_36_clk rf_ram.memory\[202\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_108_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10517_ _00261_ clknet_leaf_218_clk rf_ram.memory\[253\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_126_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05829__B _01978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11497_ _01229_ clknet_leaf_186_clk rf_ram.memory\[504\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10448_ _00192_ clknet_leaf_197_clk rf_ram.memory\[483\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_122_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_1053 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09943__A1 _04921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10379_ _00123_ clknet_leaf_99_clk rf_ram.memory\[428\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06757__A1 _02881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05564__B _01504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_88_2035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05980__A2 _01643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06379__C _01569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05717__C1 _01912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_49_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_49_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06610_ _02748_ _02782_ _02784_ _00019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07590_ _03422_ _03430_ _03431_ _00352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_88_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_66_1621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_149_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_66_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_177_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06541_ _02716_ _02726_ _02727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_87_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_146_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09260_ cpu.state.cnt_r\[3\] cpu.state.o_cnt\[2\] _04487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06472_ rf_ram.memory\[25\]\[1\] _01514_ _02667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__08682__A1 _02821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_146_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05423_ rf_ram.memory\[354\]\[0\] _01606_ _01608_ rf_ram.memory\[355\]\[0\] _01618_
+ _01619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_29_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08211_ _03787_ _03817_ _03818_ _00586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_157_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09191_ _04431_ _04439_ _04440_ _00944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_28_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_173_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_7_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_173_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08142_ rf_ram.memory\[548\]\[0\] _03775_ _03776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_16_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05354_ _01525_ _01550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_132_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08434__A1 _02971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10241__A1 _02819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06445__B1 _01607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08073_ _02761_ _03729_ _03733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_295_clk clknet_5_7__leaf_clk clknet_leaf_295_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__05739__B _01805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05285_ _01405_ _01482_ _01483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06996__A1 _03053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07024_ _02738_ _02813_ _03076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_114_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_144_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_1165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05263__A4 _01461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_1127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09934__A1 _04911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08737__A2 _04157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06748__A1 _02779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05956__C1 _01518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08975_ rf_ram.memory\[117\]\[1\] _04304_ _04306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07926_ rf_ram.memory\[458\]\[0\] _03639_ _03640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input25_I i_dbus_rdt[30] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_1000 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05971__A2 _01686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09162__A2 _04418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07857_ _03590_ _03595_ _03597_ _00453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07173__A1 _03161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_1093 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06808_ _02801_ _02894_ _02932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_39_1066 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_1223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07788_ _03355_ _03554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__05723__A2 _01918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06920__A1 _02773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09527_ cpu.immdec.imm19_12_20\[1\] _04654_ _04655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05921__C _01660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06739_ _02845_ _02881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_38_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_1206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09458_ _04605_ _01046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_164_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08409_ _03922_ _03939_ _03941_ _00661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_35_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09389_ _04567_ _01015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_149_1032 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11420_ _01152_ clknet_leaf_24_clk rf_ram.memory\[75\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_117_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_163_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05239__A1 _01434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_915 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_117_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_286_clk clknet_5_18__leaf_clk clknet_leaf_286_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_149_1098 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11351_ _01083_ clknet_leaf_258_clk cpu.immdec.imm24_20\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_162_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06987__A1 _03050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_134_2876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_134_2887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10302_ _00046_ clknet_leaf_286_clk rf_ram.memory\[51\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_131_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11282_ _01017_ clknet_leaf_244_clk net218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_104_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09925__A1 _04918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10233_ _05081_ _05107_ _05109_ _01318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_30_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10164_ _05046_ _05066_ _05067_ _01291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_7_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10095_ _02814_ _02909_ _05025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_156_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05962__A2 _01536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09571__S _03967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_6_clk_I clknet_5_2__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07164__A1 _02889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_639 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_210_clk clknet_5_25__leaf_clk clknet_leaf_210_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08900__A2 _04257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05714__A2 _01510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06911__A1 _02970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_69_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10997_ _00734_ clknet_leaf_308_clk rf_ram.memory\[549\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_96_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_44_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_320_clk_I clknet_5_5__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_44_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08664__A1 _04094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_26_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_26_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_61_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_155_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_182_563 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_155_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11618_ net68 net140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08416__A1 _02959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_277_clk clknet_5_16__leaf_clk clknet_leaf_277_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__10223__A1 _05081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06427__B1 _01793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11549_ _01281_ clknet_leaf_122_clk rf_ram.memory\[453\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06978__A1 _03018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_180_1321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xmax_cap237 _02903_ net237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_64_1148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_151_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05278__C _01366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xmax_cap248 _02760_ net248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__09916__A1 _04887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08719__A2 _04005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_59_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05402__A1 _01347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08760_ _01353_ rf_ram_if.wen1_r _04173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05972_ _02165_ _02167_ _01563_ _02168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05953__A2 _01661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09481__S _01411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_140_3003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07711_ rf_ram.memory\[3\]\[0\] _03506_ _03507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08691_ _04061_ _04129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_79_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07155__A1 _03157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_201_clk clknet_5_25__leaf_clk clknet_leaf_201_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07642_ rf_ram.memory\[387\]\[0\] _03463_ _03464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_75_1266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_178_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05705__A2 _01623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06902__A1 _02867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07573_ _03389_ _03419_ _03420_ _00346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_177_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_81_1905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_165_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09312_ _04520_ _04521_ _04522_ _02721_ _04523_ _00982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_06524_ cpu.state.init_done _02709_ _02710_ _02711_ _02712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_75_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05313__I _01508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_146_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_958 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09243_ _04471_ _04472_ _04473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_29_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06455_ rf_ram.memory\[58\]\[1\] _01661_ _01653_ rf_ram.memory\[59\]\[1\] _01655_
+ rf_ram.memory\[57\]\[1\] _02650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_28_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06130__A2 _01777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08407__A1 _03919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05406_ _01601_ _01602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_113_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06386_ rf_ram.memory\[74\]\[1\] _01808_ _01925_ rf_ram.memory\[75\]\[1\] _02580_
+ _02581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_09174_ _04397_ _04428_ _04429_ _00938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_43_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_146_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06418__B1 _01911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_915 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_268_clk clknet_5_16__leaf_clk clknet_leaf_268_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__10214__A1 _03892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08125_ _03692_ _03765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_05337_ rf_ram.memory\[522\]\[0\] _01532_ _01521_ rf_ram.memory\[523\]\[0\] _01517_
+ rf_ram.memory\[521\]\[0\] _01533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_31_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_116_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06969__A1 _02788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_79_1867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_160_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_151_3198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08056_ _03134_ _03693_ _03722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05268_ _01465_ _01466_ _01467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07630__A2 _03089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07007_ _02738_ _02909_ _03065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_12_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05199_ cpu.decode.opcode\[2\] _01399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_45_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07394__A1 _03292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06197__A2 _01719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08958_ _04269_ _04292_ _04294_ _00857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_102_Left_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_99_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07909_ _03622_ _03627_ _03629_ _00473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_118_1307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08889_ _04234_ _04251_ _04252_ _00830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07146__A1 _02761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10920_ _00664_ clknet_leaf_207_clk rf_ram.memory\[29\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08894__A1 _04234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06354__C1 _01959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_155_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10851_ _00595_ clknet_leaf_310_clk rf_ram.memory\[531\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_39_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_175_3644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07449__A2 _03101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08646__A1 _04097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10782_ _00526_ clknet_leaf_326_clk rf_ram.memory\[565\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_93_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_136_2916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06121__A2 _01500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_136_2927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_34_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09446__I0 net73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08949__A2 _04038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_259_clk clknet_5_17__leaf_clk clknet_leaf_259_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_34_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11403_ _01135_ clknet_leaf_231_clk net118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__09071__A1 net248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09566__S _04678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_10_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11334_ _01066_ clknet_leaf_216_clk cpu.immdec.imm19_12_20\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_50_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_162_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11265_ _01000_ clknet_leaf_247_clk net231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_123_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10216_ _05078_ _05098_ _05099_ _01311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_98_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11196_ _00932_ clknet_leaf_58_clk rf_ram.memory\[88\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_37_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_1176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07385__A1 _02992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_37_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10147_ _03672_ _02889_ _05057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_118_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_1228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05935__A2 _01633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10078_ _04396_ _05014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__07613__I _02800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_806 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06360__A2 _01846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_57_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_0_clk clk clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__06112__A2 _01631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06240_ _01909_ _02433_ _02434_ _02435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_26_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_274_clk_I clknet_5_16__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_991 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_115_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_131_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06171_ _01527_ _02364_ _02365_ _02366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__09062__A1 _04331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_96_2178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_96_2189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_1054 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_180_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_leaf_289_clk_I clknet_5_18__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09930_ rf_ram.memory\[341\]\[0\] _04923_ _04924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_159_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_15_Right_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_74_1775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09861_ _02794_ _03035_ _04881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_111_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08812_ _04061_ _04205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA_clkbuf_leaf_212_clk_I clknet_5_19__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05387__B1 _01555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09792_ rf_ram.memory\[80\]\[0\] _04838_ _04839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_139_1020 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05308__I _01503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09117__A2 _03692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08743_ _04160_ _04161_ _04162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05955_ rf_ram.memory\[54\]\[0\] _01661_ _01503_ _02151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07128__A1 _03123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08674_ _04094_ _04117_ _04118_ _00749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08876__A1 _04237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05886_ rf_ram.memory\[64\]\[0\] _01537_ _01551_ _02082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_178_633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07523__I _03355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_leaf_227_clk_I clknet_5_23__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07625_ rf_ram.memory\[407\]\[0\] _03452_ _03453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_24_Right_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_89_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_5_4__f_clk_I clknet_3_1_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07556_ _02806_ _03390_ _03410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_159_880 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_159_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_76_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_165_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06507_ cpu.ctrl.pc_plus_offset_cy_r _01397_ _02697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07487_ _03360_ _03365_ _03367_ _00313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_63_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_107_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07300__A1 net239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_153_3238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09226_ _04431_ _04460_ _04461_ _00958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_1_1034 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_91_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06438_ _01903_ _02631_ _02632_ _02633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_146_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_170_3552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_146_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_1024 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09157_ _02991_ _04418_ _04419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_32_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06369_ rf_ram.memory\[244\]\[1\] _01634_ _01610_ rf_ram.memory\[245\]\[1\] _01636_
+ rf_ram.memory\[247\]\[1\] _02564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_44_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08108_ _03685_ _03754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_121_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_131_2824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07603__A2 _02813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_131_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09088_ rf_ram.memory\[569\]\[0\] _04375_ _04376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08800__A1 _04167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_169_Right_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_33_Right_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_output179_I net179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_1176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08039_ _03690_ _03709_ _03711_ _00521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05927__B _02004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11050_ _00787_ clknet_leaf_10_clk rf_ram.memory\[143\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_101_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10001_ _02910_ _02992_ _04967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05378__B1 _01521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_129_2786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_129_2797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06590__A2 _02766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_1115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_157_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08867__A1 net239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_28_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_42_Right_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_54_1114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10903_ _00647_ clknet_leaf_17_clk rf_ram.memory\[185\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_58_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_1267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_157_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08619__A1 _04062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10834_ _00578_ clknet_leaf_286_clk rf_ram.memory\[53\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09292__A1 _04466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10765_ _00509_ clknet_leaf_127_clk rf_ram.memory\[465\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_27_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06493__B _02687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07842__A2 _03234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09419__I0 net90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10696_ _00440_ clknet_leaf_82_clk rf_ram.memory\[433\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_81_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05853__A1 _01951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_1210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09044__A1 _04334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_51_Right_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_50_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_164_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_65_1243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_136_Right_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_39_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_121_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_39_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_188_3879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11317_ _01050_ clknet_leaf_262_clk net82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_120_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_56_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_91_2086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11248_ _00984_ clknet_leaf_280_clk cpu.immdec.imm11_7\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_91_2097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07358__A1 _02788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11179_ _00915_ clknet_leaf_55_clk rf_ram.memory\[94\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05908__A2 _01706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_52_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_1074 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_1185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_60_Right_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05740_ rf_ram.memory\[428\]\[0\] _01724_ _01725_ rf_ram.memory\[429\]\[0\] _01811_
+ rf_ram.memory\[431\]\[0\] _01936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_188_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06318__C1 _01773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_159_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05671_ rf_ram.memory\[462\]\[0\] _01808_ _01707_ _01867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07530__A1 _03393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06333__A2 _01515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07410_ _03292_ _03316_ _03318_ _00285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08390_ _03892_ _02829_ _03930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05541__B1 _01679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_159_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07341_ rf_ram.memory\[270\]\[1\] _03274_ _03276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_98_2218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_162_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_156_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_155_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_14_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07272_ rf_ram.memory\[193\]\[1\] _03231_ _03233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_171_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_93_clk_I clknet_5_14__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_5_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_115_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_1322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09011_ _04301_ _04325_ _04327_ _00877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06223_ _01675_ _02416_ _02417_ _02418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_14_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_60_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_72_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09035__A1 net249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_76_1804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_76_1815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06154_ rf_ram.memory\[494\]\[1\] _01543_ _02349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07597__A1 _03425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_103_Right_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05747__B _01756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06085_ rf_ram.memory\[324\]\[1\] _01709_ _01656_ rf_ram.memory\[325\]\[1\] _01654_
+ rf_ram.memory\[327\]\[1\] _02280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_106_1063 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09913_ rf_ram.memory\[344\]\[0\] _04912_ _04913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_10_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_151_clk_I clknet_5_26__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09844_ _02714_ _04869_ _01168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_176_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08010__A2 _03693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_31_clk_I clknet_5_6__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09775_ net243 _04507_ _04828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06987_ _03050_ _03051_ _03052_ _00128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08726_ _04126_ _04149_ _04150_ _00769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06309__C1 _01953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08849__A1 _04205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05938_ rf_ram.memory\[41\]\[0\] _01513_ _02134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_178_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08657_ _02953_ _03945_ _04108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_68_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05869_ rf_ram.memory\[242\]\[0\] _01606_ _01625_ rf_ram.memory\[243\]\[0\] _01702_
+ rf_ram.memory\[241\]\[0\] _02065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XANTENNA_clkbuf_leaf_46_clk_I clknet_5_12__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_124_2694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_113_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07608_ _02898_ _03390_ _03442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_117_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08588_ rf_ram.memory\[167\]\[0\] _04064_ _04065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_64_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07539_ rf_ram.memory\[360\]\[1\] _03398_ _03400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_36_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_181_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_10_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_12_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10550_ _00294_ clknet_leaf_165_clk rf_ram.memory\[332\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_146_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06627__A3 _02730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_736 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05501__I _01514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09209_ net241 _04418_ _04451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_104_clk_I clknet_5_15__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_1238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09026__A1 _04331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10481_ _00225_ clknet_leaf_104_clk rf_ram.memory\[420\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_161_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_32_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08812__I _04061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07588__A1 _02889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11102_ _00838_ clknet_leaf_83_clk rf_ram.memory\[125\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_119_clk_I clknet_5_12__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_34_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11033_ _00770_ clknet_leaf_294_clk rf_ram.memory\[14\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_120_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_34_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08001__A2 _02832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_183_3787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_183_3798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09501__A2 _02899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07512__A1 _03360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06315__A2 _01711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_185_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_86_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_169_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_129_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_157_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_1231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_995 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_1156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10817_ _00561_ clknet_leaf_319_clk rf_ram.memory\[548\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_67_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08068__A2 _03729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_172_639 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10748_ _00492_ clknet_leaf_197_clk rf_ram.memory\[480\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_165_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05411__I _01518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10679_ _00423_ clknet_leaf_110_clk rf_ram.memory\[374\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_140_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_93_2126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07579__A1 _03422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput206 net206 o_ibus_adr[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_11_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput217 net217 o_ibus_adr[23] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_112_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput228 net228 o_ibus_adr[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_54_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06251__A1 _01909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_71_1712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_71_1723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06910_ rf_ram.memory\[27\]\[0\] _03001_ _03002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07890_ _03587_ _03616_ _03617_ _00466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_156_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06841_ _02935_ _02954_ _02955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09740__A2 net16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07751__A1 _03524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09560_ _04477_ _04677_ _04678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_06772_ rf_ram.memory\[512\]\[0\] _02905_ _02906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08511_ _03989_ _04014_ _01366_ _04015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05723_ rf_ram.memory\[433\]\[0\] _01918_ _01919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_136_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_77_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_188_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_19_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09491_ cpu.alu.i_rs1 _04625_ _04626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_69_1674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07503__A1 _02781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06306__A2 _01989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_69_1685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08442_ rf_ram.memory\[175\]\[1\] _03961_ _03963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_72_1066 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05514__B1 _01656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05654_ _01769_ _01847_ _01849_ _01850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_187_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_65_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_176_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08373_ _03685_ _03919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_102_2288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_175_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05585_ _01776_ _01780_ _01746_ _01781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_102_2299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_163_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07324_ rf_ram.memory\[255\]\[0\] _03265_ _03266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_156_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07806__A2 _03559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05321__I _01516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07255_ _03193_ _03219_ _03221_ _00227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_171_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06206_ _02397_ _02398_ _02399_ _02400_ _01717_ _02401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__06490__A1 _01349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_171_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_170_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07186_ _03157_ _03178_ _03179_ _00200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_42_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_1136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_131_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05477__B _01672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06137_ rf_ram.memory\[294\]\[1\] _01777_ _01778_ rf_ram.memory\[295\]\[1\] _01793_
+ rf_ram.memory\[293\]\[1\] _02332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_0_14_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08231__A2 _02866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input55_I i_ibus_rdt[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_148_3137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06068_ _01600_ _02250_ _02262_ net253 _02263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XTAP_TAPCELL_ROW_148_3148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_165_3451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_165_3462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09827_ _03668_ _02917_ _04860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07742__A1 _02788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_126_2734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_126_2745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09758_ _04804_ net22 _04817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_08709_ net235 _04078_ _04140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_55_1242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08298__A2 _03135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09689_ net126 _04767_ _04768_ net127 _04769_ _04770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_0_68_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05940__B _01563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11651_ net101 net173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__09247__A1 _03967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10602_ _00346_ clknet_leaf_154_clk rf_ram.memory\[317\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_107_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_92_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11582_ _01314_ clknet_leaf_290_clk rf_ram.memory\[23\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_135_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_458 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_1073 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10533_ _00277_ clknet_leaf_209_clk rf_ram.memory\[24\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_49_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_134_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_load_slew245_I _02812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06481__A1 rf_ram.memory\[10\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_845 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10464_ _00208_ clknet_leaf_196_clk rf_ram.memory\[262\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_161_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06490__C net254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_185_3827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10395_ _00139_ clknet_leaf_295_clk rf_ram.memory\[222\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09574__S _03967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_1208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05441__C1 _01636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07981__A1 _03651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11016_ _00753_ clknet_leaf_332_clk rf_ram.memory\[155\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_137_1310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_5_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_5_24__f_clk clknet_3_6_0_clk clknet_5_24__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__05406__I _01601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_1099 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09486__A1 _01375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_87_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_16_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_185_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_157_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_47_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_47_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_184_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09238__A1 _04463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_954 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_185_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_64_1582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_64_1593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_166_1005 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05370_ _01557_ _01565_ _01351_ _01566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_28_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_1124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07040_ _03053_ _03084_ _03086_ _00147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_125_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_113_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08991_ _04301_ _04313_ _04315_ _00869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_167_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07942_ _03619_ _03648_ _03649_ _00486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05983__B1 _01714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_1220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_1231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09713__A2 net7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_1107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07873_ _02836_ _02954_ _03607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07724__A1 _03491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_143_3045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_143_3056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09612_ _04637_ _04714_ _04716_ _01089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06824_ _02927_ _02942_ _02943_ _00074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_97_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05316__I _01496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_160_3370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09543_ _01732_ _04654_ _04665_ _01071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_78_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06755_ _02773_ _02887_ _02893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XTAP_TAPCELL_ROW_104_2328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_151_1318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_149_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09477__A1 _02703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_104_2339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05706_ rf_ram.memory\[404\]\[0\] _01509_ _01656_ rf_ram.memory\[405\]\[0\] _01763_
+ rf_ram.memory\[407\]\[0\] _01902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_149_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_188_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_148_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09474_ _04613_ _01054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_84_1958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_121_2642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_148_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06686_ _02845_ _02846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_66_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_84_1969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_121_2653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_176_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08425_ rf_ram.memory\[173\]\[1\] _03950_ _03952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_65_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05637_ rf_ram.memory\[510\]\[0\] _01631_ _01833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_4_1235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_1101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_1026 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08356_ rf_ram.memory\[182\]\[1\] _03907_ _03909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_135_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_129_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05568_ rf_ram.memory\[258\]\[0\] _01500_ _01763_ rf_ram.memory\[259\]\[0\] _01668_
+ rf_ram.memory\[257\]\[0\] _01764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_18_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07307_ rf_ram.memory\[257\]\[0\] _03254_ _03255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_116_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08287_ _03855_ _03863_ _03865_ _00615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_117_875 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08452__A2 _01496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05499_ _01518_ _01695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_33_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06463__A1 _01599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07238_ _03190_ _03210_ _03211_ _00220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_132_845 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_1219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_167_3502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08204__A2 _02992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07169_ _02915_ _02954_ _03169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10011__A2 _02839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10180_ rf_ram.memory\[202\]\[1\] _05075_ _05077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_121_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09407__B _01344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05974__B1 _01617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_180_3735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08507__A3 cpu.immdec.imm11_7\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07715__A1 _02839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_1146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_139_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08140__A1 _03757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_178_3697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_127_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_182_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_139_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11634_ net84 net157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_53_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_139_2969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_154_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_42_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11565_ _01297_ clknet_leaf_36_clk rf_ram.memory\[202\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_25_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10516_ _00260_ clknet_leaf_219_clk rf_ram.memory\[253\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_21_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11496_ _01228_ clknet_leaf_189_clk rf_ram.memory\[276\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_52_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_150_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10447_ _00191_ clknet_leaf_198_clk rf_ram.memory\[496\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_150_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_139_Left_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10378_ _00122_ clknet_leaf_99_clk rf_ram.memory\[428\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_27_1185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06757__A2 _02894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07954__A1 _03651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_1217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_88_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_88_2036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05717__B1 _01911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_49_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_49_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06390__B1 _02019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_148_Left_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_137_1184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_66_1622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05580__B _01693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06540_ _02719_ _02725_ _02726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XTAP_TAPCELL_ROW_66_1633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_1281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_1172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08131__A1 _02805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_1183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_158_775 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06471_ rf_ram.memory\[24\]\[1\] _01682_ _01550_ _02666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08682__A2 _04078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08210_ rf_ram.memory\[535\]\[0\] _03817_ _03818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05422_ rf_ram.memory\[353\]\[0\] _01617_ _01618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_09190_ rf_ram.memory\[83\]\[0\] _04439_ _04440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_161_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08141_ net241 _03765_ _03775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05353_ rf_ram.memory\[532\]\[0\] _01523_ _01516_ rf_ram.memory\[533\]\[0\] _01520_
+ rf_ram.memory\[535\]\[0\] _01549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_83_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08434__A2 _03949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08072_ _03724_ _03730_ _03732_ _00533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05284_ _01442_ cpu.bne_or_bge _01482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_114_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_157_Left_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_148_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07023_ _03053_ _03073_ _03075_ _00141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05653__C1 _01848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_141_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08198__A1 _03790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09934__A2 _03135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08974_ _04298_ _04304_ _04305_ _00862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05956__B1 _01655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_162_3410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_89_Right_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05420__A2 _01614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07925_ _02774_ _02832_ _03639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09698__A1 net129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09698__B2 net99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07856_ rf_ram.memory\[430\]\[1\] _03595_ _03597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_166_Left_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08370__A1 _03884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06807_ _02930_ _02928_ _02931_ _00069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input18_I i_dbus_rdt[24] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07787_ _03524_ _03551_ _03553_ _00427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_155_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09526_ _03967_ _04653_ _04654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_06738_ _02876_ _02878_ _02880_ _00051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_94_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08122__A1 _03754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09457_ net78 net79 _04604_ _04605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_176_561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06669_ _02829_ _02832_ _02833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_176_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08408_ rf_ram.memory\[178\]\[1\] _03939_ _03941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_98_Right_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_164_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09388_ net216 _04561_ _04564_ net217 _04567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_19_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08339_ rf_ram.memory\[240\]\[1\] _03896_ _03898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_85_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09473__I1 net88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_175_Left_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_123_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_151_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11350_ _01082_ clknet_leaf_216_clk cpu.immdec.imm24_20\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__06605__I _02780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_1005 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05649__C net253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_134_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10301_ _00045_ clknet_leaf_316_clk rf_ram.memory\[520\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_43_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05644__C1 _01519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_134_2888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_132_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11281_ _01016_ clknet_leaf_244_clk net217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08189__A1 _03668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09386__B1 _04564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10232_ rf_ram.memory\[237\]\[1\] _05107_ _05109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_131_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_7_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10163_ rf_ram.memory\[448\]\[0\] _05066_ _05067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05665__B _01860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10094_ _05017_ _05022_ _05024_ _01264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05384__C _01495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09689__A1 net126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_184_Left_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_156_1037 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07164__A2 _03158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05175__A1 _01375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_1058 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10996_ _00733_ clknet_leaf_324_clk rf_ram.memory\[549\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_57_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_139_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_44_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_128_915 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_44_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09861__A1 _02794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_26_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_61_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_61_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_167_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11617_ net67 net139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_65_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09613__A1 net250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08416__A2 _03945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_182_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_170_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11548_ _01280_ clknet_leaf_121_clk rf_ram.memory\[454\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_107_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11479_ _01211_ clknet_leaf_177_clk rf_ram.memory\[336\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xmax_cap238 _02898_ net238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_122_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_110_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_150_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_59_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07927__A1 _03619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06060__C1 _01656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05402__A2 _01478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05971_ rf_ram.memory\[26\]\[0\] _01686_ _01624_ rf_ram.memory\[27\]\[0\] _02166_
+ _02167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_07710_ net240 _02997_ _03506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_140_3004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08690_ _04126_ _04127_ _04128_ _00755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_164_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08352__A1 _03887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07641_ _02889_ _03089_ _03463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_178_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06902__A2 _02939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07572_ rf_ram.memory\[317\]\[0\] _03419_ _03420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_81_1906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09311_ _04477_ net62 _04523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_88_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06523_ _01399_ _01381_ _02711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09852__A1 _01385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_1170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_76_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05469__A2 _01509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09242_ cpu.genblk3.csr.mie_mtie cpu.genblk3.csr.mstatus_mie net66 _04472_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__06666__A1 cpu.immdec.imm11_7\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_425 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_146_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06454_ rf_ram.memory\[56\]\[1\] _01613_ _01601_ _02649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_8_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05405_ rf_ram.i_raddr\[2\] _01601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__05874__C1 _01696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_1176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09173_ rf_ram.memory\[85\]\[0\] _04428_ _04429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_155_3280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09604__A1 _04478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06385_ rf_ram.memory\[73\]\[1\] _01918_ _02580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_133_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_1284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08124_ _03757_ _03762_ _03764_ _00553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05336_ _01531_ _01532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_71_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10214__A2 _02954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06969__A2 _03040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_79_1868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_116_2552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_151_3199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08055_ _03685_ _03721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__07091__A1 _03092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05267_ cpu.genblk3.csr.mcause31 _01418_ _01386_ cpu.genblk3.csr.mcause3_0\[0\] _01466_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_98_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_141_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07006_ _03053_ _03062_ _03064_ _00135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_141_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05641__A2 _01652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05198_ cpu.ctrl.pc_plus_offset_cy_r _01397_ _01398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_101_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07256__I _03013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08591__A1 _04062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08957_ rf_ram.memory\[120\]\[1\] _04292_ _04294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07908_ rf_ram.memory\[460\]\[1\] _03627_ _03629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08888_ rf_ram.memory\[479\]\[0\] _04251_ _04252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08343__A1 _03884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07146__A2 _02911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07839_ rf_ram.memory\[411\]\[1\] _03584_ _03586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06354__B1 _01968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10850_ _00594_ clknet_leaf_306_clk rf_ram.memory\[531\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_67_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09509_ _04634_ _04639_ _04640_ _01062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06106__B1 _01679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10781_ _00525_ clknet_leaf_325_clk rf_ram.memory\[566\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_13_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_177_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_175_3645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06657__A1 _02815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_87_1105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_117_Right_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_136_2917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_136_2928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09446__I1 net74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11402_ _01134_ clknet_leaf_230_clk net117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_136_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05880__A2 _01755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09071__A2 _04005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11333_ _01065_ clknet_leaf_236_clk cpu.immdec.imm31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07082__A1 _02781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_5_21__f_clk_I clknet_3_5_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06290__C1 _01857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11264_ _00999_ clknet_leaf_247_clk net230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_28_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07909__A1 _03622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_1182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10215_ rf_ram.memory\[207\]\[0\] _05098_ _05099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11195_ _00931_ clknet_leaf_5_clk rf_ram.memory\[159\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_24_1166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08582__A1 _04058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07385__A2 _02997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06042__C1 _01610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_37_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10146_ _05049_ _05054_ _05056_ _01284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_37_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06003__C _01495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10077_ _04985_ _05011_ _05013_ _01258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10141__A1 _05049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_195_clk clknet_5_25__leaf_clk clknet_leaf_195_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08885__A2 _04248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05699__A2 _01543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_173_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05414__I _01609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_1165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_1176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10979_ _00716_ clknet_leaf_1_clk rf_ram.memory\[168\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09834__A1 _04837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06648__A1 _02813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_170_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05871__A2 _01641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06170_ rf_ram.memory\[508\]\[1\] _01644_ _01645_ rf_ram.memory\[509\]\[1\] _01636_
+ rf_ram.memory\[511\]\[1\] _02365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_25_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_1071 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_142_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_96_2179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_142_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_124_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_170_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05623__A2 _01677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06820__A1 _02799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_0_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09860_ _04877_ _04880_ _02714_ _01174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_111_2460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_74_1776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08573__A1 _02945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08811_ _04202_ _04203_ _04204_ _00800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09791_ _02945_ _04507_ _04838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_175_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08742_ _01498_ _04158_ _01506_ _04161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_178_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05954_ _02148_ _02149_ _01562_ _02150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08325__A1 _03035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_1076 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08673_ rf_ram.memory\[156\]\[0\] _04117_ _04118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05885_ _02078_ _02080_ _01928_ _02081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xclkbuf_leaf_186_clk clknet_5_28__leaf_clk clknet_leaf_186_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_152_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07624_ _03082_ _03089_ _03452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__06887__A1 _02970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05324__I _01519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07555_ _03393_ _03407_ _03409_ _00339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_75_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06639__A1 _02743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06506_ _02692_ _02693_ _02696_ _00005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_75_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07486_ rf_ram.memory\[365\]\[1\] _03365_ _03367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_5_1160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08635__I _04057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07300__A2 _02941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_153_3228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09225_ rf_ram.memory\[339\]\[0\] _04460_ _04461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_90_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05847__C1 _01725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_153_3239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06437_ rf_ram.memory\[44\]\[1\] _01633_ _01609_ rf_ram.memory\[45\]\[1\] _01607_
+ rf_ram.memory\[47\]\[1\] _02632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_63_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_170_3542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_146_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_185_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_170_3553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05862__A2 _01523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09156_ _04004_ _04418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA_clkbuf_leaf_5_clk_I clknet_5_1__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06368_ rf_ram.memory\[246\]\[1\] _01989_ _02004_ _02563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10199__A1 _02908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08107_ _03724_ _03751_ _03753_ _00547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_121_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07064__A1 _03087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05319_ _01514_ _01515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_47_1144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09087_ _02983_ _03765_ _04375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_110_clk clknet_5_15__leaf_clk clknet_leaf_110_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_131_2825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_130_921 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06299_ _01552_ _02492_ _02493_ _02494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XTAP_TAPCELL_ROW_131_2836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08038_ rf_ram.memory\[568\]\[1\] _03709_ _03711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_82_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_130_987 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06104__B _01684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10000_ _04953_ _04964_ _04966_ _01228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09989_ rf_ram.memory\[503\]\[1\] _04958_ _04960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_122_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_5_5__f_clk clknet_3_1_0_clk clknet_5_5__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_129_2787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_129_2798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_1251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_177_clk clknet_5_31__leaf_clk clknet_leaf_177_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA_clkbuf_leaf_334_clk_I clknet_5_0__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08867__A2 _04195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_170_1321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06878__A1 _02935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10902_ _00646_ clknet_leaf_17_clk rf_ram.memory\[185\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_58_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10833_ _00577_ clknet_leaf_273_clk rf_ram.memory\[540\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_168_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_156_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09816__A1 _04840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_183_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10764_ _00508_ clknet_leaf_126_clk rf_ram.memory\[465\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_39_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06493__C _01373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_884 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_164_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10695_ _00439_ clknet_leaf_83_clk rf_ram.memory\[413\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_152_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_164_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07055__A1 _02806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_101_clk clknet_5_14__leaf_clk clknet_leaf_101_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_50_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_39_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_1266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06802__A1 _02801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11316_ _01049_ clknet_leaf_262_clk net81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_61_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_56_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_56_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11247_ _00983_ clknet_leaf_279_clk cpu.immdec.imm11_7\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_91_2087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_91_2098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05409__I _01499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08555__A1 _04023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07358__A2 _03253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11178_ _00914_ clknet_leaf_57_clk rf_ram.memory\[94\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_52_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06030__A2 _01511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10129_ _05017_ _05043_ _05045_ _01278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08307__A1 _03855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10114__A1 _05017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_1302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_168_clk clknet_5_30__leaf_clk clknet_leaf_168_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__06318__B1 _01772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06869__A1 _02970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_188_954 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05670_ _01850_ _01854_ _01861_ _01865_ _01866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_148_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09807__A1 _02774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_169_1003 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07340_ _03257_ _03274_ _03275_ _00258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_128_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_98_2219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07294__A1 _03225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_14_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07271_ _03222_ _03231_ _03232_ _00232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06097__A2 _01735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_14_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09010_ rf_ram.memory\[110\]\[1\] _04325_ _04327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06222_ rf_ram.memory\[390\]\[1\] _01777_ _01778_ rf_ram.memory\[391\]\[1\] _01793_
+ rf_ram.memory\[389\]\[1\] _02417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_26_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05844__A2 _01808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09035__A2 _04339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07046__A1 _03087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_76_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_170_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06153_ _01597_ _02291_ _02347_ _02348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_TAPCELL_ROW_113_2500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_76_1816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06254__C1 _01726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08794__A1 _04167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06084_ rf_ram.memory\[326\]\[1\] _01706_ _01707_ _02279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_22_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09912_ _04911_ _02992_ _04912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05319__I _01514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08546__A1 _02764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06006__C1 _01520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09843_ cpu.state.cnt_r\[2\] _04869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_146_3098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09774_ _04637_ _04825_ _04827_ _01140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06986_ rf_ram.memory\[227\]\[0\] _03051_ _03052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08725_ rf_ram.memory\[14\]\[0\] _04149_ _04150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05937_ rf_ram.memory\[40\]\[0\] _01682_ _01601_ _02133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xclkbuf_leaf_159_clk clknet_5_27__leaf_clk clknet_leaf_159_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__10105__A1 _02800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06309__B1 _01516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08656_ _04097_ _04105_ _04107_ _00742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05868_ rf_ram.memory\[240\]\[0\] _01683_ _01684_ _02064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07607_ _03425_ _03439_ _03441_ _00359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_77_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_124_2695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_1244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08587_ _02828_ _03949_ _04064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__05532__B2 _01727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05799_ _01992_ _01994_ _01494_ _01995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_113_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07538_ _03389_ _03398_ _03399_ _00332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_165_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_88_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07285__A1 _02836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07469_ _02742_ _03355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
Xclkbuf_leaf_331_clk clknet_5_1__leaf_clk clknet_leaf_331_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_146_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_1206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05835__A2 _01755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09208_ _04434_ _04448_ _04450_ _00951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10480_ _00224_ clknet_leaf_103_clk rf_ram.memory\[420\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_106_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_44_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09139_ rf_ram.memory\[169\]\[1\] _04406_ _04408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_32_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_161_386 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07588__A2 _03390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05599__A1 _01675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11101_ _00837_ clknet_leaf_78_clk rf_ram.memory\[126\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06260__A2 _01755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_1250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_124_1175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_25_1272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11032_ _00769_ clknet_leaf_294_clk rf_ram.memory\[14\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_34_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_183_3788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06012__A2 _01511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_183_3799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05673__B _01650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_273_clk_I clknet_5_16__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06488__C rf_ram.i_raddr\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_188_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_8_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_170_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_1076 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_288_clk_I clknet_5_18__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10816_ _00560_ clknet_leaf_319_clk rf_ram.memory\[548\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_54_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_1265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_322_clk clknet_5_4__leaf_clk clknet_leaf_322_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_83_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10747_ _00491_ clknet_leaf_187_clk rf_ram.memory\[481\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_82_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_211_clk_I clknet_5_28__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05826__A2 _01537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10678_ _00422_ clknet_leaf_110_clk rf_ram.memory\[374\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_70_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07028__A1 _03053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_93_2127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_120_Left_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_65_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput207 net207 o_ibus_adr[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__08776__A1 _04170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput218 net218 o_ibus_adr[24] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_11_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput229 net229 o_ibus_adr[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA_clkbuf_leaf_226_clk_I clknet_5_23__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_71_1713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_71_1724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_1237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_142_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_103_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06840_ _02953_ _02954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_171_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_65_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_179_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06771_ _02881_ _02904_ _02905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_65_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08510_ _04010_ _04011_ _04013_ _04014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05722_ _01514_ _01918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_09490_ cpu.bne_or_bge _01342_ _01442_ _04625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_172_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_19_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_69_1675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_106_2370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07503__A2 _03101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_19_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_69_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08441_ _03953_ _03961_ _03962_ _00672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_188_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_175_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05653_ rf_ram.memory\[470\]\[0\] _01785_ _01786_ rf_ram.memory\[471\]\[0\] _01848_
+ rf_ram.memory\[469\]\[0\] _01849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_0_176_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_1078 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_175_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08372_ _03887_ _03916_ _03918_ _00647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05584_ rf_ram.memory\[298\]\[0\] _01777_ _01778_ rf_ram.memory\[299\]\[0\] _01779_
+ _01780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XTAP_TAPCELL_ROW_102_2289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_635 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07323_ _03055_ _02909_ _03265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07267__A1 _03225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_313_clk clknet_5_5__leaf_clk clknet_leaf_313_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_156_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05817__A2 _01856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07254_ rf_ram.memory\[41\]\[1\] _03219_ _03221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_182_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_30_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06205_ rf_ram.memory\[450\]\[1\] _01801_ _01811_ rf_ram.memory\[451\]\[1\] _01810_
+ rf_ram.memory\[449\]\[1\] _02400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_26_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07019__A1 _03055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_1104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07185_ rf_ram.memory\[198\]\[0\] _03178_ _03179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_108_1115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_565 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_143_1028 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08767__A1 _02945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06136_ rf_ram.memory\[292\]\[1\] _01735_ _02331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_41_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_1125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05477__C net253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_1196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06242__A2 _01787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06067_ _02253_ _02256_ _01599_ _02261_ _02262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XTAP_TAPCELL_ROW_148_3138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_148_3149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08519__A1 _02838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input48_I i_ibus_rdt[23] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_165_3452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_165_3463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09826_ _04840_ _04857_ _04859_ _01160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06545__A3 _02730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_126_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_126_2746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09757_ _04816_ _01134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__05753__A1 _01372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06969_ _02788_ _03040_ _03041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_154_1135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08708_ _04129_ _04137_ _04139_ _00762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_154_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09688_ _04740_ net30 _04769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_115_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_1134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08639_ _04061_ _04097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_11650_ net100 net172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_49_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09247__A2 net56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10601_ _00345_ clknet_leaf_155_clk rf_ram.memory\[357\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11581_ _01313_ clknet_leaf_207_clk rf_ram.memory\[23\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_304_clk clknet_5_4__leaf_clk clknet_leaf_304_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_153_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10532_ _00276_ clknet_leaf_209_clk rf_ram.memory\[24\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_80_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06481__A2 _01686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10463_ _00207_ clknet_leaf_188_clk rf_ram.memory\[273\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_150_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08758__A1 _04170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_60_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10394_ _00138_ clknet_leaf_300_clk rf_ram.memory\[222\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_20_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_185_3828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06233__A2 _01634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05441__B1 _01610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05992__A1 _01371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11015_ _00752_ clknet_leaf_323_clk rf_ram.memory\[559\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09183__A1 _04434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_95_1034 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_92_clk_I clknet_5_11__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06536__A3 _01341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_158_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07497__A1 _03360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_16_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05850__C _01362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_142_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06518__I _01411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_47_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_173_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_150_clk_I clknet_5_26__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_64_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_64_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08997__A1 _02945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_30_clk_I clknet_5_6__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_42_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_181_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_71_969 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06472__A2 _01514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_165_clk_I clknet_5_27__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08749__A1 _04126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_45_clk_I clknet_5_12__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08990_ rf_ram.memory\[114\]\[1\] _04313_ _04315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_11_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_1023 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05432__B1 _01625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07941_ rf_ram.memory\[43\]\[0\] _03648_ _03649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05983__A1 rf_ram.memory\[4\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09174__A1 _04397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07872_ _03590_ _03604_ _03606_ _00459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06202__B _01805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_108_2410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_143_3046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08921__A1 _04266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_143_3057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09611_ rf_ram.memory\[73\]\[1\] _04714_ _04716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06823_ rf_ram.memory\[287\]\[0\] _02942_ _02943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_39_1216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_103_clk_I clknet_5_15__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_160_3360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_183_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_160_3371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06754_ _02876_ _02890_ _02892_ _00055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09542_ _04478_ net41 _04650_ cpu.immdec.imm19_12_20\[5\] _04665_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_TAPCELL_ROW_104_2329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05705_ rf_ram.memory\[406\]\[0\] _01623_ _01504_ _01901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_92_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07488__A1 _02795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09473_ net86 net88 _04604_ _04613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06685_ _02730_ _02732_ _02734_ _02845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XTAP_TAPCELL_ROW_121_2643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_84_1959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_90_clk clknet_5_11__leaf_clk clknet_leaf_90_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_65_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08424_ _03919_ _03950_ _03951_ _00666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05636_ _01820_ _01824_ _01828_ _01831_ _01832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_114_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_136_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_118_clk_I clknet_5_12__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05332__I _01527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_163_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_176_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_1271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08355_ _03884_ _03907_ _03908_ _00640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05567_ _01653_ _01763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_12
XFILLER_0_34_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07306_ _02899_ _03253_ _03254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06448__C1 _01609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08286_ rf_ram.memory\[204\]\[1\] _03863_ _03865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05498_ rf_ram.memory\[336\]\[0\] _01692_ _01693_ _01694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_73_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07237_ rf_ram.memory\[422\]\[0\] _03210_ _03211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_143_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07660__A1 _03458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07168_ _03161_ _03166_ _03168_ _00193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_167_3503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_5_30__f_clk clknet_3_7_0_clk clknet_5_30__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__07412__A1 _03319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06215__A2 _01777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06119_ rf_ram.memory\[260\]\[1\] _01509_ _01668_ rf_ram.memory\[261\]\[1\] _01519_
+ rf_ram.memory\[263\]\[1\] _02314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_100_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_30_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07099_ rf_ram.memory\[48\]\[0\] _03124_ _03125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_112_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05423__B1 _01608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output154_I net154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_180_3736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07715__A2 _03496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09809_ _04837_ _04848_ _04849_ _01153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_92_1218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_2_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_81_clk clknet_5_11__leaf_clk clknet_leaf_81_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_178_3698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_1057 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_96_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06151__A1 _01768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11633_ net83 net156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_181_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_182_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08979__A1 _04298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11564_ _01296_ clknet_leaf_292_clk rf_ram.memory\[20\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_107_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_163_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_42_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07651__A1 net239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06454__A2 _01613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10515_ _00259_ clknet_leaf_191_clk rf_ram.memory\[270\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11495_ _01227_ clknet_leaf_189_clk rf_ram.memory\[276\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_134_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_21_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_150_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10446_ _00190_ clknet_leaf_198_clk rf_ram.memory\[496\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_110_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07403__A1 _03289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10377_ _00121_ clknet_leaf_209_clk rf_ram.memory\[22\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06801__I _02819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_88_2026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06022__B _01506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05417__I _01508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_88_2037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_172_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05861__B _01494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_49_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_1623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_66_1634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_172_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_38_1293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_72_clk clknet_5_8__leaf_clk clknet_leaf_72_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08131__A2 _03765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_1146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06470_ _02662_ _02664_ _01493_ _02665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_34_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_134_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_68_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05421_ _01513_ _01617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_173_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07890__A1 _03587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08140_ _03757_ _03772_ _03774_ _00559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05352_ rf_ram.memory\[534\]\[0\] _01532_ _01505_ _01548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_16_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08071_ rf_ram.memory\[562\]\[1\] _03730_ _03732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_71_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06445__A2 _01605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05283_ _01442_ _01480_ _01452_ _01481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_144_1101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_71_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07022_ rf_ram.memory\[245\]\[1\] _03073_ _03075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05653__B1 _01786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_1253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_122_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_1188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08973_ rf_ram.memory\[117\]\[0\] _04304_ _04305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_162_3400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_162_3411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07924_ _03622_ _03636_ _03638_ _00479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05327__I _01509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07855_ _03587_ _03595_ _03596_ _00452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06806_ rf_ram.memory\[291\]\[1\] _02928_ _02931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07786_ rf_ram.memory\[416\]\[1\] _03551_ _03553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09525_ _01491_ _04652_ _04653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_06737_ rf_ram.memory\[517\]\[1\] _02878_ _02880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_17_1322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_leaf_63_clk clknet_5_8__leaf_clk clknet_leaf_63_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_93_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_66_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06668_ _02831_ _02832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_09456_ _01411_ _04604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_164_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05619_ _01768_ _01796_ _01814_ net253 _01815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_08407_ _03919_ _03939_ _03940_ _00660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_163_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06599_ rf_ram.memory\[234\]\[0\] _02776_ _02777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09387_ _04566_ _01014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_34_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08338_ _03884_ _03896_ _03897_ _00634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08269_ _03852_ _03853_ _03854_ _00608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06436__A2 _01530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_116_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_160_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06107__B _01746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10300_ _00044_ clknet_leaf_316_clk rf_ram.memory\[520\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05644__B1 _01668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_134_2878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11280_ _01015_ clknet_leaf_245_clk net216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_134_2889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_131_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10231_ _05078_ _05107_ _05108_ _01317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08189__A2 _03072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09386__B2 net216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_max_cap248_I _02760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output79_I net79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10162_ _02831_ _02904_ _05066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_100_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_7_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05947__A1 _01903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09138__A1 _04397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10093_ rf_ram.memory\[310\]\[1\] _05022_ _05024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_22_1072 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_92_1026 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_187_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05175__A2 _01376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10995_ _00732_ clknet_leaf_313_clk rf_ram.memory\[539\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_54_clk clknet_5_9__leaf_clk clknet_leaf_54_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09310__A1 _01491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06124__A1 _01674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_155_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_44_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09861__A2 _03035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_1071 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_26_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07872__A1 _03590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_182_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_61_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_61_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11616_ net96 net169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_37_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09613__A2 _04507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_1107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07624__A1 _03082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06427__A2 _01677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11547_ _01279_ clknet_leaf_121_clk rf_ram.memory\[454\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_41_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_123_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_151_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06017__B _01506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_150_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_1248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11478_ _01210_ clknet_leaf_175_clk rf_ram.memory\[337\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_111_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_1318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10429_ _00173_ clknet_leaf_222_clk rf_ram.memory\[488\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_122_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_59_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06060__B1 _01763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05970_ rf_ram.memory\[25\]\[0\] _01514_ _02166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__05147__I _01349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_1037 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_140_3005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_1258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07640_ _03458_ _03460_ _03462_ _00371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_73_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07571_ _02935_ _02960_ _03419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_45_clk clknet_5_12__leaf_clk clknet_leaf_45_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09310_ _01491_ _04013_ _03967_ _04522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_06522_ _01442_ _01376_ _01405_ _01375_ _02710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_81_1907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_119_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_1111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09241_ _01418_ _03989_ _04471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06453_ _01526_ _02646_ _02647_ _02648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_145_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06666__A2 cpu.immdec.imm11_7\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07863__A1 _02774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05404_ _01599_ _01600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_51_1290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05874__B1 _01793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09172_ _03071_ _04418_ _04428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_155_3270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06384_ rf_ram.memory\[72\]\[1\] _01922_ _01551_ _02579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_173_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_161_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_155_3281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_145_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09604__A2 cpu.immdec.imm30_25\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_185_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08123_ rf_ram.memory\[552\]\[1\] _03762_ _03764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_43_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06418__A2 _01706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05335_ _01530_ _01531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_44_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_1217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_116_2553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08054_ _03690_ _03718_ _03720_ _00527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_79_1869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05266_ _01409_ _01464_ _01465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_43_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07005_ rf_ram.memory\[224\]\[1\] _03062_ _03064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_12_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05766__B _01564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05197_ _01389_ _01396_ _01397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_113_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08040__A1 net235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08956_ _04266_ _04292_ _04293_ _00856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input30_I i_dbus_rdt[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07907_ _03619_ _03627_ _03628_ _00472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08887_ _03672_ _02909_ _04251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_98_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09540__A1 _04478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07838_ _03554_ _03584_ _03585_ _00446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_169_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07769_ _03521_ _03541_ _03542_ _00420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05562__C1 _01715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_36_clk clknet_5_6__leaf_clk clknet_leaf_36_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09508_ rf_ram.memory\[279\]\[0\] _04639_ _04640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_1066 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_175_3635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10780_ _00524_ clknet_leaf_325_clk rf_ram.memory\[566\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_39_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_1174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_175_3646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_1099 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06657__A2 _02822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09439_ _04595_ _01037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_23_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_137_779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_136_2918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_136_2929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11401_ _01133_ clknet_leaf_227_clk net116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_152_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06409__A2 _01510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11332_ _01064_ clknet_leaf_240_clk cpu.genblk3.csr.timer_irq_r vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_132_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07082__A2 _02911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09359__A1 net233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06290__B1 _01931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05676__B _01805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11263_ _00998_ clknet_leaf_251_clk net229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_28_1281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_1172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10214_ _03892_ _02954_ _05098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_24_1145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05395__C _01564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11194_ _00930_ clknet_leaf_4_clk rf_ram.memory\[159\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_101_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06042__B1 _01608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10145_ rf_ram.memory\[452\]\[1\] _05054_ _05056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_37_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_37_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09662__I net120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10076_ rf_ram.memory\[308\]\[1\] _05011_ _05013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09531__A1 _04526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06300__B _01956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_186_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_159_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05553__C1 _01625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_27_clk clknet_5_3__leaf_clk clknet_leaf_27_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_58_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08098__A1 _02787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10978_ _00715_ clknet_leaf_1_clk rf_ram.memory\[168\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_70_1165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06648__A2 _02815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05856__B1 _01959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06526__I net65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05430__I _01514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09598__A1 _04478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_993 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_1202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_145_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_41_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_1115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06820__A2 _02939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08022__A1 _03686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_74_1766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_81_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_111_2461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_74_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08810_ rf_ram.memory\[138\]\[0\] _04203_ _04204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08573__A2 _03945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09770__A1 net243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09790_ _04396_ _04837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__05387__A2 _01538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08741_ _02718_ _04158_ _04160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XPHY_EDGE_ROW_183_Right_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05953_ rf_ram.memory\[58\]\[0\] _01661_ _01653_ rf_ram.memory\[59\]\[0\] _01655_
+ rf_ram.memory\[57\]\[0\] _02149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__08325__A2 _03072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08672_ _02838_ _04078_ _04117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_75_1032 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05884_ rf_ram.memory\[74\]\[0\] _01808_ _01925_ rf_ram.memory\[75\]\[0\] _02079_
+ _02080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__05605__I _01661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1065 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07623_ _03425_ _03449_ _03451_ _00365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_5_Right_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_75_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_18_clk clknet_5_2__leaf_clk clknet_leaf_18_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_159_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_157_3310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08916__I _04061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07554_ rf_ram.memory\[31\]\[1\] _03407_ _03409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_119_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_158_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06505_ _01409_ _02695_ _02696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_187_1318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07485_ _03356_ _03365_ _03366_ _00312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07836__A1 _02822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_880 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05847__B1 _01811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_153_3229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09224_ _03319_ _02866_ _04460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_134_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06436_ rf_ram.memory\[46\]\[1\] _01530_ _02631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_161_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05311__A2 _01502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05340__I _01508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_170_3543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09589__A1 _03967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_170_3554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06367_ _02550_ _02554_ _02558_ _02561_ _02562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_09155_ _04401_ _04415_ _04417_ _00931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_32_703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_15_Left_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10199__A2 _03902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08106_ rf_ram.memory\[555\]\[1\] _03751_ _03753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05318_ _01513_ _01514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__08261__A1 _03230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_911 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06298_ rf_ram.memory\[166\]\[1\] _01958_ _01520_ rf_ram.memory\[167\]\[1\] _01516_
+ rf_ram.memory\[165\]\[1\] _02493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_09086_ _04367_ _04372_ _04374_ _00905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_131_2826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_1156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_1036 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_131_2837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08037_ _03686_ _03709_ _03710_ _00520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_47_1178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05249_ _01428_ _01441_ _01446_ _01448_ _01449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_130_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_47_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05378__A2 _01532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06575__A1 _01562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09988_ _04950_ _04958_ _04959_ _01223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_157_1100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_157_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08939_ net245 _04038_ _04283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_output234_I net234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_150_Right_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_129_2788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_24_Left_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_129_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06327__A1 _01951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05515__I _01613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06120__B _01526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_28_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_169_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_168_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10901_ _00645_ clknet_leaf_20_clk rf_ram.memory\[184\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06878__A2 _02844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_79_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_184_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_157_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10832_ _00576_ clknet_leaf_273_clk rf_ram.memory\[540\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_79_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_184_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_67_666 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10763_ _00507_ clknet_leaf_125_clk rf_ram.memory\[466\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10694_ _00438_ clknet_leaf_91_clk rf_ram.memory\[413\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_152_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_33_Left_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_164_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_152_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_164_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07055__A2 _02869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_39_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11315_ _01048_ clknet_leaf_267_clk net80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_120_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06802__A2 _02889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_1109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_120_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_56_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11246_ _00982_ clknet_leaf_258_clk cpu.immdec.imm11_7\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_91_2088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06014__C _01564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06566__A1 _01496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11177_ _00913_ clknet_leaf_62_clk rf_ram.memory\[95\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_42_Left_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08510__B _04013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1016 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_1165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10128_ rf_ram.memory\[475\]\[1\] _05043_ _05045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_98_1076 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_1206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10059_ rf_ram.memory\[507\]\[0\] _05002_ _05003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06030__B _01552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_1314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05526__C1 _01713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_188_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_98_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05541__A2 _01687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_175_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09807__A2 _04004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07818__A1 _03554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_51_Left_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_169_1037 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_85_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07270_ rf_ram.memory\[193\]\[0\] _03231_ _03232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_14_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06221_ rf_ram.memory\[388\]\[1\] _01846_ _02416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_26_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06152_ net252 _02319_ _02346_ _02347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__08243__A1 _03820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_76_1806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_76_1817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_113_2501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_170_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10050__A1 _04982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06254__B1 _01725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06083_ _02266_ _02270_ _02274_ _02277_ _02278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__09991__A1 _02727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_7_clk clknet_5_0__leaf_clk clknet_leaf_7_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_106_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09911_ _02814_ _04911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_106_1054 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06006__B1 _01516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08546__A2 _02867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09842_ _02714_ _04620_ _01167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09773_ rf_ram.memory\[269\]\[1\] _04825_ _04827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06985_ _02766_ _02889_ _03051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_146_3099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08724_ _02971_ _03945_ _04149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05936_ _01903_ _02130_ _02131_ _02132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__10105__A2 _02992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05780__A2 _01915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05335__I _01530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08655_ rf_ram.memory\[160\]\[1\] _04105_ _04107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_7_1201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05867_ rf_ram.memory\[244\]\[0\] _01634_ _01610_ rf_ram.memory\[245\]\[0\] _01636_
+ rf_ram.memory\[247\]\[0\] _02063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_89_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07606_ rf_ram.memory\[314\]\[1\] _03439_ _03441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_178_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_117_1172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_124_2696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_178_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08586_ _04062_ _04059_ _04063_ _00716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05798_ rf_ram.memory\[162\]\[0\] _01958_ _01520_ rf_ram.memory\[163\]\[0\] _01993_
+ _01994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_178_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07537_ rf_ram.memory\[360\]\[0\] _03398_ _03399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_64_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_162_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08482__A1 _03991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_1234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07468_ _03326_ _03352_ _03354_ _00307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07285__A2 _03083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09207_ rf_ram.memory\[6\]\[1\] _04448_ _04450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06419_ _02611_ _02613_ _01928_ _02614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_161_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07399_ rf_ram.memory\[248\]\[1\] _03310_ _03312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09138_ _04397_ _04406_ _04407_ _00924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_output184_I net184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09069_ _04334_ _04361_ _04363_ _00899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06796__A1 _02921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06115__B _01756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_163_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11100_ _00836_ clknet_leaf_78_clk rf_ram.memory\[126\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_102_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_187_3870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_130_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_1240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_1120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11031_ _00768_ clknet_leaf_59_clk rf_ram.memory\[89\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05954__B _01562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_34_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06548__A1 _01353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_183_3789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05771__A2 _01523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_185_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06720__A1 _02797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_1200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_184_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_157_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10815_ _00559_ clknet_leaf_297_clk rf_ram.memory\[54\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_83_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_1255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10746_ _00490_ clknet_leaf_197_clk rf_ram.memory\[481\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_27_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05287__A1 _01341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06009__C _01494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_137_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10677_ _00421_ clknet_leaf_116_clk rf_ram.memory\[393\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_36_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_3_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08225__A1 _03823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_93_2128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05848__C _01717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10032__A1 _04985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput208 net208 o_ibus_adr[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__09973__A1 _04921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_1210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput219 net219 o_ibus_adr[25] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_65_1075 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_1205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_120_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05995__C1 _01521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_71_1714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_71_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11229_ _00965_ clknet_leaf_257_clk cpu.bufreg.i_sh_signed vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09725__B2 net107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06539__A1 _02723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_175_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_175_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06770_ _02903_ _02904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_136_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_1100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10099__A1 _05017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_4_clk_I clknet_5_1__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05721_ rf_ram.memory\[432\]\[0\] _01915_ _01916_ _01917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_136_1036 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_69_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_1193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_78_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_106_2360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_106_2371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08440_ rf_ram.memory\[175\]\[0\] _03961_ _03962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_69_1687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05652_ _01617_ _01848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__05514__A2 _01709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06711__A1 _02826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_1188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_86_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_176_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08371_ rf_ram.memory\[185\]\[1\] _03916_ _03918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_105_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05583_ rf_ram.memory\[297\]\[0\] _01697_ _01779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_74_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09498__S _01491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07322_ _03260_ _03262_ _03264_ _00251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_74_956 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_162_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_18_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_74_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07253_ _03190_ _03219_ _03220_ _00226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_73_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11620__I net70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_30_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06204_ rf_ram.memory\[448\]\[1\] _01649_ _01756_ _02399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_14_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07019__A2 _03072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07184_ _02738_ _02806_ _03178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_121_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_5_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10023__A1 _04950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09964__A1 _03445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06135_ _02327_ _02329_ _01790_ _02330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_clkbuf_leaf_333_clk_I clknet_5_4__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08767__A2 _04152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_160_1321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06778__A1 _02764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_1137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_100_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06066_ _02257_ _02258_ _02259_ _02260_ _01670_ _02261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XTAP_TAPCELL_ROW_148_3139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08519__A2 _03949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09716__A1 _04781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_165_3453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_165_3464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09825_ rf_ram.memory\[249\]\[1\] _04857_ _04859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_126_2736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09756_ net117 _04766_ _04760_ net118 _04815_ _04816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_06968_ _03039_ _03040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_154_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06950__A1 _03018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_1318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08707_ rf_ram.memory\[152\]\[1\] _04137_ _04139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05919_ rf_ram.memory\[124\]\[0\] _01799_ _01931_ rf_ram.memory\[125\]\[0\] _01786_
+ rf_ram.memory\[127\]\[0\] _02115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_69_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09687_ _04760_ _04768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_06899_ _02970_ _02993_ _02994_ _00098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_55_1233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08638_ _04094_ _04095_ _04096_ _00735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_55_1266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_1146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_167_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05505__A2 _01537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06702__A1 _02775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08569_ rf_ram.memory\[170\]\[0\] _04051_ _04052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_77_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10600_ _00344_ clknet_leaf_155_clk rf_ram.memory\[357\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_181_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11580_ _01312_ clknet_leaf_34_clk rf_ram.memory\[207\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_92_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_181_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05269__A1 _01363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_146_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10531_ _00275_ clknet_leaf_192_clk rf_ram.memory\[266\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_18_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09404__B1 _04539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10462_ _00206_ clknet_leaf_189_clk rf_ram.memory\[273\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_126_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_32_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06769__A1 _02716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10393_ _00137_ clknet_leaf_33_clk rf_ram.memory\[223\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_185_3829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09707__A1 _04781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11014_ _00751_ clknet_leaf_323_clk rf_ram.memory\[559\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_159_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_8_Left_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07194__A1 _02813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_240_clk clknet_5_21__leaf_clk clknet_leaf_240_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_5_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06941__A1 _02738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_99_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_158_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08694__A1 _02983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_16_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_158_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_68_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_129_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_185_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05901__C1 _01763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_173_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_172_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_144_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_64_1584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08446__A1 _03953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_64_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10253__A1 _02825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08997__A2 _04303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_1096 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10729_ _00473_ clknet_leaf_51_clk rf_ram.memory\[460\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_183_1310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_1115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_126_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_153_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10005__A1 _04953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09946__A1 _04918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07940_ _02781_ _02869_ _03648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05983__A2 _01643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07871_ rf_ram.memory\[408\]\[1\] _03604_ _03606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_108_2400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_231_clk clknet_5_23__leaf_clk clknet_leaf_231_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09610_ _04634_ _04714_ _04715_ _01088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_108_2411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06822_ _02909_ _02941_ _02942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_143_3047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_1255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_143_3058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06393__C1 _01912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_160_3361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09541_ _01354_ _04654_ _04664_ _01070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_160_3372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06753_ rf_ram.memory\[515\]\[1\] _02890_ _02892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05704_ _01898_ _01899_ _01629_ _01900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__07488__A2 _02815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09472_ _04612_ _01053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_176_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06684_ _02843_ _02844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_121_2644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_149_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08423_ rf_ram.memory\[173\]\[0\] _03950_ _03951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_47_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05635_ _01603_ _01829_ _01830_ _01831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_148_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_1141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08354_ rf_ram.memory\[182\]\[0\] _03907_ _03908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_175_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05566_ rf_ram.memory\[256\]\[0\] _01644_ _01526_ _01762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_163_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10244__A1 _02727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_298_clk clknet_5_7__leaf_clk clknet_leaf_298_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__06448__B1 _01607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07305_ _02940_ _03253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_144_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_1158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08285_ _03852_ _03863_ _03864_ _00614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05497_ _01550_ _01693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_116_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06999__A1 _03050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07236_ _02806_ _03040_ _03210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_171_460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_272_clk_I clknet_5_16__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_85_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_131_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07167_ rf_ram.memory\[483\]\[1\] _03166_ _03168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_167_3504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input60_I i_ibus_rdt[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06118_ rf_ram.memory\[262\]\[1\] _01662_ _01504_ _02313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07412__A2 _02972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07098_ _02921_ _02946_ _03124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_121_1102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_30_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_287_clk_I clknet_5_18__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06049_ rf_ram.memory\[361\]\[1\] _01617_ _02244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_79_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05974__A2 _01633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_180_3737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07176__A1 _03157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09808_ rf_ram.memory\[74\]\[0\] _04848_ _04849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_222_clk clknet_5_22__leaf_clk clknet_leaf_222_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA_clkbuf_leaf_210_clk_I clknet_5_25__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09739_ _04739_ _04804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_2_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08676__A1 _04097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05523__I _01686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_225_clk_I clknet_5_23__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_178_3699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_155_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_5_15__f_clk_I clknet_3_3_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11632_ net82 net155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08428__A1 _02822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_289_clk clknet_5_18__leaf_clk clknet_leaf_289_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_53_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11563_ _01295_ clknet_leaf_292_clk rf_ram.memory\[20\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07100__A1 _03123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_92_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_42_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10514_ _00258_ clknet_leaf_190_clk rf_ram.memory\[270\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07651__A2 _03089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11494_ _01226_ clknet_leaf_137_clk rf_ram.memory\[296\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_134_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_126_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_150_633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_21_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09928__A1 _04921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10445_ _00189_ clknet_leaf_185_clk rf_ram.memory\[484\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_1023 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08600__A1 _04058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10376_ _00120_ clknet_leaf_209_clk rf_ram.memory\[22\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_27_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06303__B _01494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05965__A2 _01682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_88_2027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_213_clk clknet_5_19__leaf_clk clknet_leaf_213_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_88_2038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05717__A2 _01706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06914__A1 _02775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06390__A2 _01808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08667__A1 _02959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_66_1624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_158_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05433__I _01563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_157_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06142__A2 _01799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05420_ rf_ram.memory\[352\]\[0\] _01614_ _01615_ _01616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_158_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09467__I0 net83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10226__A1 _05078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05351_ _01495_ _01534_ _01546_ _01547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_127_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_161_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09092__A1 net238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_172_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08070_ _03721_ _03730_ _03731_ _00532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05282_ _01342_ cpu.alu.i_rs1 _01479_ _01480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__05248__A4 _01388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09919__A1 _04884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07021_ _03050_ _03073_ _03074_ _00140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_114_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_1210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_70_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_178_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_1243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08972_ _03071_ _04303_ _04304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06213__B _01693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05956__A2 _01508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05608__I _01640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_162_3401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_162_3412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07923_ rf_ram.memory\[441\]\[1\] _03636_ _03638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07158__A1 _03161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_204_clk clknet_5_24__leaf_clk clknet_leaf_204_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07854_ rf_ram.memory\[430\]\[0\] _03595_ _03596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05169__B1 _01367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05708__A2 _01634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06805_ _02825_ _02930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_39_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07785_ _03521_ _03551_ _03552_ _00426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_79_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06381__A2 _01531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09524_ _01419_ _04647_ _04652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_78_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06736_ _02873_ _02878_ _02879_ _00050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05343__I _01516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09455_ _04603_ _01045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_176_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06667_ _02736_ _02830_ _02831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_8_1170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06133__A2 _01787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07330__A1 _03257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_563 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08406_ rf_ram.memory\[178\]\[0\] _03939_ _03940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05618_ _01600_ _01803_ _01813_ _01814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_148_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09386_ net215 _04561_ _04564_ net216 _04566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06598_ _02766_ _02775_ _02776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_149_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05892__A1 _01972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08337_ rf_ram.memory\[240\]\[0\] _03896_ _03897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05549_ rf_ram.memory\[282\]\[0\] _01687_ _01696_ rf_ram.memory\[283\]\[0\] _01744_
+ _01745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_TAPCELL_ROW_138_2960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_163_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_145_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08268_ rf_ram.memory\[197\]\[0\] _03853_ _03854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08830__A1 net246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_91_clk_I clknet_5_11__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07219_ rf_ram.memory\[260\]\[1\] _03198_ _03200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_134_2879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08199_ _03798_ _02984_ _03811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_14_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_631 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10230_ rf_ram.memory\[237\]\[0\] _05107_ _05108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_89_Left_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_30_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10161_ _05049_ _05063_ _05065_ _01290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06123__B _01349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_7_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05518__I _01513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10092_ _05014_ _05022_ _05023_ _01263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_156_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08897__A1 net243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_69_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_97_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_164_clk_I clknet_5_27__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_98_Left_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06109__C1 _01625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08649__A1 _04094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10994_ _00731_ clknet_leaf_313_clk rf_ram.memory\[539\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_57_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09310__A2 _04013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_44_clk_I clknet_5_12__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06124__A2 _02306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_44_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_44_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_61_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_179_clk_I clknet_5_29__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10208__A1 _05081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_61_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11615_ net95 net168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_65_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_154_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_59_clk_I clknet_5_9__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11546_ _01278_ clknet_leaf_44_clk rf_ram.memory\[475\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07624__A2 _03089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05635__A1 _01603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_180_1313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_102_clk_I clknet_5_15__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11477_ _01209_ clknet_leaf_168_clk rf_ram.memory\[337\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_34_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_123_666 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_150_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10428_ _00172_ clknet_leaf_184_clk rf_ram.memory\[488\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_123_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_164_Right_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_59_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10359_ _00103_ clknet_leaf_210_clk rf_ram.memory\[27\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06033__B _01505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05428__I _01518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05938__A2 _01513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_117_clk_I clknet_5_14__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07560__A1 _03393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07570_ _03393_ _03416_ _03418_ _00345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_88_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06521_ cpu.state.cnt_r\[1\] cpu.state.cnt_r\[0\] cpu.state.cnt_r\[3\] cpu.state.cnt_r\[2\]
+ _02709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_38_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_81_1908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_158_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06115__A2 _01755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07312__A1 _02904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_186_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_173_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09240_ _04466_ _04468_ _04470_ _00963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_75_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06452_ rf_ram.memory\[60\]\[1\] _01633_ _01609_ rf_ram.memory\[61\]\[1\] _01635_
+ rf_ram.memory\[63\]\[1\] _02647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XANTENNA__06666__A3 _02730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07863__A2 _02869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05403_ _01347_ _01346_ _01598_ _01599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_90_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09171_ _04401_ _04425_ _04427_ _00937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_29_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09065__A1 net237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06383_ _01972_ _02576_ _02577_ _02578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_155_3271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_155_3282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_145_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08122_ _03754_ _03762_ _03763_ _00552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05334_ _01499_ _01530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__07615__A2 _03446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_79_1859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_116_2543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08053_ rf_ram.memory\[565\]\[1\] _03718_ _03720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_43_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_116_2554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05265_ _01333_ cpu.decode.co_ebreak _01337_ _01464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_3_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_109_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07004_ _03050_ _03062_ _03063_ _00134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05196_ cpu.decode.opcode\[0\] cpu.decode.opcode\[1\] _01392_ _01394_ _01395_ _01396_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_109_1085 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_131_Right_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07379__A1 _03292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_995 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_1073 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08040__A2 _03693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05929__A2 _01922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08955_ rf_ram.memory\[120\]\[0\] _04292_ _04293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07906_ rf_ram.memory\[460\]\[0\] _03627_ _03628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08886_ _04237_ _04248_ _04250_ _00829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08879__A1 _04234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input23_I i_dbus_rdt[29] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07837_ rf_ram.memory\[411\]\[0\] _03584_ _03585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09540__A2 net40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06354__A2 _01614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07551__A1 _02909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_1072 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07768_ rf_ram.memory\[393\]\[0\] _03541_ _03542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05562__B1 _01654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09507_ _02958_ _03083_ _04639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06719_ _02798_ _02729_ _02730_ _02867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_67_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_177_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07699_ _03491_ _03497_ _03499_ _00393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06106__A2 _01687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_1078 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_175_3636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_177_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_175_3647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09438_ net69 net70 _04593_ _04595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_93_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_136_2919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09369_ _04556_ _01006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06118__B _01504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11400_ _01132_ clknet_leaf_227_clk net115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_151_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08803__A1 net243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_145_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11331_ _01063_ clknet_leaf_191_clk rf_ram.memory\[279\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_50_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05957__B _01525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11262_ _00997_ clknet_leaf_251_clk net228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_120_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_1140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_30_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10213_ _05081_ _05095_ _05097_ _01310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_11193_ _00929_ clknet_leaf_39_clk rf_ram.memory\[8\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10144_ _05046_ _05054_ _05055_ _01283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_37_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_37_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10075_ _04982_ _05011_ _05012_ _01257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09531__A2 net37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_5_30__f_clk_I clknet_3_7_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05553__B1 _01678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_1100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08098__A2 _03729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10977_ _00714_ clknet_leaf_289_clk rf_ram.memory\[16\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09295__A1 _04463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_183_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_183_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09047__A1 _04331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06028__B _01505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1024 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11529_ _01261_ clknet_leaf_205_clk rf_ram.memory\[30\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_29_1057 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06281__A1 _01951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_150_3190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06542__I _02727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_123_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_111_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_74_1767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_111_2462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_74_1778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09770__A2 _03253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xload_slew243 _02843_ net243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
Xload_slew254 _01361_ net254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_08740_ _04157_ _04159_ _00774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05952_ rf_ram.memory\[56\]\[0\] _01613_ _01601_ _02148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_139_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08671_ _04097_ _04114_ _04116_ _00748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05883_ rf_ram.memory\[73\]\[0\] _01918_ _02079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__07533__A1 _03389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06336__A2 _01531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07622_ rf_ram.memory\[352\]\[1\] _03449_ _03451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_108_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_178_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_36_1039 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_76_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07553_ _03389_ _03407_ _03408_ _00338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_157_3311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11623__I net73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_159_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06504_ _01408_ _02694_ _02695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_76_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07484_ rf_ram.memory\[365\]\[0\] _03365_ _03366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07836__A2 _03559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_146_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_158_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09223_ _04434_ _04457_ _04459_ _00957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_91_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06435_ _01569_ _02618_ _02629_ net251 _02630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_0_119_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09154_ rf_ram.memory\[159\]\[1\] _04415_ _04417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_99_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_173_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_170_3544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06366_ _01951_ _02559_ _02560_ _02561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_173_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_170_3555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_161_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08105_ _03721_ _03751_ _03752_ _00546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05317_ _01512_ _01497_ _01513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_114_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09085_ rf_ram.memory\[98\]\[1\] _04372_ _04374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_130_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06297_ rf_ram.memory\[164\]\[1\] _01523_ _02492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08261__A2 _02844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_131_2827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_131_2838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08036_ rf_ram.memory\[568\]\[0\] _03709_ _03710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05248_ _01442_ _01447_ cpu.alu.cmp_r _01388_ _01448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_141_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05179_ _01377_ _01379_ _00002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09761__A2 net23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09987_ rf_ram.memory\[503\]\[0\] _04958_ _04959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07772__A1 _03008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08938_ _04269_ _04280_ _04282_ _00849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06401__B _01746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_129_2789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_1231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output227_I net227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08869_ _04234_ _04239_ _04240_ _00822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_93_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10900_ _00644_ clknet_leaf_18_clk rf_ram.memory\[184\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_28_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_1106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10831_ _00575_ clknet_leaf_312_clk rf_ram.memory\[541\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_39_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10762_ _00506_ clknet_leaf_124_clk rf_ram.memory\[466\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_149_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_11_Right_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_67_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_165_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_95_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10693_ _00437_ clknet_leaf_80_clk rf_ram.memory\[434\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_125_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05687__B _01693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_1258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_95_2170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06263__A1 _01350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11314_ _01047_ clknet_leaf_267_clk net79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_39_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_56_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11245_ _00981_ clknet_leaf_292_clk rf_ram.memory\[63\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_20_Right_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09201__A1 _04431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_91_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09752__A2 net20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_1022 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11176_ _00912_ clknet_leaf_56_clk rf_ram.memory\[95\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_101_1144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10127_ _05014_ _05043_ _05044_ _01277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_98_1099 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_175_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10058_ _02821_ _03158_ _05002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07515__A1 _03356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06318__A2 _01711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05526__B1 _01721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_72_1239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09268__A1 _01418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_987 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_155_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_14_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06220_ _02412_ _02414_ _01790_ _02415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08752__I _04057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_143_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06151_ _01768_ _02334_ _02345_ net253 _02346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_41_534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_76_1807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_113_2502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_76_1818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06082_ _01603_ _02275_ _02276_ _02277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__09991__A2 _02801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_123_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09910_ _04887_ _04908_ _04910_ _01194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_22_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_186_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_111_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09841_ _02714_ _01384_ _01166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07754__A1 _03521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09772_ _04634_ _04825_ _04826_ _01139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05765__B1 _01959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06984_ _03013_ _03050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_119_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08723_ _04129_ _04146_ _04148_ _00768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05935_ rf_ram.memory\[44\]\[0\] _01633_ _01609_ rf_ram.memory\[45\]\[0\] _01607_
+ rf_ram.memory\[47\]\[0\] _02131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XANTENNA__06309__A2 _01683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08654_ _04094_ _04105_ _04106_ _00741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05866_ rf_ram.memory\[246\]\[0\] _01989_ _02004_ _02062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_14_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07605_ _03422_ _03439_ _03440_ _00358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_178_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08585_ rf_ram.memory\[168\]\[1\] _04059_ _04063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_89_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_124_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05797_ rf_ram.memory\[161\]\[0\] _01664_ _01993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_113_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_1184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_166_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_1075 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07536_ _02728_ _03390_ _03398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_14_1123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_187_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_147_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_36_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_147_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_48_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07467_ rf_ram.memory\[32\]\[1\] _03352_ _03354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_48_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09206_ _04431_ _04448_ _04449_ _00950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06418_ rf_ram.memory\[122\]\[1\] _01706_ _01911_ rf_ram.memory\[123\]\[1\] _02612_
+ _02613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XANTENNA__06493__A1 _02519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07398_ _03289_ _03310_ _03311_ _00280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_44_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09137_ rf_ram.memory\[169\]\[0\] _04406_ _04407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06349_ rf_ram.memory\[194\]\[1\] _01801_ _01811_ rf_ram.memory\[195\]\[1\] _01725_
+ rf_ram.memory\[193\]\[1\] _02544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_103_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09068_ rf_ram.memory\[0\]\[1\] _04361_ _04363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_32_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_956 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06796__A2 _02923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07993__A1 _03654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08019_ _03690_ _03697_ _03699_ _00513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_187_3860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_187_3871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_5_13__f_clk clknet_3_3_0_clk clknet_5_13__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_11030_ _00767_ clknet_leaf_48_clk rf_ram.memory\[89\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_1165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_34_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06131__B _01746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_51_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05220__A2 _01418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08170__A1 _03787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_157_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_1115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06720__A2 _02867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10814_ _00558_ clknet_leaf_297_clk rf_ram.memory\[54\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_68_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_1148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_138_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_172_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10745_ _00489_ clknet_leaf_50_clk rf_ram.memory\[456\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_137_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_840 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_11_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05287__A2 _01484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10676_ _00420_ clknet_leaf_116_clk rf_ram.memory\[393\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_153_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_180_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_180_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_93_2118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_93_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_1032 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput209 net209 o_ibus_adr[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_105_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07984__A1 _03672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05995__B1 _01517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_71_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11228_ _00964_ clknet_leaf_240_clk cpu.genblk3.csr.o_new_irq vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_4
XTAP_TAPCELL_ROW_71_1726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_177_1318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07736__A1 _02813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11159_ _00895_ clknet_leaf_66_clk rf_ram.memory\[101\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09489__A1 _02690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05720_ _01550_ _01916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_76_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_1003 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_106_2361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_157_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_19_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_69_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05651_ rf_ram.memory\[468\]\[0\] _01846_ _01847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_19_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_69_1688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_106_2372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_86_1991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08370_ _03884_ _03916_ _03917_ _00646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05582_ _01695_ _01778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_129_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_73_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07321_ rf_ram.memory\[272\]\[1\] _03262_ _03264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_58_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_45_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07252_ rf_ram.memory\[41\]\[0\] _03219_ _03220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_128_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_1111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_30_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_171_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_143_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06203_ rf_ram.memory\[452\]\[1\] _01724_ _01725_ rf_ram.memory\[453\]\[1\] _01811_
+ rf_ram.memory\[455\]\[1\] _02398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_27_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_30_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_147_1144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07183_ _03161_ _03175_ _03177_ _00199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_60_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06216__B _01746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06227__A1 _01603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06134_ rf_ram.memory\[290\]\[1\] _01785_ _01786_ rf_ram.memory\[291\]\[1\] _02328_
+ _02329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_41_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09964__A2 _02829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06778__A2 _02830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07975__A1 _03651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06065_ rf_ram.memory\[370\]\[1\] _01500_ _01519_ rf_ram.memory\[371\]\[1\] _01664_
+ rf_ram.memory\[369\]\[1\] _02260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_44_1149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07727__A1 _03488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_165_3454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_165_3465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09824_ _04837_ _04857_ _04858_ _01159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06967_ _02797_ _02830_ _03039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_09755_ _04804_ net21 _04815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_126_2737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05753__A3 _01948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05918_ rf_ram.memory\[126\]\[0\] _01770_ _02114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08706_ _04126_ _04137_ _04138_ _00761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09686_ _04766_ _04767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_06898_ rf_ram.memory\[280\]\[0\] _02993_ _02994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_94_1283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_179_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_178_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08637_ rf_ram.memory\[162\]\[0\] _04095_ _04096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_55_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05849_ _02036_ _02039_ _01350_ _02044_ _02045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__06163__B1 _01696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06702__A2 _02846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08568_ net247 _03949_ _04051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_37_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07519_ rf_ram.memory\[322\]\[0\] _03386_ _03387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_182_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_37_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08499_ _04004_ _04005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_119_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_88_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10530_ _00274_ clknet_leaf_192_clk rf_ram.memory\[266\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06466__A1 _01903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_64_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_91_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05674__C1 _01726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10461_ _00205_ clknet_leaf_43_clk rf_ram.memory\[474\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_162_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_70_Left_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_122_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10392_ _00136_ clknet_leaf_33_clk rf_ram.memory\[223\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_32_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_1216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07966__A1 _03654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05965__B _01601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05441__A2 _01634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09707__A2 net5 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_159_1015 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11013_ _00750_ clknet_leaf_3_clk rf_ram.memory\[156\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_102_1283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07194__A2 _02832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06941__A2 _02972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08143__A1 _03754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_386 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_16_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_169_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08694__A2 _04078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09891__A1 _02922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05901__B1 _01656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09643__A1 _04637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_64_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_101_2280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_172_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_64_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10728_ _00472_ clknet_leaf_119_clk rf_ram.memory\[460\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_71_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_109_Left_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_183_1322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10659_ _00403_ clknet_leaf_117_clk rf_ram.memory\[398\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_67_1149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06209__A1 _01368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07957__A1 _02903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05432__A2 _01623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06090__C1 _01713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_1074 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07709__A1 _03491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07870_ _03587_ _03604_ _03605_ _00458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05166__I _01347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08382__A1 _03919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_108_2401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_108_2412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06821_ _02940_ _02941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_143_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_143_3059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06393__B1 _01925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09540_ _04478_ net40 _04650_ cpu.csr_imm _04664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_TAPCELL_ROW_160_3362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06752_ _02873_ _02890_ _02891_ _00054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_160_3373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05703_ rf_ram.memory\[410\]\[0\] _01801_ _01726_ rf_ram.memory\[411\]\[0\] _01721_
+ rf_ram.memory\[409\]\[0\] _01899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_09471_ net85 net86 _04604_ _04612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06683_ _02750_ _02786_ _02843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_78_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_148_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_121_2645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_176_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08422_ net243 _03949_ _03950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06696__A1 _02826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05634_ rf_ram.memory\[486\]\[0\] _01623_ _01688_ rf_ram.memory\[487\]\[0\] _01678_
+ rf_ram.memory\[485\]\[0\] _01830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_176_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_65_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08353_ _03008_ _03903_ _03907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05565_ rf_ram.memory\[260\]\[0\] _01509_ _01668_ rf_ram.memory\[261\]\[0\] _01519_
+ rf_ram.memory\[263\]\[0\] _01761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XANTENNA__09634__A1 _04524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11631__I net81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07304_ _03225_ _03250_ _03252_ _00245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_178_Right_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10244__A2 _02958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08284_ rf_ram.memory\[204\]\[0\] _03863_ _03864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05496_ _01682_ _01692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_132_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07235_ _03193_ _03207_ _03209_ _00219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_132_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_171_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_81_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09398__B1 _04564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_116_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07166_ _03157_ _03166_ _03167_ _00192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05671__A2 _01808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07948__A1 _03651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06117_ _02310_ _02311_ _01629_ _02312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_30_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07097_ _03013_ _03123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA_input53_I i_ibus_rdt[28] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05423__A2 _01606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06081__C1 _01702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06620__A1 _02723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06048_ rf_ram.memory\[360\]\[1\] _01614_ _01615_ _02243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_125_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_180_3727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_1266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_180_3738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09807_ _02774_ _04004_ _04848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07999_ _02742_ _03685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_158_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_2_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09738_ _04803_ _01128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_97_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_2_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_119_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09873__A1 _02713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09669_ _04737_ _03976_ _04752_ _04753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_139_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06687__A1 _02844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_167_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_139_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11631_ net81 net154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_77_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05895__C1 _01773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_46_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08428__A2 _02869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09625__A1 _04637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_166_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_182_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_145_Right_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_11562_ _01294_ clknet_leaf_79_clk rf_ram.memory\[447\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_65_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_42_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10513_ _00257_ clknet_leaf_217_clk rf_ram.memory\[254\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_150_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11493_ _01225_ clknet_leaf_137_clk rf_ram.memory\[296\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_165_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_load_slew243_I _02843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_165_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_21_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10444_ _00188_ clknet_leaf_186_clk rf_ram.memory\[484\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05662__A2 _01787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_3_clk_I clknet_5_1__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_150_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07939__A1 _03622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10375_ _00119_ clknet_leaf_279_clk rf_ram.memory\[230\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_131_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_1057 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_88_2028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_88_2039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05178__A1 _01369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10171__A1 _05049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06914__A2 _02801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_172_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_332_clk_I clknet_5_4__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_66_1625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08667__A2 _04078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_66_1636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_103_2320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_158_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06678__A1 _02836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_1175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_1321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_83_1950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_68_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_157_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09467__I1 net84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_117_Left_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_173_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05350_ _01535_ _01541_ _01542_ _01545_ _01495_ _01546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_172_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_112_Right_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09092__A2 _04339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05638__C1 _01636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05281_ _01342_ _01478_ _01479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_154_995 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_126_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07020_ rf_ram.memory\[245\]\[0\] _03073_ _03074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_12_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05653__A2 _01785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_49_Right_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_109_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_1109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_87_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06063__C1 _01519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06602__A1 _02748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08971_ _04037_ _04303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XPHY_EDGE_ROW_126_Left_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05810__C1 _01679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_162_3402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07922_ _03619_ _03636_ _03637_ _00478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08355__A1 _03884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07853_ _02971_ _03234_ _03595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__05169__A1 _01353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11626__I net76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06804_ _02927_ _02928_ _02929_ _00068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07784_ rf_ram.memory\[416\]\[0\] _03551_ _03552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08107__A1 _03724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_58_Right_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_78_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06735_ rf_ram.memory\[517\]\[0\] _02878_ _02879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09523_ _03992_ net45 _04651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_116_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09855__A1 _02713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_176_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06669__A1 _02829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09454_ net77 net78 _04593_ _04603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_66_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_176_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06666_ cpu.immdec.imm11_7\[3\] cpu.immdec.imm11_7\[4\] _02730_ _02830_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_148_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_135_Left_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05617_ _01806_ _01807_ _01809_ _01812_ _01658_ _01813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_08405_ net236 _03903_ _03939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_176_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09385_ _04565_ _01013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09607__A1 _04643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06597_ net247 _02775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA_clkbuf_5_7__f_clk_I clknet_3_1_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08336_ _03309_ _02946_ _03896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_163_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05548_ rf_ram.memory\[281\]\[0\] _01697_ _01744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_138_2950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_138_2961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07094__A1 _03087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08267_ _03230_ _02795_ _03853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_140_clk clknet_5_27__leaf_clk clknet_leaf_140_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_05479_ _01602_ _01675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_105_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08830__A2 _02832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_1301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_67_Right_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_116_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07218_ _03190_ _03198_ _03199_ _00212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06841__A1 _02935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05644__A2 _01509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_171_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08198_ _03790_ _03808_ _03810_ _00581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_15_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07149_ rf_ram.memory\[497\]\[1\] _03154_ _03156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_144_Left_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06404__B _01602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10160_ rf_ram.memory\[44\]\[1\] _05063_ _05065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_30_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_7_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10091_ rf_ram.memory\[310\]\[0\] _05022_ _05023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08346__A1 _02731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08897__A2 _03547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_173_1310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_76_Right_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_57_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_48_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06109__B1 _01678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_186_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10993_ _00730_ clknet_leaf_308_clk rf_ram.memory\[529\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_153_Left_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_69_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_44_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_182_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_26_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11614_ net94 net167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_53_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05883__A2 _01918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_108_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_85_Right_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_128_1109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11545_ _01277_ clknet_leaf_44_clk rf_ram.memory\[475\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_131_clk clknet_5_24__leaf_clk clknet_leaf_131_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_40_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06293__C1 _01610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11476_ _01208_ clknet_leaf_175_clk rf_ram.memory\[338\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_64_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_162_Left_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_33_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10427_ _00171_ clknet_leaf_220_clk rf_ram.memory\[501\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_104_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06314__B _01916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_59_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10358_ _00102_ clknet_leaf_210_clk rf_ram.memory\[27\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06060__A2 _01500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10289_ _00033_ clknet_leaf_121_clk rf_ram.memory\[476\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_1141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_100_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_94_Right_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10144__A1 _05046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_198_clk clknet_5_28__leaf_clk clknet_leaf_198_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_164_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06899__A1 _02970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_271_clk_I clknet_5_16__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05444__I _01499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_171_Left_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_88_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05571__A1 _01674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09837__A1 cpu.mem_bytecnt\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06520_ _02700_ _02706_ _02708_ _00004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_87_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_81_1909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07312__A2 _03253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10937__D cpu.o_wdata0 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06451_ rf_ram.memory\[62\]\[1\] _01530_ _02646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_158_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_1162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_286_clk_I clknet_5_18__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_146_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_1270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05402_ _01347_ _01478_ _01598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_29_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09170_ rf_ram.memory\[86\]\[1\] _04425_ _04427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05874__A2 _01863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06382_ rf_ram.memory\[76\]\[1\] _01649_ _01912_ rf_ram.memory\[77\]\[1\] _01925_
+ rf_ram.memory\[79\]\[1\] _02577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_7_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09065__A2 _03945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_155_3272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08121_ rf_ram.memory\[552\]\[0\] _03762_ _03763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_43_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05333_ rf_ram.memory\[520\]\[0\] _01524_ _01528_ _01529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07076__A1 _03092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06208__C net254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_122_clk clknet_5_15__leaf_clk clknet_leaf_122_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_16_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_154_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_71_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08052_ _03686_ _03718_ _03719_ _00526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06284__C1 _01911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05626__A2 _01626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_116_2544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_141_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05264_ _01462_ _01463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_25_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_116_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07003_ rf_ram.memory\[224\]\[0\] _03062_ _03063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_141_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05195_ cpu.decode.opcode\[2\] cpu.decode.opcode\[0\] cpu.decode.opcode\[1\] _01395_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_109_1075 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06036__C1 _01539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_45_1085 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_224_clk_I clknet_5_22__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08954_ _02991_ _04038_ _04292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_44_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07905_ _02787_ _02832_ _03627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08885_ rf_ram.memory\[419\]\[1\] _04248_ _04250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_99_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_189_clk clknet_5_29__leaf_clk clknet_leaf_189_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_98_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07836_ _02822_ _03559_ _03584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_239_clk_I clknet_5_21__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05354__I _01525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07551__A2 _02997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input16_I i_dbus_rdt[22] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07767_ _02752_ _03481_ _03541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_155_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_155_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_149_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09506_ _04637_ _04635_ _04638_ _01061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_39_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_1132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06718_ _02865_ _02866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_56_1181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07698_ rf_ram.memory\[382\]\[1\] _03497_ _03499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_67_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08500__A1 _02953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_175_3637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_175_3648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06649_ rf_ram.memory\[346\]\[0\] _02816_ _02817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09437_ _04594_ _01036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_93_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09368_ net206 _04549_ _04552_ net207 _04556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_75_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07067__A1 _02915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08319_ _03309_ _02923_ _03885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_113_clk clknet_5_15__leaf_clk clknet_leaf_113_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_35_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09299_ rf_ram.memory\[66\]\[0\] _04514_ _04515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_118_995 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_23_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08803__A2 _03945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06814__A1 _02935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11330_ _01062_ clknet_leaf_191_clk rf_ram.memory\[279\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_144_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11261_ _00996_ clknet_leaf_250_clk net227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__06290__A2 _01799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_max_cap253_I _01568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output84_I net84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08567__A1 _04026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05529__I _01714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10212_ rf_ram.memory\[442\]\[1\] _05095_ _05097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_127_1197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_120_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11192_ _00928_ clknet_leaf_39_clk rf_ram.memory\[8\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06042__A2 _01606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10143_ rf_ram.memory\[452\]\[0\] _05054_ _05055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_37_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08319__A1 _03309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10074_ rf_ram.memory\[308\]\[0\] _05011_ _05012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_89_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09819__A1 _04837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_1270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10976_ _00713_ clknet_leaf_289_clk rf_ram.memory\[16\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_84_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05856__A2 _01940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_183_876 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_155_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_65_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_104_clk clknet_5_15__leaf_clk clknet_leaf_104_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_109_984 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11528_ _01260_ clknet_leaf_168_clk rf_ram.memory\[350\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_124_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_184_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_150_3180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11459_ _01191_ clknet_leaf_167_clk rf_ram.memory\[345\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06044__B _01615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_1241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06018__C1 _01521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05439__I _01518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08558__A1 _02865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_111_2452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_74_1768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_111_2463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07230__A1 _03193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06033__A2 _01502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_74_1779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xload_slew244 _02821_ net244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_187_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input8_I i_dbus_rdt[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05951_ _01526_ _02145_ _02146_ _02147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__10117__A1 _05014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08670_ rf_ram.memory\[157\]\[1\] _04114_ _04116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05882_ rf_ram.memory\[72\]\[0\] _01922_ _01551_ _02078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_clkbuf_leaf_90_clk_I clknet_5_11__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08730__A1 _03134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07621_ _03422_ _03449_ _03450_ _00364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_36_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_178_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07552_ rf_ram.memory\[31\]\[0\] _03407_ _03408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_177_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_157_3312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06503_ cpu.state.init_done cpu.genblk3.csr.o_new_irq _02694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07297__A1 _03222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07483_ _02844_ _03101_ _03365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_75_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_159_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_119_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09222_ rf_ram.memory\[349\]\[1\] _04457_ _04459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05847__A2 _01801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06434_ _01350_ _02623_ _02628_ _02629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_173_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_146_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_1196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_1051 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07049__A1 _03092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09153_ _04397_ _04415_ _04416_ _00930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06365_ rf_ram.memory\[230\]\[1\] _01940_ _01959_ rf_ram.memory\[231\]\[1\] _01968_
+ rf_ram.memory\[229\]\[1\] _02560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XTAP_TAPCELL_ROW_170_3545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_170_3556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08104_ rf_ram.memory\[555\]\[0\] _03751_ _03752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_44_565 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_146_1028 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05316_ _01496_ _01512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
X_09084_ _04364_ _04372_ _04373_ _00904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06296_ _01674_ _02477_ _02490_ _01362_ _02491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_71_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_131_2828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08035_ _02991_ _03693_ _03709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06272__A2 _01515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_1158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05247_ _01342_ _01447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_141_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_163_clk_I clknet_5_30__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05178_ _01369_ rf_ram.rdata\[0\] _01378_ _01379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA_clkbuf_leaf_43_clk_I clknet_5_13__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07221__A1 _02752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06024__A2 _01524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09986_ _02915_ _03083_ _04958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07772__A2 _03496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10108__A1 rf_ram.memory\[312\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08937_ rf_ram.memory\[399\]\[1\] _04280_ _04282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_178_clk_I clknet_5_31__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_1210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08868_ rf_ram.memory\[130\]\[0\] _04239_ _04240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_99_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_58_clk_I clknet_5_9__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_1205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08721__A1 _04126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07819_ rf_ram.memory\[413\]\[1\] _03572_ _03574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_28_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05535__A1 _01368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_101_clk_I clknet_5_14__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_1313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08799_ rf_ram.memory\[140\]\[0\] _04196_ _04197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_93_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10830_ _00574_ clknet_leaf_274_clk rf_ram.memory\[541\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_95_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_149_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10761_ _00505_ clknet_leaf_120_clk rf_ram.memory\[477\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_334_clk clknet_5_0__leaf_clk clknet_leaf_334_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_94_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_164_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05838__A2 _01531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10692_ _00436_ clknet_leaf_81_clk rf_ram.memory\[434\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_116_clk_I clknet_5_14__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_137_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05968__B _01493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07739__I _03359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_50_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_1247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_95_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11313_ _01046_ clknet_leaf_263_clk net78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_95_2171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_39_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_1269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_946 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11244_ _00980_ clknet_leaf_292_clk rf_ram.memory\[63\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_121_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_56_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11175_ _00911_ clknet_leaf_63_clk rf_ram.memory\[96\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07474__I _02747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10126_ rf_ram.memory\[475\]\[0\] _05043_ _05044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05774__A1 _01951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10057_ _04985_ _04999_ _05001_ _01250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_54_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_72_1218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05722__I _01514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_175_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07279__A1 _03225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_325_clk clknet_5_4__leaf_clk clknet_leaf_325_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10959_ _00696_ clknet_leaf_297_clk rf_ram.memory\[49\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_46_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_85_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06487__C1 _01714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_152_3220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05878__B _01597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_170_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06239__C1 _01931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08779__A1 _04167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06150_ _01600_ _02339_ _02344_ _02345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_108_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_76_1808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_0_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_76_1819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_113_2503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06254__A2 _01724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07451__A1 _03323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06081_ rf_ram.memory\[342\]\[1\] _01623_ _01688_ rf_ram.memory\[343\]\[1\] _01702_
+ rf_ram.memory\[341\]\[1\] _02276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_0_22_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_110_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_1180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_106_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06006__A2 _01523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07203__A1 _03161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09840_ _04867_ _04868_ _02714_ _01165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_111_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08951__A1 _04266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09771_ rf_ram.memory\[269\]\[0\] _04825_ _04826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06983_ _03018_ _03047_ _03049_ _00127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_77_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08722_ rf_ram.memory\[89\]\[1\] _04146_ _04148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05934_ rf_ram.memory\[46\]\[0\] _01530_ _02130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08703__A1 _04129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08653_ rf_ram.memory\[160\]\[0\] _04105_ _04106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05865_ _02049_ _02053_ _02057_ _02060_ _02061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_179_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11634__I net84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07604_ rf_ram.memory\[314\]\[0\] _03439_ _03440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_117_1141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05796_ rf_ram.memory\[160\]\[0\] _01846_ _01956_ _01992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08584_ _04061_ _04062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_48_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_124_2698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_1016 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07535_ _03393_ _03395_ _03397_ _00331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_152_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_316_clk clknet_5_5__leaf_clk clknet_leaf_316_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_64_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07466_ _03323_ _03352_ _03353_ _00306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_92_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06417_ rf_ram.memory\[121\]\[1\] _01918_ _02612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_09205_ rf_ram.memory\[6\]\[0\] _04448_ _04449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07397_ rf_ram.memory\[248\]\[0\] _03310_ _03311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_17_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_1269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09136_ net249 _04067_ _04406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_72_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06348_ rf_ram.memory\[192\]\[1\] _01649_ _01650_ _02543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_32_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09067_ _04331_ _04361_ _04362_ _00898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06245__A2 _01922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06279_ rf_ram.memory\[148\]\[1\] _01523_ _02474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_60_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08018_ rf_ram.memory\[572\]\[1\] _03697_ _03699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_187_3861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_187_3872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_1310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06412__B _01916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_34_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_34_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_1188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09969_ _03672_ _02946_ _04947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_51_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05508__A1 _01603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06181__A1 _01600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10813_ _00557_ clknet_leaf_318_clk rf_ram.memory\[550\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_0_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_307_clk clknet_5_4__leaf_clk clknet_leaf_307_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_0_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_149_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10744_ _00488_ clknet_leaf_49_clk rf_ram.memory\[456\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_165_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_97_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_152_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_137_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07681__A1 _03458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_11_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06484__A2 _01640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10675_ _00419_ clknet_leaf_113_clk rf_ram.memory\[394\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_180_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_82_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07469__I _02742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_1034 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_93_2119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_180_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07433__A1 _03326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_1089 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_65_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07984__A2 _02866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_181_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_121_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09186__A1 _04431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11227_ _00963_ clknet_leaf_153_clk rf_ram.memory\[319\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_71_1716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_71_1727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07736__A2 _03496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08933__A1 _04269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11158_ _00894_ clknet_leaf_66_clk rf_ram.memory\[101\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10109_ _05017_ _05031_ _05033_ _01270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_11089_ _00826_ clknet_leaf_25_clk rf_ram.memory\[128\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_145_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_159_Right_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_37_1135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05650_ _01536_ _01846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_106_2362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_172_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_19_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_69_1678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_106_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_69_1689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_86_1992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05581_ _01686_ _01777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_169_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07320_ _03257_ _03262_ _03263_ _00250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_129_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_1071 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07251_ _02752_ _02869_ _03219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_183_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_156_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07672__A1 _02904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06475__A2 _01530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_183_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06202_ rf_ram.memory\[454\]\[1\] _01804_ _01805_ _02397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_30_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_116_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07182_ rf_ram.memory\[1\]\[1\] _03175_ _03177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_14_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_1100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_26_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_1107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_171_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06133_ rf_ram.memory\[289\]\[1\] _01787_ _02328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_131_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07424__A1 _03319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06064_ rf_ram.memory\[368\]\[1\] _01666_ _01526_ _02259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_111_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11629__I net79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_165_3455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08924__A1 _02838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_165_3466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09823_ rf_ram.memory\[249\]\[0\] _04857_ _04858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_182_3780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09754_ _04814_ _01133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_20_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06966_ _03018_ _03036_ _03038_ _00121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_126_2738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08705_ rf_ram.memory\[152\]\[0\] _04137_ _04138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05917_ _02110_ _02112_ _01928_ _02113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_20_1194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05790__C _01349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09685_ _04739_ _01401_ _04733_ _04766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_06897_ _02958_ _02992_ _02993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_119_1258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_93_clk clknet_5_14__leaf_clk clknet_leaf_93_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_90_1115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_126_Right_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08636_ _02893_ _04067_ _04095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_96_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05848_ _02040_ _02041_ _02042_ _02043_ _01717_ _02044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_08567_ _04026_ _04048_ _04050_ _00710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_138_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05779_ _01972_ _01973_ _01974_ _01975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_77_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09101__A1 _04367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07518_ _03319_ _02894_ _03386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08498_ _02736_ _02867_ _04004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_88_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07663__A1 _03455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07449_ _02946_ _03101_ _03343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_36_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06407__B _01660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05674__B1 _01725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05311__B _01506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_1077 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10460_ _00204_ clknet_leaf_43_clk rf_ram.memory\[474\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_161_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_165_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06218__A2 _01787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09119_ _04364_ _04393_ _04394_ _00918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_103_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_1218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10391_ _00135_ clknet_leaf_275_clk rf_ram.memory\[224\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_60_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_103_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06921__I _03008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06142__B _01602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08915__A1 _04266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11012_ _00749_ clknet_leaf_29_clk rf_ram.memory\[156\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_159_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_1314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_5_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_172_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_84_clk clknet_5_10__leaf_clk clknet_leaf_84_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09340__A1 cpu.ctrl.pc vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09340__B2 net213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_16_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09891__A2 _03035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_185_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08583__I _02747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_64_1586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_101_2270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_64_1597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_101_2281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10727_ _00471_ clknet_leaf_54_clk rf_ram.memory\[444\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_32_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06457__A2 _01661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_165_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_153_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06317__B _01505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10658_ _00402_ clknet_leaf_117_clk rf_ram.memory\[398\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07406__A1 _03100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06209__A2 _02376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10589_ _00333_ clknet_leaf_159_clk rf_ram.memory\[360\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07957__A2 _03158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05875__C _01860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09159__A1 _04397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06090__B1 _01715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_1150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_147_3130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05447__I _01508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08906__A1 _04237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_108_2402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06820_ _02799_ _02939_ _02940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XTAP_TAPCELL_ROW_108_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_143_3049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_1208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05196__A2 cpu.decode.opcode\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06751_ rf_ram.memory\[515\]\[0\] _02890_ _02891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_92_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_160_3363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_160_3374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_75_clk clknet_5_10__leaf_clk clknet_leaf_75_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_78_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05702_ rf_ram.memory\[408\]\[0\] _01614_ _01615_ _01898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06682_ _02826_ _02840_ _02842_ _00033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09470_ _04611_ _01052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_176_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_149_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08421_ _03902_ _03949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_TAPCELL_ROW_121_2646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_148_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05633_ rf_ram.memory\[484\]\[0\] _01735_ _01829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_118_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_175_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05353__C1 _01520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_1144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_1239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08352_ _03887_ _03904_ _03906_ _00639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_86_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05564_ rf_ram.memory\[262\]\[0\] _01662_ _01504_ _01760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_74_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07303_ rf_ram.memory\[258\]\[1\] _03250_ _03252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07645__A1 _03458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06448__A2 _01661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05495_ _01685_ _01690_ _01629_ _01691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08283_ _03230_ _02788_ _03863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_6_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07234_ rf_ram.memory\[423\]\[1\] _03207_ _03209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05131__B cpu.decode.co_ebreak vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07165_ rf_ram.memory\[483\]\[0\] _03166_ _03167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_131_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06116_ rf_ram.memory\[266\]\[1\] _01652_ _01654_ rf_ram.memory\[267\]\[1\] _01715_
+ rf_ram.memory\[265\]\[1\] _02311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XANTENNA__06741__I net241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08070__A1 _03721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07096_ _03092_ _03120_ _03122_ _00167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_112_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06081__B1 _01688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06047_ _02239_ _02241_ _01620_ _02242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_140_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input46_I i_ibus_rdt[21] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_180_3728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_180_3739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09806_ _04840_ _04845_ _04847_ _01152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07998_ _03654_ _03682_ _03684_ _00507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09737_ net111 _04790_ _04791_ net112 _04802_ _04803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_06949_ rf_ram.memory\[232\]\[1\] _03026_ _03028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_2_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_1106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_66_clk clknet_5_8__leaf_clk clknet_leaf_66_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09668_ net120 _03975_ net123 _04752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_179_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_167_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09873__A2 _01413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08619_ _04062_ _04082_ _04084_ _00728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_output202_I net202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06687__A2 _02846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09599_ _04700_ _04704_ _04707_ _04708_ _01084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_16_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_139_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05895__B1 _01772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11630_ net80 net153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_46_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_167_779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_46_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_1318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_166_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07636__A1 _03008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06439__A2 _01613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11561_ _01293_ clknet_leaf_53_clk rf_ram.memory\[447\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_135_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_25_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10512_ _00256_ clknet_leaf_220_clk rf_ram.memory\[254\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_162_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11492_ _01224_ clknet_leaf_220_clk rf_ram.memory\[503\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_150_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10443_ _00187_ clknet_leaf_221_clk rf_ram.memory\[497\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08061__A1 _03724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_1059 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10374_ _00118_ clknet_leaf_278_clk rf_ram.memory\[230\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_1178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_5_24__f_clk_I clknet_3_6_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_88_2029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_1070 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08578__I _02742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_57_clk clknet_5_9__leaf_clk clknet_leaf_57_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__06127__A1 _01769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_103_2310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_1188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_66_1626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_73_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_87_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_1285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06678__A2 _02839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07875__A1 _03587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_1198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_83_1940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06047__B _01620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05638__B1 _01610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05280_ cpu.csr_imm _01478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_153_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_125_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_125_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05886__B _01551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08052__A1 _03686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06063__B1 _01664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08970_ _04301_ _04299_ _04302_ _00861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_87_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05810__B1 _01793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07921_ rf_ram.memory\[441\]\[0\] _03636_ _03637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_162_3403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09552__A1 _04478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07852_ _03590_ _03592_ _03594_ _00451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06366__A1 _01951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10162__A2 _02904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06803_ rf_ram.memory\[291\]\[0\] _02928_ _02929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput1 i_dbus_ack net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_07783_ net237 _03234_ _03551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_78_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_48_clk clknet_5_12__leaf_clk clknet_leaf_48_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_39_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09522_ _04649_ _04650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_06734_ _02795_ _02846_ _02878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_149_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09855__A2 _01418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06669__A2 _02832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09453_ _04602_ _01044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06665_ _02828_ _02829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__05326__C1 _01521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_1150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08404_ _03922_ _03936_ _03938_ _00659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05616_ rf_ram.memory\[312\]\[0\] _01666_ _01810_ rf_ram.memory\[313\]\[0\] _01811_
+ rf_ram.memory\[315\]\[0\] _01812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_59_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09384_ net214 _04561_ _04564_ net215 _04565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_148_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06596_ _02773_ _02726_ _02774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__07618__A1 _03425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_1069 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08335_ _03887_ _03893_ _03895_ _00633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05547_ rf_ram.memory\[280\]\[0\] _01692_ _01684_ _01743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_129_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_138_2951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_138_2962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_173_3598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08266_ _03685_ _03852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_05478_ _01349_ _01674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_117_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07217_ rf_ram.memory\[260\]\[0\] _03198_ _03199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_160_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06841__A2 _02954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09268__B _01366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05796__B _01956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08197_ rf_ram.memory\[538\]\[1\] _03808_ _03810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_160_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07148_ _03123_ _03154_ _03155_ _00186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_30_633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09791__A1 _02945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07079_ _03087_ _03111_ _03112_ _00160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_7_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10090_ _03445_ _03009_ _05022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08346__A2 _02797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_173_1322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05565__C1 _01519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_39_clk clknet_5_7__leaf_clk clknet_leaf_39_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_97_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_48_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10992_ _00729_ clknet_leaf_307_clk rf_ram.memory\[529\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05580__A2 _01692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07857__A1 _03590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_919 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05550__I _01563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11613_ net93 net166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_61_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_182_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_0_clk_I clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11544_ _01276_ clknet_leaf_117_clk rf_ram.memory\[438\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08282__A1 _03855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06293__B1 _01608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05635__A3 _01830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11475_ _01207_ clknet_leaf_175_clk rf_ram.memory\[338\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_150_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08034__A1 _03690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10426_ _00170_ clknet_leaf_220_clk rf_ram.memory\[501\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09782__A1 _04634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_59_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10357_ _00101_ clknet_leaf_292_clk rf_ram.memory\[2\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06596__A1 _02773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10288_ _00032_ clknet_leaf_123_clk rf_ram.memory\[476\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09534__A1 _04526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_1197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_178_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05571__A2 _01751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09837__A2 _01385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07848__A1 _02813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_186_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_180_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06450_ _02633_ _02637_ _02641_ _02644_ _02645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_111_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05460__I _01655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_29_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05401_ _01369_ _01595_ _01596_ _01597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_84_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06381_ rf_ram.memory\[78\]\[1\] _01531_ _02576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_28_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_155_3273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05332_ _01527_ _01528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_08120_ _02728_ _03729_ _03762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_83_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08273__A1 _03230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_1288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06284__B1 _01912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05263_ cpu.state.cnt_r\[3\] _01460_ _01386_ _01461_ _01462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_08051_ rf_ram.memory\[565\]\[0\] _03718_ _03719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_148_1070 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_116_2545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_153_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_116_2556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_142_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07002_ _03055_ _02904_ _03062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_142_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_40_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08025__A1 _02813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05194_ _01380_ _01393_ cpu.branch_op _01394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_133_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_141_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06036__B1 _01540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06587__A1 _02743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08953_ _04269_ _04289_ _04291_ _00855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11637__I net88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09525__A1 _01491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07904_ _03622_ _03624_ _03626_ _00471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08884_ _04234_ _04248_ _04249_ _00828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_138_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07835_ _03557_ _03581_ _03583_ _00445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_155_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07766_ _03524_ _03538_ _03540_ _00419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05562__A2 _01652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_2_clk_I clknet_5_1__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09505_ rf_ram.memory\[289\]\[1\] _04635_ _04638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06717_ _02779_ _02759_ _02865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_116_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07697_ _03488_ _03497_ _03498_ _00392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_116_1058 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08500__A2 _04005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_175_3638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09436_ net68 net69 _04593_ _04594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_175_3649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06648_ _02813_ _02815_ _02816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06511__A1 cpu.alu.i_rs1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_1079 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_23_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09367_ _04555_ _01005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06579_ _02760_ _02761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_118_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08318_ _03685_ _03884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__07067__A2 _02972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09298_ net239 _04507_ _04514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_62_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06814__A2 _02904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08249_ rf_ram.memory\[528\]\[1\] _03840_ _03842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06415__B _01790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11260_ _00995_ clknet_leaf_250_clk net224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA_clkbuf_leaf_331_clk_I clknet_5_1__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10211_ _05078_ _05095_ _05096_ _01309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_162_1078 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_max_cap246_I _02780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11191_ _00927_ clknet_leaf_57_clk rf_ram.memory\[90\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_140_1321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06578__A1 _02750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output77_I net77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10142_ _03672_ _02883_ _05054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput190 net190 o_ext_rs2[28] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_98_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09516__A1 _04524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08319__A2 _02923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10073_ _03445_ _03134_ _05011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__09017__I _04057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_wire249_I _02751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05553__A2 _01634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06750__A1 _02881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10975_ _00712_ clknet_leaf_8_clk rf_ram.memory\[170\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_134_1169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_1266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_5_0__f_clk clknet_3_0_0_clk clknet_5_0__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_84_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_563 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09687__I _04760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08255__A1 _03823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_170_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_68_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_25_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10062__A1 _04985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11527_ _01259_ clknet_leaf_168_clk rf_ram.memory\[350\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_124_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_163_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_78_1850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08007__A1 _03690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_150_3181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11458_ _01190_ clknet_leaf_138_clk rf_ram.memory\[263\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_111_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06018__B1 _01517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_110_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08558__A2 _03158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10409_ _00153_ clknet_leaf_129_clk rf_ram.memory\[38\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_111_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11389_ _01121_ clknet_leaf_225_clk net103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__06569__A1 _02738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_74_1769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_111_2453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_111_2464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xload_slew245 _02812_ net245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__05241__A1 _01343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09507__A1 _02958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05950_ rf_ram.memory\[60\]\[0\] _01633_ _01609_ rf_ram.memory\[61\]\[0\] _01635_
+ rf_ram.memory\[63\]\[0\] _02146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XANTENNA__05792__A2 _01523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_1036 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_139_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05881_ _01972_ _02075_ _02076_ _02077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_108_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07620_ rf_ram.memory\[352\]\[0\] _03449_ _03450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08730__A2 _04152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1057 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05544__A2 _01626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1079 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07551_ _02909_ _02997_ _03407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_157_3302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_159_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_157_3313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06502_ cpu.state.cnt_r\[2\] _01386_ _01471_ _02693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_07482_ _03360_ _03362_ _03364_ _00311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09221_ _04431_ _04457_ _04458_ _00956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_33_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_118_215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06433_ _02624_ _02625_ _02626_ _02627_ _01978_ _02628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_57_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_173_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08246__A1 _03798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09152_ rf_ram.memory\[159\]\[0\] _04415_ _04416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_133_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06364_ rf_ram.memory\[228\]\[1\] _01523_ _02559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_127_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_135_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_170_3546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_170_3557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08103_ _02780_ _03729_ _03751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_114_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05315_ _01510_ _01511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_71_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_154_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06295_ _02480_ _02483_ _02486_ _02489_ _01349_ _02490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_09083_ rf_ram.memory\[98\]\[0\] _04372_ _04373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_163_1310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_140_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_82_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_47_1148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08034_ _03690_ _03706_ _03708_ _00519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_131_2829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05246_ _01442_ _01443_ _01445_ _01446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_114_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_130_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05177_ rf_ram.regzero _01378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_101_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08450__B _03967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07845__I _03359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07221__A2 _03040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09985_ _04953_ _04955_ _04957_ _01222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_0_880 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_1073 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08936_ _04266_ _04280_ _04281_ _00848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_23_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_99_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08867_ net239 _04195_ _04239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_93_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_1109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07818_ _03554_ _03572_ _03573_ _00438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_58_1255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_28_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07580__I _03359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_28_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08798_ _02787_ _04195_ _04196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07749_ _03521_ _03529_ _03530_ _00412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_output115_I net115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_94_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08485__A1 _03953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10760_ _00504_ clknet_leaf_120_clk rf_ram.memory\[477\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_39_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09419_ net90 net91 _02707_ _04585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_48_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10691_ _00435_ clknet_leaf_91_clk rf_ram.memory\[414\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_168_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_165_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_125_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_875 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09985__A1 _04953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_180_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06145__B _01805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_270_clk_I clknet_5_16__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11312_ _01045_ clknet_leaf_265_clk net77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_95_2161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_95_2172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_39_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_160_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05984__B _01525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11243_ _00979_ clknet_leaf_60_clk rf_ram.memory\[66\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_56_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_56_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11174_ _00910_ clknet_leaf_62_clk rf_ram.memory\[96\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_285_clk_I clknet_5_18__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_270_clk clknet_5_16__leaf_clk clknet_leaf_270_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10125_ net244 _02832_ _05043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_101_1146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06971__A1 _03014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10056_ rf_ram.memory\[34\]\[1\] _04999_ _05001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_37_1306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05526__A2 _01709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_11_Left_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_187_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_174_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10958_ _00695_ clknet_leaf_296_clk rf_ram.memory\[49\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_58_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_223_clk_I clknet_5_29__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06039__C _01362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06487__B1 _01635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_183_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10889_ _00633_ clknet_leaf_301_clk rf_ram.memory\[217\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_186_1321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_152_3210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08228__A1 _03820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_152_3221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_26_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_171_847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10035__A1 _04982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06239__B1 _01911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_238_clk_I clknet_5_21__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_76_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_113_2504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06080_ rf_ram.memory\[340\]\[1\] _01537_ _02275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_112_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_9_Right_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09728__A1 net107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08400__A1 _03892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05214__A1 net134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_261_clk clknet_5_17__leaf_clk clknet_leaf_261_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_EDGE_ROW_107_Right_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09770_ net243 _03253_ _04825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06982_ rf_ram.memory\[426\]\[1\] _03047_ _03049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_3_6_0_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05765__A2 _01958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06962__A1 _03035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08721_ _04126_ _04146_ _04147_ _00767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05933_ _01569_ _02117_ _02128_ net251 _02129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_0_179_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09900__A1 _04887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_128_2780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08652_ net237 _04067_ _04105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05864_ _01951_ _02058_ _02059_ _02060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__06714__A1 _02820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07603_ _02935_ _02813_ _03439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_178_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08583_ _02747_ _04061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_77_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05795_ _01552_ _01988_ _01990_ _01991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_77_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_89_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06190__A2 _01787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_124_2699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07534_ rf_ram.memory\[321\]\[1\] _03395_ _03397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_88_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_1196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07465_ rf_ram.memory\[32\]\[0\] _03352_ _03353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_29_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_174_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09204_ _02805_ _03035_ _04448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06416_ rf_ram.memory\[120\]\[1\] _01915_ _01916_ _02611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_45_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_63_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07396_ _03309_ _02992_ _03310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_146_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_134_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09135_ _04401_ _04403_ _04405_ _00923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06347_ rf_ram.memory\[196\]\[1\] _01709_ _01721_ rf_ram.memory\[197\]\[1\] _01713_
+ rf_ram.memory\[199\]\[1\] _02542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_161_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09066_ rf_ram.memory\[0\]\[0\] _04361_ _04362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06278_ _02470_ _02472_ _01494_ _02473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_115_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08017_ _03686_ _03697_ _03698_ _00512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_13_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05229_ cpu.alu.i_rs1 cpu.alu.add_cy_r _01429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_187_3862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_187_3873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_1232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_124_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_130_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_60_1145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_90_2080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_34_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_252_clk clknet_5_20__leaf_clk clknet_leaf_252_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_34_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09968_ _04921_ _04944_ _04946_ _01216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05756__A2 _01501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06953__A1 _03014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_51_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08919_ _02794_ _03559_ _04271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_output232_I net232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_51_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09899_ rf_ram.memory\[263\]\[1\] _04902_ _04904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_99_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06166__C1 _01702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05823__I _01695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10812_ _00556_ clknet_leaf_318_clk rf_ram.memory\[550\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_67_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_0_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06469__B1 _01624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05979__B _01525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10743_ _00487_ clknet_leaf_128_clk rf_ram.memory\[43\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_67_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07130__A1 _03126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_137_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_97_2201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06654__I _02819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10674_ _00418_ clknet_leaf_116_clk rf_ram.memory\[394\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_36_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_152_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09958__A1 _04921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_1057 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_50_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08630__A1 _02794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_181_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_142_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05995__A2 _01511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11226_ _00962_ clknet_leaf_153_clk rf_ram.memory\[319\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_121_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_71_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_71_1728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_243_clk clknet_5_21__leaf_clk clknet_leaf_243_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_11157_ _00893_ clknet_leaf_63_clk rf_ram.memory\[102\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05747__A2 _01755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10108_ rf_ram.memory\[312\]\[1\] _05031_ _05033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11088_ _00825_ clknet_leaf_295_clk rf_ram.memory\[12\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_145_3080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_145_3091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10039_ rf_ram.memory\[305\]\[0\] _04990_ _04991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_136_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_76_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_1185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_1147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_19_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_69_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_1027 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_106_2363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06172__A2 _01755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_106_2374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_162_clk_I clknet_5_30__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_176_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_175_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_187_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05580_ rf_ram.memory\[296\]\[0\] _01692_ _01693_ _01776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_86_1993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_175_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10256__A1 _02819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05889__B _01978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_42_clk_I clknet_5_13__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07121__A1 _02829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07250_ _03193_ _03216_ _03218_ _00225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_128_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_177_clk_I clknet_5_31__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_875 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05683__A1 _01368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06201_ _02392_ _02393_ _02394_ _02395_ _01658_ _02396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__10008__A1 _04950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09949__A1 net248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07181_ _03157_ _03175_ _03176_ _00198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_30_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_48_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06132_ rf_ram.memory\[288\]\[1\] _01782_ _01783_ _02327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_48_1243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_57_clk_I clknet_5_9__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07424__A2 _02844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_100_clk_I clknet_5_14__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_1313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06063_ rf_ram.memory\[372\]\[1\] _01536_ _01664_ rf_ram.memory\[373\]\[1\] _01519_
+ rf_ram.memory\[375\]\[1\] _02258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_83_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07188__A1 _03161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09822_ _03309_ _02984_ _04857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_165_3456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08924__A2 _04038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_165_3467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06935__A1 _03018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_115_clk_I clknet_5_15__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_182_3770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09753_ net116 _04766_ _04760_ net117 _04813_ _04814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XTAP_TAPCELL_ROW_182_3781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06965_ rf_ram.memory\[22\]\[1\] _03036_ _03038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_126_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11645__I net126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_126_2739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08704_ _02991_ _04078_ _04137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05916_ rf_ram.memory\[122\]\[0\] _01706_ _01911_ rf_ram.memory\[123\]\[0\] _02111_
+ _02112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XANTENNA__06148__C1 _01811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08688__A1 _02812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06739__I _02845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09684_ _04763_ _04736_ _04764_ _04765_ _01112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_158_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06896_ _02991_ _02992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_08635_ _04057_ _04094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_05847_ rf_ram.memory\[194\]\[0\] _01801_ _01811_ rf_ram.memory\[195\]\[0\] _01725_
+ rf_ram.memory\[193\]\[0\] _02043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_167_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_167_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_96_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06163__A2 _01687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07360__A1 _03257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08566_ rf_ram.memory\[509\]\[1\] _04048_ _04050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05778_ rf_ram.memory\[132\]\[0\] _01649_ _01912_ rf_ram.memory\[133\]\[0\] _01925_
+ rf_ram.memory\[135\]\[0\] _01974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_76_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05910__A2 _01915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07517_ _03360_ _03383_ _03385_ _00325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05799__B _01494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08497_ _03956_ _04001_ _04003_ _00687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_91_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_639 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07448_ _03326_ _03340_ _03342_ _00299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_130_1172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_107_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06320__C1 _01931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07379_ _03292_ _03297_ _03299_ _00273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_134_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09118_ rf_ram.memory\[575\]\[0\] _04393_ _04394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10390_ _00134_ clknet_leaf_275_clk rf_ram.memory\[224\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08612__A1 _04058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09049_ _04334_ _04349_ _04351_ _00891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_130_563 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05977__A2 _01640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07179__A1 _02899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11011_ _00748_ clknet_leaf_3_clk rf_ram.memory\[157\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_225_clk clknet_5_23__leaf_clk clknet_leaf_225_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__06926__A1 _02975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_1174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05981__C _01562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08679__A1 _04094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09340__A2 _03991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06154__A2 _01543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_16_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08864__I _04061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05901__A2 _01709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10238__A1 _02825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_775 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_173_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07103__A1 _03126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_101_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_64_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_101_2282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10726_ _00470_ clknet_leaf_78_clk rf_ram.memory\[444\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_64_1598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_1107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_126_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10657_ _00401_ clknet_leaf_106_clk rf_ram.memory\[380\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_152_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_141_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07406__A2 _03135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08603__A1 net241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06209__A3 _02403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_180_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10588_ _00332_ clknet_leaf_159_clk rf_ram.memory\[360\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_23_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_121_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_147_3120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_1027 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_147_3131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_142_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_216_clk clknet_5_22__leaf_clk clknet_leaf_216_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_76_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11209_ _00945_ clknet_leaf_47_clk rf_ram.memory\[83\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_108_2403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07590__A1 _03422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06393__A2 _01719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06750_ _02881_ _02889_ _02890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_160_3364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_162_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_160_3375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05701_ _01603_ _01895_ _01896_ _01897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_78_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06681_ rf_ram.memory\[476\]\[1\] _02840_ _02842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06145__A2 _01804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07342__A1 _03260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08420_ _03922_ _03946_ _03948_ _00665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_121_2636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05632_ _01825_ _01827_ _01620_ _01828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__05353__B1 _01516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_121_2647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_1231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08351_ rf_ram.memory\[181\]\[1\] _03904_ _03906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05563_ _01757_ _01758_ _01629_ _01759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07302_ _03222_ _03250_ _03251_ _00244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_11_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_74_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08282_ _03855_ _03860_ _03862_ _00613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05494_ rf_ram.memory\[346\]\[0\] _01687_ _01688_ rf_ram.memory\[347\]\[0\] _01689_
+ _01690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__08842__A1 _04202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07233_ _03190_ _03207_ _03208_ _00218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_4_Left_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_14_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07164_ _02889_ _03158_ _03166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_30_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06115_ rf_ram.memory\[264\]\[1\] _01755_ _01756_ _02310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07095_ rf_ram.memory\[502\]\[1\] _03120_ _03122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_112_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_563 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_184_3810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06046_ rf_ram.memory\[354\]\[1\] _01606_ _01608_ rf_ram.memory\[355\]\[1\] _02240_
+ _02241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_1_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_207_clk clknet_5_24__leaf_clk clknet_leaf_207_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_22_1246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06369__C1 _01636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06908__A1 _02975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_180_3729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09570__A2 _04678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input39_I i_ibus_rdt[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09805_ rf_ram.memory\[75\]\[1\] _04845_ _04847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07997_ rf_ram.memory\[466\]\[1\] _03682_ _03684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06384__A2 _01922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06948_ _03014_ _03026_ _03027_ _00114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09736_ _04781_ net15 _04802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_2_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05373__I _01568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_1180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09667_ _04747_ _04736_ _04750_ _04751_ _01109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_97_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06879_ rf_ram.memory\[301\]\[0\] _02980_ _02981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_94_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06136__A2 _01735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07333__A1 _03055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08618_ rf_ram.memory\[163\]\[1\] _04082_ _04084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09873__A3 _03989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09598_ _04478_ cpu.immdec.imm24_20\[3\] _04700_ _04708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_49_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_171_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_167_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_167_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08549_ rf_ram.memory\[119\]\[0\] _04039_ _04040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_46_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09086__A1 _04367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_166_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_182_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11560_ _01292_ clknet_leaf_112_clk rf_ram.memory\[448\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07636__A2 _03089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10511_ _00255_ clknet_leaf_194_clk rf_ram.memory\[271\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_107_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11491_ _01223_ clknet_leaf_221_clk rf_ram.memory\[503\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_92_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10442_ _00186_ clknet_leaf_221_clk rf_ram.memory\[497\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06932__I _02747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_21_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_1124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_1173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_131_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10373_ _00117_ clknet_leaf_276_clk rf_ram.memory\[231\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_60_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06375__A2 _01989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_1036 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_1231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_66_1627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_103_2311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_68_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_83_1941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_185_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09077__A1 _03668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06328__B _01551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07627__A2 _03452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08824__A1 _04205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10709_ _00453_ clknet_leaf_97_clk rf_ram.memory\[430\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_43_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_181_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_631 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_52_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_70_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_1213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_1273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_178_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_51_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05458__I _01653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07920_ _02983_ _03547_ _03636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09001__A1 _04301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_162_3404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07851_ rf_ram.memory\[410\]\[1\] _03592_ _03594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09552__A2 net44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07563__A1 _03389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06802_ _02801_ _02889_ _02928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07782_ _03524_ _03548_ _03550_ _00425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xinput2 i_dbus_rdt[0] net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05193__I cpu.decode.co_ebreak vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09521_ _03967_ _04648_ _04649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06733_ _02876_ _02874_ _02877_ _00049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_79_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_155_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06118__A2 _01662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09452_ net76 net77 _04593_ _04602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__05326__B1 _01517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06664_ _02779_ _02793_ _02828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_52_1217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08403_ rf_ram.memory\[209\]\[1\] _03936_ _03938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05877__A1 _01768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_19_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05615_ _01635_ _01811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_09383_ _04539_ _04564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__09068__A1 rf_ram.memory\[0\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06595_ _01512_ _01498_ _02773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XTAP_TAPCELL_ROW_177_3680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_176_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05142__B _01344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08334_ rf_ram.memory\[217\]\[1\] _03893_ _03895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07618__A2 _03446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_458 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08009__I _03692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05546_ _01739_ _01741_ _01620_ _01742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08815__A1 net249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_163_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_7_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_49_Left_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_144_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_138_2952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_138_2963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08265_ _03823_ _03849_ _03851_ _00607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_85_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_173_3599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05477_ _01600_ _01639_ _01672_ net253 _01673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_74_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07216_ _02883_ _02941_ _03198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_41_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08196_ _03787_ _03808_ _03809_ _00580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_171_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_162_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_42_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07147_ rf_ram.memory\[497\]\[0\] _03154_ _03155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09240__A1 _04466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05368__I _01563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06054__A1 _01527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09791__A2 _04507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07078_ rf_ram.memory\[492\]\[0\] _03111_ _03112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_125_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06029_ rf_ram.memory\[564\]\[1\] _01538_ _01555_ rf_ram.memory\[565\]\[1\] _01554_
+ rf_ram.memory\[567\]\[1\] _02224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XTAP_TAPCELL_ROW_7_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_58_Left_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_96_1100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06357__A2 _01515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05565__B1 _01668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09719_ _04766_ _04790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__06109__A2 _01634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10991_ _00728_ clknet_leaf_338_clk rf_ram.memory\[163\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_48_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07306__A1 _02899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06927__I _02742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_96_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09059__A1 _04334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_167_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_1075 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11612_ net92 net165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_67_Left_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_61_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08806__A1 rf_ram.memory\[13\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_5_19__f_clk clknet_3_4_0_clk clknet_5_19__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_182_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_167_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_154_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11543_ _01275_ clknet_leaf_53_clk rf_ram.memory\[438\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_25_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_163_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11474_ _01206_ clknet_leaf_202_clk rf_ram.memory\[33\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_123_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_956 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10425_ _00169_ clknet_leaf_208_clk rf_ram.memory\[48\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_61_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10356_ _00100_ clknet_leaf_206_clk rf_ram.memory\[2\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_59_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_76_Left_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_20_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10287_ _00031_ clknet_leaf_122_clk rf_ram.memory\[455\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09534__A2 net38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07545__A1 _03393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06348__A2 _01649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09298__A1 net239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07848__A2 _03559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_85_Left_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_186_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_115_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_185_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_146_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_1250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05400_ cpu.immdec.imm24_20\[3\] _01367_ _01596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_29_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06380_ _01368_ _02547_ _02574_ _01597_ _02575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_29_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_1245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_127_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_155_3274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05331_ _01526_ _01527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_84_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05897__B _01684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08273__A2 _02889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08050_ _03071_ _03693_ _03718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05262_ cpu.decode.op26 _01337_ _01461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_98_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_116_2546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07001_ _03053_ _03059_ _03061_ _00133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_24_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_116_2557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_133_2860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05193_ cpu.decode.co_ebreak _01393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__08025__A2 _03693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_133_2871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_94_Left_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_12_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_45_1065 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_987 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08952_ rf_ram.memory\[121\]\[1\] _04289_ _04291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08499__I _04004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07903_ rf_ram.memory\[444\]\[1\] _03624_ _03626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08883_ rf_ram.memory\[419\]\[0\] _04248_ _04249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07536__A1 _02728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_1318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07834_ rf_ram.memory\[432\]\[1\] _03581_ _03583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_155_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07765_ rf_ram.memory\[394\]\[1\] _03538_ _03540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_179_3720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_155_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11653__I net103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_1150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_149_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06716_ _02826_ _02862_ _02864_ _00045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09504_ _04400_ _04637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_07696_ rf_ram.memory\[382\]\[0\] _03497_ _03498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_177_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_177_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09435_ _01411_ _04593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_78_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06647_ _02814_ _02815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_175_3639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_1178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_23_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_43_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09366_ net205 _04549_ _04552_ net206 _04555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_23_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06578_ _02750_ _02759_ _02760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_129_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08317_ _03855_ _03881_ _03883_ _00627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_152_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05529_ _01714_ _01725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_12
XFILLER_0_90_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09297_ _04466_ _04511_ _04513_ _00977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_133_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08248_ _03820_ _03840_ _03841_ _00600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_105_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_172_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_1111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_921 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08179_ _03798_ _02960_ _03799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__09213__A1 _04434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_162_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06027__A1 _01495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10210_ rf_ram.memory\[442\]\[0\] _05095_ _05096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_127_1188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09764__A2 net25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11190_ _00926_ clknet_leaf_57_clk rf_ram.memory\[90\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10141_ _05049_ _05051_ _05053_ _01282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xoutput180 net180 o_ext_rs2[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__06431__B _01923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput191 net191 o_ext_rs2[29] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__05250__A2 _01382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09516__A2 net57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10072_ _04985_ _05008_ _05010_ _01256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07527__A1 _03389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06750__A2 _02889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_173_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_1137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10974_ _00711_ clknet_leaf_336_clk rf_ram.memory\[170\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_97_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_1272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_167_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_183_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_182_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06266__A1 _01372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11526_ _01258_ clknet_leaf_144_clk rf_ram.memory\[308\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_135_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xwire252 _01734_ net252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_123_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_151_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_68_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_78_1840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_1851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09204__A1 _02805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11457_ _01189_ clknet_leaf_195_clk rf_ram.memory\[263\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_150_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_180_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_68_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10408_ _00152_ clknet_leaf_130_clk rf_ram.memory\[38\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_141_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09755__A2 net21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11388_ _01120_ clknet_leaf_224_clk net102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__07766__A1 _03524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06569__A2 _02752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_111_2454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10339_ _00083_ clknet_leaf_180_clk rf_ram.memory\[285\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_111_2465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_1298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09507__A2 _03083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07518__A1 _03319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05880_ rf_ram.memory\[76\]\[0\] _01755_ _01912_ rf_ram.memory\[77\]\[0\] _02019_
+ rf_ram.memory\[79\]\[0\] _02076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__08191__A1 _03787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1036 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_1069 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07550_ _03393_ _03404_ _03406_ _00337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_157_3303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06501_ cpu.ctrl.pc cpu.ctrl.pc_plus_4_cy_r _02692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_88_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_157_3314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07481_ rf_ram.memory\[328\]\[1\] _03362_ _03364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_76_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09691__A1 _04740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09220_ rf_ram.memory\[349\]\[0\] _04457_ _04458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_29_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06432_ rf_ram.memory\[98\]\[1\] _01785_ _01857_ rf_ram.memory\[99\]\[1\] _01772_
+ rf_ram.memory\[97\]\[1\] _02627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_124_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_173_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_3_2_0_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09151_ _02908_ _04077_ _04415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06363_ _02555_ _02557_ _01494_ _02558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_72_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_161_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_135_2900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_1053 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08246__A2 _02946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_135_2911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_185_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_170_3547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08102_ _03724_ _03748_ _03750_ _00545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05420__B _01615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05314_ _01509_ _01510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_72_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_170_3558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10053__A2 _02894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09082_ net239 _04339_ _04372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_47_1105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06294_ _02487_ _02488_ _01928_ _02489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_86_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_1322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06235__C _01670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08033_ rf_ram.memory\[56\]\[1\] _03706_ _03708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05245_ cpu.bne_or_bge _01443_ _01444_ _01445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_115_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput60 i_ibus_rdt[5] net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_13_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05480__A2 _01543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09746__A2 net18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05176_ _01353_ rf_ram_if.rdata0\[1\] _01377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_101_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07757__A1 _02991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11648__I net129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09984_ rf_ram.memory\[275\]\[1\] _04955_ _04957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_122_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08935_ rf_ram.memory\[399\]\[0\] _04280_ _04281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_36_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_1182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08866_ _04237_ _04235_ _04238_ _00821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input21_I i_dbus_rdt[27] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07817_ rf_ram.memory\[413\]\[0\] _03572_ _03573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_98_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_28_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08797_ _04077_ _04195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_TAPCELL_ROW_28_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07748_ rf_ram.memory\[377\]\[0\] _03529_ _03530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_95_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07679_ _03455_ _03485_ _03486_ _00386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_149_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09682__A1 _04740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_164_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09418_ _04584_ _01027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_109_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10690_ _00434_ clknet_leaf_91_clk rf_ram.memory\[414\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_133_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_137_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09349_ _04545_ _00997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_47_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06426__B _01783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_145_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07101__I _03017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11311_ _01044_ clknet_leaf_266_clk net76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_106_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07996__A1 _03651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_95_2162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_1249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05471__A2 _01666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11242_ _00978_ clknet_leaf_59_clk rf_ram.memory\[66\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_56_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_56_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11173_ _00909_ clknet_leaf_70_clk rf_ram.memory\[97\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06161__B _01693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10124_ _05017_ _05040_ _05042_ _01276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_105_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10055_ _04982_ _04999_ _05000_ _01249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08173__A1 _02881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07920__A1 _02983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10957_ _00007_ clknet_leaf_281_clk rf_ram.regzero vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_57_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10888_ _00632_ clknet_leaf_301_clk rf_ram.memory\[217\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_73_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_152_3211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_155_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_152_3222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_183_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09976__A2 _04951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11509_ _01241_ clknet_leaf_143_clk rf_ram.memory\[326\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_113_2505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_1_clk_I clknet_5_1__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_110_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_1085 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_186_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08400__A2 _02761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_1057 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05466__I _01661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06411__A1 _01909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06981_ _03014_ _03047_ _03048_ _00126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06962__A2 _03009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08720_ rf_ram.memory\[89\]\[0\] _04146_ _04147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05932_ _01350_ _02122_ _02127_ _02128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__08164__A1 _03787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_128_2770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08651_ _04097_ _04102_ _04104_ _00740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05863_ rf_ram.memory\[230\]\[0\] _01940_ _01959_ rf_ram.memory\[231\]\[0\] _01968_
+ rf_ram.memory\[229\]\[0\] _02059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XTAP_TAPCELL_ROW_128_2781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07602_ _03425_ _03436_ _03438_ _00357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08582_ _04058_ _04059_ _04060_ _00715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05794_ rf_ram.memory\[166\]\[0\] _01989_ _01520_ rf_ram.memory\[167\]\[0\] _01516_
+ rf_ram.memory\[165\]\[0\] _01990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_7_1205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_1143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07533_ _03389_ _03395_ _03396_ _00330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_7_1238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_1176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_330_clk_I clknet_5_1__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_77_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_146_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_158_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07464_ _02921_ _02904_ _03352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_146_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_158_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06415_ _02607_ _02609_ _01790_ _02610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_88_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09203_ _04434_ _04445_ _04447_ _00949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_162_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_146_355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07395_ _02765_ _03309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__09416__A1 _04466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09134_ rf_ram.memory\[91\]\[1\] _04403_ _04405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06346_ rf_ram.memory\[198\]\[1\] _01808_ _01805_ _02541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_115_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09065_ net237 _03945_ _04361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06277_ rf_ram.memory\[146\]\[1\] _01958_ _01953_ rf_ram.memory\[147\]\[1\] _02471_
+ _02472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_71_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_103_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08016_ rf_ram.memory\[572\]\[0\] _03697_ _03698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06650__A1 _02743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05228_ _01375_ _01411_ _01428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_103_948 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_1200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_187_3863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_187_3874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_130_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_1244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05159_ _01361_ _01362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_90_2070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_1108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_34_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09967_ rf_ram.memory\[295\]\[1\] _04944_ _04946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_34_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08918_ _04269_ _04267_ _04270_ _00841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08687__I _04057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_51_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08155__A1 _03757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09898_ _04884_ _04902_ _04903_ _01189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08849_ _04205_ _04225_ _04227_ _00815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06166__B1 _01688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_1053 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07902__A1 _03619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_185_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_169_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10811_ _00555_ clknet_leaf_324_clk rf_ram.memory\[551\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_0_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09655__A1 net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_981 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_0_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10742_ _00486_ clknet_leaf_131_clk rf_ram.memory\[43\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_32_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05677__C1 _01811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_165_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_97_2202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_180_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10673_ _00417_ clknet_leaf_109_clk rf_ram.memory\[376\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05141__A1 _01343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_5_18__f_clk_I clknet_3_4_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_11_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_11_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_173_Right_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_36_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05692__A2 _01787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07969__A1 _03651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_775 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08630__A2 _03765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06641__A1 _02748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11225_ _00961_ clknet_leaf_152_clk rf_ram.memory\[329\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_120_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_102_970 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_71_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08394__A1 _03922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11156_ _00892_ clknet_leaf_63_clk rf_ram.memory\[102\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10107_ _05014_ _05031_ _05032_ _01269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_11087_ _00824_ clknet_leaf_295_clk rf_ram.memory\[12\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_179_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08146__A1 _02888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_145_3081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10038_ net248 _02801_ _04990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_145_3092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_153_1310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_106_2364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_106_2375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_147_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09646__A1 _01409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_86_1994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07121__A2 _02911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05668__C1 _01778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06200_ rf_ram.memory\[456\]\[1\] _01724_ _01725_ rf_ram.memory\[457\]\[1\] _01726_
+ rf_ram.memory\[459\]\[1\] _02395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XPHY_EDGE_ROW_140_Right_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_6_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09949__A2 _02815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06880__A1 _02970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07180_ rf_ram.memory\[1\]\[0\] _03175_ _03176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05683__A2 _01845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_30_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_30_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_171_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06131_ _02323_ _02325_ _01746_ _02326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_54_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_2_921 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06632__A1 _02743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06062_ rf_ram.memory\[374\]\[1\] _01662_ _01504_ _02257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_112_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08385__A1 _02959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09821_ _04840_ _04854_ _04856_ _01158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_165_3457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_158_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_182_3771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09752_ _04804_ net20 _04813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_182_3782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06964_ _03014_ _03036_ _03037_ _00120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_126_2729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08703_ _04129_ _04134_ _04136_ _00760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05915_ rf_ram.memory\[121\]\[0\] _01918_ _02111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__06148__B1 _01810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06895_ _02716_ _02811_ _02991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_09683_ net1 net29 _04736_ _04765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08688__A2 _04078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09885__A1 _04887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06699__A1 _02820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09840__B _02714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08634_ _04062_ _04091_ _04093_ _00734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_94_1275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05846_ rf_ram.memory\[192\]\[0\] _01649_ _01650_ _02042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_179_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_77_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09637__A1 _04524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05777_ rf_ram.memory\[134\]\[0\] _01531_ _01973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08565_ _04023_ _04048_ _04049_ _00709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_7_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07516_ rf_ram.memory\[362\]\[1\] _03383_ _03385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_76_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08496_ rf_ram.memory\[359\]\[1\] _04001_ _04003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_30_Left_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_9_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07447_ rf_ram.memory\[331\]\[1\] _03340_ _03342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_64_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_174_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_162_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_284_clk_I clknet_5_18__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_170_clk clknet_5_31__leaf_clk clknet_leaf_170_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_64_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06320__B1 _01911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_1270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_1281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05674__A2 _01724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07378_ rf_ram.memory\[250\]\[1\] _03297_ _03299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_73_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_162_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09117_ _02908_ _03692_ _04393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06329_ rf_ram.memory\[209\]\[1\] _01515_ _02524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_72_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_92_2110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05426__A2 _01614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_299_clk_I clknet_5_7__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09048_ rf_ram.memory\[103\]\[1\] _04349_ _04351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_130_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_20_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output175_I net175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06423__C _01660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11010_ _00747_ clknet_leaf_3_clk rf_ram.memory\[157\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08376__A1 _03919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07179__A2 _02997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10183__A1 _02916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_222_clk_I clknet_5_22__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_1142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_1321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_1275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08128__A1 _03754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09876__A1 _03309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_169_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05898__C1 _01645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09628__A1 _04643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_83_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06665__I _02828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_184_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_67_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08300__A1 _03852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_64_1588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_101_2272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10725_ _00469_ clknet_leaf_119_clk rf_ram.memory\[461\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_32_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_101_2283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_64_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_919 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10656_ _00400_ clknet_leaf_106_clk rf_ram.memory\[380\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_181_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10587_ _00331_ clknet_leaf_164_clk rf_ram.memory\[321\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_140_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08603__A2 _04067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_1000 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_133_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06090__A2 _01709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08367__A1 _03887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_147_3121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_147_3132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11208_ _00944_ clknet_leaf_47_clk rf_ram.memory\[83\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_43_1174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10174__A1 _05046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11139_ _00875_ clknet_leaf_72_clk rf_ram.memory\[111\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_108_2404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08119__A1 _03757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05744__I _01640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09867__A1 _02838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05700_ rf_ram.memory\[412\]\[0\] _01634_ _01702_ rf_ram.memory\[413\]\[0\] _01608_
+ rf_ram.memory\[415\]\[0\] _01896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XTAP_TAPCELL_ROW_160_3365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06680_ _02820_ _02840_ _02841_ _00032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_155_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05631_ rf_ram.memory\[482\]\[0\] _01777_ _01696_ rf_ram.memory\[483\]\[0\] _01826_
+ _01827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_149_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_121_2637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09619__A1 _04643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_121_2648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10229__A2 _02844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08350_ _03884_ _03904_ _03905_ _00638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05562_ rf_ram.memory\[266\]\[0\] _01652_ _01654_ rf_ram.memory\[267\]\[0\] _01715_
+ rf_ram.memory\[265\]\[0\] _01758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_0_59_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07301_ rf_ram.memory\[258\]\[0\] _03250_ _03251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_50_1145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08281_ rf_ram.memory\[194\]\[1\] _03860_ _03862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_152_clk clknet_5_26__leaf_clk clknet_leaf_152_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_05493_ rf_ram.memory\[345\]\[0\] _01626_ _01689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__06302__B1 _01953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07232_ rf_ram.memory\[423\]\[0\] _03207_ _03208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06853__A1 _02930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_1208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05656__A2 _01787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_61_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_132_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07163_ _03161_ _03163_ _03165_ _00191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_119_2599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05408__A2 _01537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06114_ _01527_ _02307_ _02308_ _02309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_07094_ _03087_ _03120_ _03121_ _00166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_124_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_164_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06045_ rf_ram.memory\[353\]\[1\] _01617_ _02240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__06081__A2 _01623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_184_3811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08358__A1 net235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06369__B1 _01610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09804_ _04837_ _04845_ _04846_ _01151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_157_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07996_ _03651_ _03682_ _03683_ _00506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09735_ _04801_ _01127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06947_ rf_ram.memory\[232\]\[0\] _03026_ _03027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_105_Left_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_97_805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_158_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_2_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09666_ net1 net24 _04736_ _04751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06878_ _02935_ _02844_ _02980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08530__A1 _04026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07333__A2 _02917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08617_ _04058_ _04082_ _04083_ _00727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_96_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05829_ _02022_ _02024_ _01978_ _02025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_96_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09597_ _03992_ net47 _04707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_77_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05895__A2 _01711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08548_ net235 _04038_ _04039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_46_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_148_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_148_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_181_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_143_clk clknet_5_27__leaf_clk clknet_leaf_143_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08479_ _03967_ _03992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_64_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10510_ _00254_ clknet_leaf_194_clk rf_ram.memory\[271\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11490_ _01222_ clknet_leaf_181_clk rf_ram.memory\[275\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_165_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10441_ _00185_ clknet_leaf_224_clk rf_ram.memory\[485\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_163_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_162_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_21_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06057__C1 _01646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08597__A1 _04062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_1114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10372_ _00116_ clknet_leaf_276_clk rf_ram.memory\[231\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06072__A2 _01683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_884 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_130_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10156__A1 _05049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_41_clk_I clknet_5_13__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07021__A1 _03050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_176_clk_I clknet_5_30__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_142_3040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09849__A1 _02713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_56_clk_I clknet_5_9__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08521__A1 _03953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_103_2312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_1107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_150_1313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_158_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_87_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_73_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_83_1942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05886__A2 _01537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09077__A2 _02984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_157_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_1230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_134_clk clknet_5_24__leaf_clk clknet_leaf_134_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_83_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05638__A2 _01644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10708_ _00452_ clknet_leaf_101_clk rf_ram.memory\[430\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_114_clk_I clknet_5_15__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_125_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_183_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_102_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10639_ _00383_ clknet_leaf_96_clk rf_ram.memory\[403\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_141_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_148_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_140_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06063__A2 _01536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_129_clk_I clknet_5_13__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05810__A2 _01677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10147__A1 _03672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_18_Right_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_20_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_162_3405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07012__A1 _02738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07850_ _03587_ _03592_ _03593_ _00450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05474__I rf_ram.i_raddr\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08760__A1 _01353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_1034 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06801_ _02819_ _02927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_07781_ rf_ram.memory\[437\]\[1\] _03548_ _03550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_78_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput3 i_dbus_rdt[10] net3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09520_ _01419_ _04647_ _02709_ _04648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_06732_ rf_ram.memory\[518\]\[1\] _02874_ _02877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_116_1219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08512__A1 _01353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06663_ _02826_ _02823_ _02827_ _00029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09451_ _04601_ _01043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_91_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08402_ _03919_ _03936_ _03937_ _00658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05614_ _01714_ _01810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_176_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_87_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06594_ _02748_ _02770_ _02772_ _00015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09382_ _04563_ _01012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_87_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_27_Right_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_177_3681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_164_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_86_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_188_1022 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_74_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07079__A1 _03087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_163_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08333_ _03884_ _03893_ _03894_ _00632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_74_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05545_ rf_ram.memory\[274\]\[0\] _01623_ _01688_ rf_ram.memory\[275\]\[0\] _01740_
+ _01741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
Xclkbuf_leaf_125_clk clknet_5_13__leaf_clk clknet_leaf_125_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_157_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08815__A2 _04195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_163_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06287__C1 _01610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06826__A1 _02930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_138_2953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08264_ rf_ram.memory\[205\]\[1\] _03849_ _03851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05629__A2 _01692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05476_ _01648_ _01659_ _01660_ _01671_ _01672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_116_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_138_2964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_1185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_172_773 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_41_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07215_ _03193_ _03195_ _03197_ _00211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08195_ rf_ram.memory\[538\]\[0\] _03808_ _03809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_41_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07146_ _02761_ _02911_ _03154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_131_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_851 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07251__A1 _02752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07077_ _02788_ _02911_ _03111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_36_Right_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input51_I i_ibus_rdt[26] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06028_ rf_ram.memory\[566\]\[1\] _01532_ _01505_ _02223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_125_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05801__A2 _01664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_113_Left_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06211__C1 _01773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08751__A1 _04129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_87_2020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07979_ _03672_ _02917_ _03673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09718_ _04789_ _01122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_10990_ _00727_ clknet_leaf_339_clk rf_ram.memory\[163\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_48_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07306__A2 _03253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09649_ _04735_ _04736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_167_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_45_Right_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_167_534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06429__B _02004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05333__B _01528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05868__A2 _01683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11611_ net91 net164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_38_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_1162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_116_clk clknet_5_14__leaf_clk clknet_leaf_116_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_33_1173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_122_Left_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_61_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_154_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11542_ _01274_ clknet_leaf_111_clk rf_ram.memory\[373\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_108_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_598 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07490__A1 _03356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06293__A2 _01606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11473_ _01205_ clknet_leaf_202_clk rf_ram.memory\[33\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06164__B _01620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05559__I _01613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10424_ _00168_ clknet_leaf_208_clk rf_ram.memory\[48\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_104_840 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_33_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_54_Right_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06045__A2 _01617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10355_ _00099_ clknet_leaf_178_clk rf_ram.memory\[280\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_59_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10286_ _00030_ clknet_leaf_112_clk rf_ram.memory\[455\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10129__A1 _05017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_131_Left_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_44_1280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05294__I _01409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_63_Right_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09298__A2 _04507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05859__A2 _01664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_150_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_111_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_107_clk clknet_5_15__leaf_clk clknet_leaf_107_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_28_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_127_921 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_1273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06808__A1 _02801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06269__C1 _01953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05330_ _01525_ _01526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_84_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07949__I _03359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_155_3275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_160_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_118_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05261_ cpu.decode.op22 _01460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__06284__A2 _01799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07000_ rf_ram.memory\[225\]\[1\] _03059_ _03061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_25_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_72_Right_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_116_2547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_116_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_142_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05192_ _01391_ net134 _01392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_98_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_109_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_133_2861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_133_2872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07233__A1 _03190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06036__A2 _01544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08981__A1 _04301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08951_ _04266_ _04289_ _04290_ _00854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_161_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05795__A1 _01552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07902_ _03619_ _03624_ _03625_ _00470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08882_ net240 _03547_ _04248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__07536__A2 _03390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07833_ _03554_ _03581_ _03582_ _00444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_81_Right_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_5_25__f_clk clknet_3_6_0_clk clknet_5_25__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07764_ _03521_ _03538_ _03539_ _00418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_179_3710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_179_3721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_1005 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09503_ _04634_ _04635_ _04636_ _01060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06715_ rf_ram.memory\[520\]\[1\] _02862_ _02864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_155_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07695_ _02917_ _03496_ _03497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_56_1173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09434_ _04592_ _01035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06646_ _02736_ _02799_ _02814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_52_1037 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_43_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_23_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09365_ _04554_ _01004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_23_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06577_ _02719_ _02758_ _02759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_47_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08316_ rf_ram.memory\[220\]\[1\] _03881_ _03883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06763__I _02898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05528_ _01643_ _01724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_7_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09296_ rf_ram.memory\[64\]\[1\] _04511_ _04513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_34_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_90_Right_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08247_ rf_ram.memory\[528\]\[0\] _03840_ _03841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06275__A2 _01846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05459_ _01513_ _01655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_62_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_144_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_1101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_160_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08178_ _02845_ _03798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_127_1145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_120_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07129_ rf_ram.memory\[4\]\[1\] _03142_ _03144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_101_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10140_ rf_ram.memory\[453\]\[1\] _05051_ _05053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_28_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06432__C1 _01772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08972__A1 _03071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05786__A1 _01909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput170 net170 o_ext_rs2[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput181 net181 o_ext_rs2[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_98_1218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput192 net192 o_ext_rs2[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_10071_ rf_ram.memory\[508\]\[1\] _05008_ _05010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08724__A1 _02971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05538__A1 _01347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_187_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_337_clk clknet_5_0__leaf_clk clknet_leaf_337_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10973_ _00710_ clknet_leaf_221_clk rf_ram.memory\[509\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_70_1104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_183_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_987 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_773 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07463__A1 _03326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11525_ _01257_ clknet_leaf_145_clk rf_ram.memory\[308\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_135_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11456_ _01188_ clknet_leaf_283_clk rf_ram.memory\[18\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_78_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_150_3172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_78_1852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09204__A2 _03035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_150_3183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07215__A1 _03193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06018__A2 _01511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_1218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10407_ _00151_ clknet_leaf_121_clk rf_ram.memory\[390\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_123_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11387_ _01119_ clknet_leaf_224_clk net101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_81_1255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08963__A1 _04269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10338_ _00082_ clknet_leaf_173_clk rf_ram.memory\[285\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_111_2455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_111_2466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10269_ _00013_ clknet_leaf_282_clk rf_ram.memory\[241\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07518__A2 _02894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_1016 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_178_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06848__I _02959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_187_Right_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_152_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_328_clk clknet_5_4__leaf_clk clknet_leaf_328_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_88_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09140__A1 _04401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06500_ _01376_ _02691_ _01400_ net131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_07480_ _03356_ _03362_ _03363_ _00310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_157_3304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_1100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_88_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_157_3315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_876 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09691__A2 net31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_159_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06431_ rf_ram.memory\[96\]\[1\] _01915_ _01923_ _02626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05701__A1 _01603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06362_ rf_ram.memory\[226\]\[1\] _01958_ _01953_ rf_ram.memory\[227\]\[1\] _02556_
+ _02557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_17_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09150_ _04401_ _04412_ _04414_ _00929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_56_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_135_2901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_1111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_135_2912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08101_ rf_ram.memory\[556\]\[1\] _03748_ _03750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05313_ _01508_ _01509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_12
XTAP_TAPCELL_ROW_170_3548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07454__A1 _02775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_146_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_170_3559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06293_ rf_ram.memory\[138\]\[1\] _01606_ _01608_ rf_ram.memory\[139\]\[1\] _01610_
+ rf_ram.memory\[137\]\[1\] _02488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_09081_ _04367_ _04369_ _04371_ _00903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_142_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05244_ cpu.alu.i_rs1 _01439_ _01342_ _01444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08032_ _03686_ _03706_ _03707_ _00518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_130_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput50 i_ibus_rdt[25] net50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput61 i_ibus_rdt[6] net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_3_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_142_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05175_ _01375_ _01376_ net130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_12_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07757__A2 _03496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08954__A1 _02991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09983_ _04950_ _04955_ _04956_ _01221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08934_ _02953_ _03559_ _04280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_122_1075 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_36_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_36_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08706__A1 _04126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08865_ rf_ram.memory\[409\]\[1\] _04235_ _04238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_99_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11664__I net115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_1235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07816_ _02959_ _03559_ _03572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_165_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08796_ _04170_ _04192_ _04194_ _00795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_28_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input14_I i_dbus_rdt[20] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_28_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07747_ _02983_ _03496_ _03529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_319_clk clknet_5_5__leaf_clk clknet_leaf_319_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_EDGE_ROW_154_Right_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_95_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09131__A1 net244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07678_ rf_ram.memory\[402\]\[0\] _03485_ _03486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_149_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_0_Right_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09417_ net87 net90 _02707_ _04584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07693__A1 _03491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06629_ _02800_ _02801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_48_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_94_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_47_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09348_ net228 _03991_ _04540_ net229 _04545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_30_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09279_ _04501_ _00971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_35_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_1206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11310_ _01043_ clknet_leaf_266_clk net75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_50_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_62_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_95_2163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09198__A1 _04434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_max_cap251_I net252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11241_ _00977_ clknet_leaf_23_clk rf_ram.memory\[64\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_output82_I net82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06442__B _01563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06405__C1 _01656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05759__A1 _01951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11172_ _00908_ clknet_leaf_70_clk rf_ram.memory\[97\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_105_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_140_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_5_0__f_clk_I clknet_3_0_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_73_1760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10123_ rf_ram.memory\[438\]\[1\] _05040_ _05042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06420__A2 _01770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_1026 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_1283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10054_ rf_ram.memory\[34\]\[0\] _04999_ _05000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08173__A2 _02917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06184__A1 _01769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05572__I _01660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07920__A2 _03547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05392__C1 _01554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_121_Right_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10956_ _00694_ clknet_leaf_6_clk rf_ram.memory\[188\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_168_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06487__A2 _01661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10887_ _00631_ clknet_leaf_207_clk rf_ram.memory\[21\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_183_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_152_3212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_171_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_152_3223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07436__A1 _03323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_1318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06239__A2 _01706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_136_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11508_ _01240_ clknet_leaf_169_clk rf_ram.memory\[327\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_80_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_151_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_145_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09189__A1 net242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_130_2820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11439_ _01171_ clknet_leaf_241_clk cpu.mem_bytecnt\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_81_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_123_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08936__A1 _04266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_1059 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_1069 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06980_ rf_ram.memory\[426\]\[0\] _03047_ _03048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_185_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input6_I i_dbus_rdt[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05931_ _02123_ _02124_ _02125_ _02126_ _01978_ _02127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_08650_ rf_ram.memory\[161\]\[1\] _04102_ _04104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_128_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05862_ rf_ram.memory\[228\]\[0\] _01523_ _02058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_128_2782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05482__I _01617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07601_ rf_ram.memory\[354\]\[1\] _03436_ _03438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_117_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05383__C1 _01517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08581_ rf_ram.memory\[168\]\[0\] _04059_ _04060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_89_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05793_ _01640_ _01989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_07532_ rf_ram.memory\[321\]\[0\] _03395_ _03396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_113_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_117_1188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_1079 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_88_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_187_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_76_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07463_ _03326_ _03349_ _03351_ _00305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_146_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09202_ rf_ram.memory\[70\]\[1\] _04445_ _04447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06414_ rf_ram.memory\[114\]\[1\] _01856_ _01857_ rf_ram.memory\[115\]\[1\] _02608_
+ _02609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_173_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07394_ _03292_ _03306_ _03308_ _00279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_134_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09133_ _04397_ _04403_ _04404_ _00922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_115_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06345_ _02538_ _02539_ _01860_ _02540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_127_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08742__B _01506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06276_ rf_ram.memory\[145\]\[1\] _01664_ _02471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_60_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09064_ _04334_ _04358_ _04360_ _00897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05989__A1 net252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05227_ _01426_ _01427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08015_ _02839_ _03693_ _03697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_103_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_38_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_163_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_187_3864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_1148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05158_ _01353_ _01354_ _01355_ _01360_ _01361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_40_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_90_2071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06402__A2 _01785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09966_ _04918_ _04944_ _04945_ _01215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_34_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08968__I _04061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08917_ rf_ram.memory\[439\]\[1\] _04267_ _04270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_51_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09897_ rf_ram.memory\[263\]\[0\] _04902_ _04903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_96_clk clknet_5_14__leaf_clk clknet_leaf_96_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_58_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08848_ rf_ram.memory\[133\]\[1\] _04225_ _04227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_output120_I net120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_1065 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_58_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08779_ _04167_ _04183_ _04184_ _00788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09104__A1 _04364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10810_ _00554_ clknet_leaf_324_clk rf_ram.memory\[551\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_170_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_68_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09655__A2 net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07666__A1 _02866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06469__A2 _01605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10741_ _00485_ clknet_leaf_51_clk rf_ram.memory\[457\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_149_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_165_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05677__B1 _01810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_991 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10672_ _00416_ clknet_leaf_114_clk rf_ram.memory\[376\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_97_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_11_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07418__A1 _02866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_11_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_1026 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_20_clk clknet_5_3__leaf_clk clknet_leaf_20_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_23_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_133_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_1036 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_121_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_75_1800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06172__B _01756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05567__I _01653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08918__A1 _04269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11224_ _00960_ clknet_leaf_152_clk rf_ram.memory\[329\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_102_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_71_1719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11155_ _00891_ clknet_leaf_66_clk rf_ram.memory\[103\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10106_ rf_ram.memory\[312\]\[0\] _05031_ _05032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11086_ _00823_ clknet_leaf_24_clk rf_ram.memory\[130\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08146__A2 _03765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05516__B _01602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10037_ _04985_ _04987_ _04989_ _01242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_145_3082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_145_3093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_187_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_153_1322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05365__C1 _01539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_106_2365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_106_2376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05380__A2 _01502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_86_1995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_169_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_123_2690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10939_ rf_ram_if.rtrig0 clknet_leaf_278_clk rf_ram_if.rtrig1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_151_1090 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05668__B1 _01848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_155_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_39_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_1147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06066__C _01670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05683__A3 _01878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_1115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_11_clk clknet_5_2__leaf_clk clknet_leaf_11_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_182_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_30_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06130_ rf_ram.memory\[298\]\[1\] _01777_ _01778_ rf_ram.memory\[299\]\[1\] _02324_
+ _02325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_26_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_1159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08082__A1 _03724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_121_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06061_ _02254_ _02255_ _01658_ _02256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__08909__A1 _04234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08385__A2 _03903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09820_ rf_ram.memory\[259\]\[1\] _04854_ _04856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_165_3458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09751_ _04812_ _01132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06963_ rf_ram.memory\[22\]\[0\] _03036_ _03037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_182_3772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_78_clk clknet_5_11__leaf_clk clknet_leaf_78_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08702_ rf_ram.memory\[39\]\[1\] _04134_ _04136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05426__B _01615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05914_ rf_ram.memory\[120\]\[0\] _01915_ _01916_ _02110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06148__A1 rf_ram.memory\[312\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09682_ _04740_ _03980_ _04764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06894_ _02975_ _02988_ _02990_ _00097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08633_ rf_ram.memory\[549\]\[1\] _04091_ _04093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_55_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_55_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05845_ rf_ram.memory\[196\]\[0\] _01724_ _01721_ rf_ram.memory\[197\]\[0\] _01713_
+ rf_ram.memory\[199\]\[0\] _02041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XANTENNA__07896__A1 _03619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_1287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_169_Left_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_7_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08564_ rf_ram.memory\[509\]\[0\] _04048_ _04049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05776_ _01615_ _01972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__09637__A2 net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07515_ _03356_ _03383_ _03384_ _00324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07648__A1 _03455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08495_ _03953_ _04001_ _04002_ _00686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_175_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_64_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_36_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_1141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_88_1003 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07446_ _03323_ _03340_ _03341_ _00298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_147_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_107_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07377_ _03289_ _03297_ _03298_ _00272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_134_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_1293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09116_ _04367_ _04390_ _04392_ _00917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_150_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08073__A1 _02761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06328_ rf_ram.memory\[208\]\[1\] _01537_ _01551_ _02523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_92_2100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_178_Left_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_92_2111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07820__A1 _03557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09047_ _04331_ _04349_ _04350_ _00890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06259_ rf_ram.memory\[420\]\[1\] _01666_ _01810_ rf_ram.memory\[421\]\[1\] _01646_
+ rf_ram.memory\[423\]\[1\] _02454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_142_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_130_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10183__A2 _03902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09949_ net248 _02815_ _04935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
Xclkbuf_leaf_69_clk clknet_5_8__leaf_clk clknet_leaf_69_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_102_1287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09325__A1 _04463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09876__A2 _02954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_187_Left_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07887__A1 _03590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_87_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05898__B1 _01646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_1063 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_16_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05362__A2 _01532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_68_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_157_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_0_clk_I clknet_5_1__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10724_ _00468_ clknet_leaf_118_clk rf_ram.memory\[461\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_55_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_101_2273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06311__A1 _02494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_64_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_1079 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10655_ _00399_ clknet_leaf_40_clk rf_ram.memory\[3\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07777__I _03039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08064__A1 _03721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10586_ _00330_ clknet_leaf_164_clk rf_ram.memory\[321\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_140_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07811__A1 net236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05297__I rf_ram.i_raddr\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_146_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_51_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_121_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_1142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_147_3122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_142_1078 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09564__A1 _03992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11207_ _00943_ clknet_leaf_16_clk rf_ram.memory\[179\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_147_3133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06378__A1 _01600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_1216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11138_ _00874_ clknet_leaf_71_clk rf_ram.memory\[111\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_5_6__f_clk clknet_3_1_0_clk clknet_5_6__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_78_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_108_2405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11069_ _00806_ clknet_leaf_15_clk rf_ram.memory\[135\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_0_clk clknet_5_1__leaf_clk clknet_leaf_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09867__A2 _02921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_160_3366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07878__A1 _02916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05630_ rf_ram.memory\[481\]\[0\] _01697_ _01826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__05353__A2 _01523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05760__I _01526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06550__A1 cpu.immdec.imm11_7\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_121_2638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_148_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_121_2649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_176_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05561_ rf_ram.memory\[264\]\[0\] _01755_ _01756_ _01757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_129_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_188_1226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_18_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_73_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07300_ net239 _02941_ _03250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_157_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08280_ _03852_ _03860_ _03861_ _00612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05492_ _01624_ _01688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_46_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07231_ _02829_ _03040_ _03207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_172_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07162_ rf_ram.memory\[496\]\[1\] _03163_ _03165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_81_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_125_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06113_ rf_ram.memory\[268\]\[1\] _01644_ _01645_ rf_ram.memory\[269\]\[1\] _01646_
+ rf_ram.memory\[271\]\[1\] _02308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_0_140_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07093_ rf_ram.memory\[502\]\[0\] _03120_ _03121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_112_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_184_3801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06044_ rf_ram.memory\[352\]\[1\] _01614_ _01615_ _02239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_140_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_565 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_184_3812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08358__A2 _03903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09803_ rf_ram.memory\[75\]\[0\] _04845_ _04846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07995_ rf_ram.memory\[466\]\[0\] _03682_ _03683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09307__A1 _04466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09734_ net110 _04790_ _04791_ net111 _04800_ _04801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_06946_ _02728_ _02766_ _03026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05592__A2 _01787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_1160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_2_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09665_ net123 _04737_ _04749_ _04740_ _04750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_97_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06877_ _02975_ _02977_ _02979_ _00091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_94_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08616_ rf_ram.memory\[163\]\[0\] _04082_ _04083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_94_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_173_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05828_ rf_ram.memory\[210\]\[0\] _01804_ _02019_ rf_ram.memory\[211\]\[0\] _02023_
+ _02024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__06541__A1 _02716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09596_ _04703_ _04704_ _04705_ _04706_ _01083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_82_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08547_ _04037_ _04038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_49_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05759_ _01951_ _01952_ _01954_ _01955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_77_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_46_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_163_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08478_ _03990_ _03991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_119_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_175_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07429_ _02923_ _03101_ _03331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_134_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_169_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_150_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10440_ _00184_ clknet_leaf_224_clk rf_ram.memory\[485\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_21_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06057__B1 _01645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_21_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_1310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_131_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10371_ _00115_ clknet_leaf_276_clk rf_ram.memory\[232\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_33_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_131_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05568__C1 _01668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_142_3030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06780__A1 _02909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05583__A2 _01697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_142_3041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_1244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_66_1618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_103_2313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_1179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_83_1943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05740__C1 _01811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08285__A1 _03852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10092__A1 _05014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10707_ _00451_ clknet_leaf_88_clk rf_ram.memory\[410\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_166_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_1264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08037__A1 _03686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10638_ _00382_ clknet_leaf_97_clk rf_ram.memory\[403\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_52_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09785__A1 _02787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10569_ _00313_ clknet_leaf_172_clk rf_ram.memory\[365\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_24_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_1139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_121_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10147__A2 _02889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06360__B _01956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05755__I _01693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_162_3406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07012__A2 _02917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_283_clk_I clknet_5_18__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06800_ _02876_ _02924_ _02926_ _00067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07780_ _03521_ _03548_ _03549_ _00424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06771__A1 _02881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput4 i_dbus_rdt[11] net4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06731_ _02825_ _02876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_09450_ net75 net76 _04593_ _04601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__05704__B _01629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06662_ rf_ram.memory\[347\]\[1\] _02823_ _02827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05326__A2 _01511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_298_clk_I clknet_5_7__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05490__I _01499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08401_ rf_ram.memory\[209\]\[0\] _03936_ _03937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_118_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05613_ rf_ram.memory\[314\]\[0\] _01808_ _01650_ _01809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_176_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09381_ net212 _04561_ _04552_ net214 _04563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06593_ rf_ram.memory\[233\]\[1\] _02770_ _02772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_177_3682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08332_ rf_ram.memory\[217\]\[0\] _03893_ _03894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_157_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05544_ rf_ram.memory\[273\]\[0\] _01626_ _01740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_35_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_1131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_188_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_leaf_221_clk_I clknet_5_22__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06287__B1 _01636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08263_ _03820_ _03849_ _03850_ _00606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05475_ _01663_ _01665_ _01667_ _01669_ _01670_ _01671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XTAP_TAPCELL_ROW_138_2954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_138_2965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_166_1321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07214_ rf_ram.memory\[261\]\[1\] _03195_ _03197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08194_ _02812_ _02846_ _03808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_41_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_41_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07145_ _03126_ _03151_ _03153_ _00185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_43_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_236_clk_I clknet_5_22__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_30_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07076_ _03092_ _03108_ _03110_ _00159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07251__A2 _02869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11667__I net118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06027_ _01495_ _02216_ _02221_ _02222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_22_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_7_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input44_I i_ibus_rdt[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06211__B1 _01772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_87_2010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09581__B _04678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07978_ _02831_ _03672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_87_2021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06762__A1 _02750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05565__A2 _01509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09717_ net104 _04767_ _04768_ net105 _04788_ _04789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_06929_ _02752_ _02801_ _03015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09700__A1 _04740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09648_ net1 _04734_ _04735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06496__I _01376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06514__A1 _01388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_1000 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_1022 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09579_ _01391_ _01469_ _04646_ _04690_ _04692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_78_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11610_ net90 net163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08267__A1 _03230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_182_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_26_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_61_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_182_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09600__I net48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_61_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11541_ _01273_ clknet_leaf_110_clk rf_ram.memory\[373\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_25_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08019__A1 _03690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11472_ _01204_ clknet_leaf_169_clk rf_ram.memory\[340\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_80_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10423_ _00167_ clknet_leaf_185_clk rf_ram.memory\[502\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_61_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_33_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10354_ _00098_ clknet_leaf_177_clk rf_ram.memory\[280\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_104_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05253__A1 _01385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_59_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10285_ _00029_ clknet_leaf_142_clk rf_ram.memory\[347\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_1101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06180__B _01660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_168_Right_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08742__A2 _04158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05556__A2 _01631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05524__B _01707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06505__A1 _01409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_96_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_1166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_736 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08258__A1 _03820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10065__A1 _04982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06269__B1 _01968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06808__A2 _02894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_155_3265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_155_3276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05260_ _01436_ _01437_ _01459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_126_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_172_3590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_142_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_116_2548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_141_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05191_ _01390_ _01391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_TAPCELL_ROW_116_2559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_148_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_133_2862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_133_2873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08430__A1 _03953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_991 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05244__A1 cpu.alu.i_rs1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_leaf_291_clk clknet_5_18__leaf_clk clknet_leaf_291_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_110_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06441__B1 _01607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_1213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08950_ rf_ram.memory\[121\]\[0\] _04289_ _04290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_110_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_1089 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06992__A1 _03055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07901_ rf_ram.memory\[444\]\[0\] _03624_ _03625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08881_ _04237_ _04245_ _04247_ _00827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_138_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_135_Right_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07832_ rf_ram.memory\[432\]\[0\] _03581_ _03582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05547__A2 _01692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06744__A1 _02873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07763_ rf_ram.memory\[394\]\[0\] _03538_ _03539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_179_3711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09502_ rf_ram.memory\[289\]\[0\] _04635_ _04636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_179_3722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06714_ _02820_ _02862_ _02863_ _00044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08497__A1 _03956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05434__B _01629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_177_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07694_ _03100_ _03496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_09433_ net67 net68 _02707_ _04592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_63_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_78_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_1065 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06645_ _02812_ _02813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_177_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_160_clk_I clknet_5_27__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09364_ net204 _04549_ _04552_ net205 _04554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_43_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06576_ _02756_ _02757_ _02758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XTAP_TAPCELL_ROW_23_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_23_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08315_ _03852_ _03881_ _03882_ _00626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05527_ rf_ram.memory\[330\]\[0\] _01706_ _01602_ _01723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_clkbuf_leaf_40_clk_I clknet_5_7__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09295_ _04463_ _04511_ _04512_ _00976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_117_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08246_ _03798_ _02946_ _03840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_7_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05458_ _01653_ _01654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_12
XFILLER_0_117_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_175_clk_I clknet_5_31__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08177_ _03790_ _03795_ _03797_ _00573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_31_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05389_ rf_ram.memory\[562\]\[0\] _01544_ _01554_ rf_ram.memory\[563\]\[0\] _01555_
+ rf_ram.memory\[561\]\[0\] _01585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_132_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_31_945 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07128_ _03123_ _03142_ _03143_ _00178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_leaf_55_clk_I clknet_5_9__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_1265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_140_1313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_282_clk clknet_5_19__leaf_clk clknet_leaf_282_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__06432__B1 _01857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07059_ _03092_ _03097_ _03099_ _00153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08972__A2 _04303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput160 net160 o_ext_rs1[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__06983__A1 _03018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput171 net171 o_ext_rs2[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput182 net182 o_ext_rs2[20] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput193 net193 o_ext_rs2[30] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_10070_ _04982_ _05008_ _05009_ _01255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_100_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_102_Right_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09921__A1 _04887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_54_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08724__A2 _03945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_113_clk_I clknet_5_15__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_173_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_97_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_1241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_186_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08488__A1 net248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10972_ _00709_ clknet_leaf_221_clk rf_ram.memory\[509\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_138_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07115__I _03134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_128_clk_I clknet_5_13__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10047__A1 _04985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09988__A1 _04950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_65_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06175__B _01504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_1023 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11524_ _01256_ clknet_leaf_198_clk rf_ram.memory\[508\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06266__A3 _02460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11455_ _01187_ clknet_leaf_283_clk rf_ram.memory\[18\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_124_969 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_78_1842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_78_1853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_1201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_150_3173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_123_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_150_3184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_5_31__f_clk clknet_3_7_0_clk clknet_5_31__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10406_ _00150_ clknet_leaf_121_clk rf_ram.memory\[390\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_33_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08412__A1 _03919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_980 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11386_ _01118_ clknet_leaf_224_clk net100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_104_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05226__A1 _01388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_273_clk clknet_5_16__leaf_clk clknet_leaf_273_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10337_ _00081_ clknet_leaf_135_clk rf_ram.memory\[303\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_103_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_111_2456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06974__A1 _02781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05777__A2 _01531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_111_2467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_178_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10268_ _00012_ clknet_leaf_282_clk rf_ram.memory\[241\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09912__A1 _04911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06726__A1 _02826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10199_ _02908_ _03902_ _05089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_108_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_159_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_157_3305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_157_3316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06430_ rf_ram.memory\[100\]\[1\] _01863_ _01848_ rf_ram.memory\[101\]\[1\] _01696_
+ rf_ram.memory\[103\]\[1\] _02625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_159_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06864__I _02819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_174_3630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_173_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_173_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_56_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10038__A1 net248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06361_ rf_ram.memory\[225\]\[1\] _01515_ _02556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_173_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_135_2902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08100_ _03721_ _03748_ _03749_ _00544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05312_ _01496_ _01497_ _01508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_09080_ rf_ram.memory\[57\]\[1\] _04369_ _04371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_170_3549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07454__A2 _02815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08651__A1 _04097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06292_ rf_ram.memory\[136\]\[1\] _01922_ _01923_ _02487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_44_569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08031_ rf_ram.memory\[56\]\[0\] _03706_ _03707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_25_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05243_ cpu.alu.i_rs1 _01439_ _01443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput40 i_ibus_rdt[15] net40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_126_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput51 i_ibus_rdt[26] net51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput62 i_ibus_rdt[7] net62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_130_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05174_ cpu.state.i_ctrl_misalign _01376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_101_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06414__B1 _01857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_264_clk clknet_5_17__leaf_clk clknet_leaf_264_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08954__A2 _04038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09982_ rf_ram.memory\[275\]\[0\] _04955_ _04956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_122_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05768__A2 _01664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08933_ _04269_ _04277_ _04279_ _00847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_23_1140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_36_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09903__A1 _04884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08864_ _04061_ _04237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__06717__A1 _02779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06178__C1 _01668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_58_1214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07815_ _03557_ _03569_ _03571_ _00437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08795_ rf_ram.memory\[139\]\[1\] _04192_ _04194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05925__C1 _01679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_150_Left_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07390__A1 _02752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06193__A2 _01543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_28_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07746_ _03524_ _03526_ _03528_ _00411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_28_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_168_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09131__A2 _04005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07677_ _02923_ _03481_ _03485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_94_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09416_ _04466_ _04581_ _04583_ _01026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_181_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_177_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06628_ _02797_ _02799_ _02800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_177_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10029__A1 _04982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09347_ _04544_ _00996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06559_ _02739_ _02743_ _02744_ _00008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_164_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_1144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09278_ cpu.genblk3.csr.mcause3_0\[1\] _04500_ _04497_ _04501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08642__A1 _02828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08229_ rf_ram.memory\[532\]\[1\] _03828_ _03830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_90_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_95_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_160_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11240_ _00976_ clknet_leaf_23_clk rf_ram.memory\[64\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_132_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09442__I0 net71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10201__A1 _05078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_255_clk clknet_5_20__leaf_clk clknet_leaf_255_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_56_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06405__B1 _01654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05339__B _01506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11171_ _00907_ clknet_leaf_304_clk rf_ram.memory\[569\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_56_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06956__A1 _02766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output75_I net75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10122_ _05014_ _05040_ _05041_ _01275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_73_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_73_1761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_1240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10053_ _02868_ _02894_ _04999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_41_1295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_1061 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_187_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05392__B1 _01555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_775 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10955_ _00693_ clknet_leaf_6_clk rf_ram.memory\[188\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_35_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07133__A1 _03123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06684__I _02843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08881__A1 _04237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06341__C1 _01925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10886_ _00630_ clknet_leaf_208_clk rf_ram.memory\[21\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_112_1223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_1320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_186_1313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_155_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_14_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_14_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_152_3213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_845 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_152_3224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_183_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_171_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11507_ _01239_ clknet_5_30__leaf_clk rf_ram.memory\[327\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_151_530 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_80_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_184_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09189__A2 _04418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11438_ _01170_ clknet_leaf_241_clk cpu.state.o_cnt\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_130_2810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09433__I0 net67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06352__C _01362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_246_clk clknet_5_21__leaf_clk clknet_leaf_246_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_145_1098 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11369_ _01101_ clknet_leaf_218_clk cpu.decode.opcode\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__09436__S _04593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05930_ rf_ram.memory\[98\]\[0\] _01785_ _01857_ rf_ram.memory\[99\]\[0\] _01772_
+ rf_ram.memory\[97\]\[0\] _02126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_119_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05763__I _01695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_178_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05861_ _02054_ _02056_ _01494_ _02057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_179_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_128_2772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07372__A1 _03289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06175__A2 _01662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_128_2783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07600_ _03422_ _03436_ _03437_ _00356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_117_1101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08580_ net250 _03949_ _04059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05792_ rf_ram.memory\[164\]\[0\] _01523_ _01988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05383__B1 _01521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05922__A2 _01641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_1220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10259__A1 _02916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07531_ _03319_ _02899_ _03395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_18_1231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_159_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07462_ rf_ram.memory\[367\]\[1\] _03349_ _03351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05712__B _01907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08872__A1 _02787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09201_ _04431_ _04445_ _04446_ _00948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_147_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05686__A1 _01769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06413_ rf_ram.memory\[113\]\[1\] _01787_ _02608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_29_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_174_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_1218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07393_ rf_ram.memory\[265\]\[1\] _03306_ _03308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_1229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09132_ rf_ram.memory\[91\]\[0\] _04403_ _04404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06344_ rf_ram.memory\[202\]\[1\] _01662_ _01636_ rf_ram.memory\[203\]\[1\] _01645_
+ rf_ram.memory\[201\]\[1\] _02539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XANTENNA__08624__A1 _04062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09063_ rf_ram.memory\[100\]\[1\] _04358_ _04360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_142_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06275_ rf_ram.memory\[144\]\[1\] _01846_ _01956_ _02470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_103_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08014_ _03690_ _03694_ _03696_ _00511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05226_ _01388_ _01425_ _01426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_170_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_38_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_38_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06262__C _01717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_187_3865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09854__B cpu.mem_bytecnt\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05157_ _01357_ _01359_ _01360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__06938__A1 _03014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_1314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_90_2072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09965_ rf_ram.memory\[295\]\[0\] _04944_ _04945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08916_ _04061_ _04269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_51_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09896_ _02828_ _03253_ _04902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_51_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09352__A2 _03991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08847_ _04202_ _04225_ _04226_ _00814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06166__A2 _01623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08778_ rf_ram.memory\[142\]\[0\] _04183_ _04184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_71_1200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_185_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07729_ _03491_ _03515_ _03517_ _00405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_138_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_184_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_68_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_149_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_0_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10740_ _00484_ clknet_leaf_51_clk rf_ram.memory\[457\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08863__A1 _04234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07666__A2 _03089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10671_ _00415_ clknet_leaf_116_clk rf_ram.memory\[395\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_137_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_97_2204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_11_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07418__A2 _03101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08615__A1 _02888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_11_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_146_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_168_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_152_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_23_528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_75_1801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_160_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11223_ _00959_ clknet_leaf_176_clk rf_ram.memory\[339\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_228_clk clknet_5_23__leaf_clk clknet_leaf_228_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_121_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09040__A1 net250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06929__A1 _02752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11154_ _00890_ clknet_leaf_66_clk rf_ram.memory\[103\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_5_27__f_clk_I clknet_3_6_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10105_ _02800_ _02992_ _05031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_11085_ _00822_ clknet_leaf_27_clk rf_ram.memory\[130\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_41_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10036_ rf_ram.memory\[326\]\[1\] _04987_ _04989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_145_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_145_3094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06157__A2 _01683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05365__B1 _01540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_1139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_106_2366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_169_950 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07106__A1 _03123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_175_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_123_2680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_86_1996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_169_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10938_ _00677_ clknet_leaf_259_clk rf_ram.i_raddr\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08854__A1 _04205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_184_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_151_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10869_ _00613_ clknet_leaf_36_clk rf_ram.memory\[194\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_38_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_1213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06363__B _01494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06060_ rf_ram.memory\[378\]\[1\] _01500_ _01763_ rf_ram.memory\[379\]\[1\] _01656_
+ rf_ram.memory\[377\]\[1\] _02255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_1_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_169_3540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_219_clk clknet_5_22__leaf_clk clknet_leaf_219_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__05840__A1 _01972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09582__A2 _04678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07593__A1 _02935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06396__A2 _01770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_165_3459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09750_ net115 _04790_ _04791_ net116 _04811_ _04812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_06962_ _03035_ _03009_ _03036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_20_1121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_182_3773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05913_ _02106_ _02108_ _01790_ _02109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_08701_ _04126_ _04134_ _04135_ _00759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09681_ cpu.bufreg2.o_sh_done_r _04763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06893_ rf_ram.memory\[300\]\[1\] _02988_ _02990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06148__A2 _01666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07345__A1 _03257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08632_ _04058_ _04091_ _04092_ _00733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05844_ rf_ram.memory\[198\]\[0\] _01808_ _01805_ _02040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_90_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08563_ _02915_ _02960_ _04048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05775_ _01955_ _01962_ _01966_ _01970_ _01971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07514_ rf_ram.memory\[362\]\[0\] _03383_ _03384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_76_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08494_ rf_ram.memory\[359\]\[0\] _04001_ _04002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08845__A1 _02794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06257__C _01658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07445_ rf_ram.memory\[331\]\[0\] _03340_ _03341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_9_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_175_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06320__A2 _01856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_135_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_1250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_174_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07376_ rf_ram.memory\[250\]\[0\] _03297_ _03298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_73_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09115_ rf_ram.memory\[93\]\[1\] _04390_ _04392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06327_ _01951_ _02520_ _02521_ _02522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_127_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_162_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08073__A2 _03729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_92_2101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_92_2112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09046_ rf_ram.memory\[103\]\[0\] _04349_ _04350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_115_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06258_ rf_ram.memory\[422\]\[1\] _01940_ _01805_ _02453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_60_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05209_ cpu.state.cnt_r\[1\] cpu.state.cnt_r\[0\] cpu.state.cnt_r\[3\] cpu.state.cnt_r\[2\]
+ _01409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_0_102_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06189_ rf_ram.memory\[472\]\[1\] _01782_ _01783_ _02384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_25_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_99_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_111_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_1144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09948_ _04921_ _04932_ _04934_ _01208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09879_ rf_ram.memory\[239\]\[1\] _04890_ _04892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_5_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_169_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09089__A1 _04364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_68_1660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_16_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_68_1671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05352__B _01505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_165_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10723_ _00467_ clknet_leaf_78_clk rf_ram.memory\[445\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_101_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_181_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_64_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10654_ _00398_ clknet_leaf_40_clk rf_ram.memory\[3\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_125_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_152_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10585_ _00329_ clknet_leaf_160_clk rf_ram.memory\[361\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09261__A1 cpu.mem_bytecnt\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07811__A2 _03234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09013__A1 rf_ram.memory\[10\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11206_ _00942_ clknet_leaf_17_clk rf_ram.memory\[179\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09564__A2 net51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_147_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_147_3134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_1165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07575__A1 _03393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11137_ _00873_ clknet_leaf_75_clk rf_ram.memory\[112\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05527__B _01602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_108_2406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11068_ _00805_ clknet_leaf_13_clk rf_ram.memory\[136\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07327__A1 _03260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_125_2720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10019_ rf_ram.memory\[505\]\[1\] _04976_ _04978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_160_3367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07878__A2 _03234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_121_2639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06550__A2 _02730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_1250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_157_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05560_ _01601_ _01756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_169_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_1223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08827__A1 _04202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_1148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05491_ _01686_ _01687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__06302__A2 _01958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07230_ _03193_ _03204_ _03206_ _00217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_129_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_171_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_171_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07161_ _03157_ _03163_ _03164_ _00190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_27_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05488__I _01550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06112_ rf_ram.memory\[270\]\[1\] _01631_ _02307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07092_ _02915_ _03009_ _03120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_2_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06043_ _01603_ _02236_ _02237_ _02238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_140_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09004__A1 _04298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_184_3802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_184_3813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_160_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_140_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_61_1243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09555__A2 _02709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07566__A1 _02795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06369__A2 _01634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09802_ net246 _04004_ _04845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_10_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07994_ _03672_ _02923_ _03682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07208__I _03017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06945_ _03018_ _03023_ _03025_ _00113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09733_ _04781_ net14 _04800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__07318__A1 _02958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06876_ rf_ram.memory\[282\]\[1\] _02977_ _02979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_2_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09664_ _04737_ _04748_ _04749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_94_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_1074 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_179_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08615_ _02888_ _04067_ _04082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_55_1036 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05827_ rf_ram.memory\[209\]\[0\] _01515_ _02023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_09595_ cpu.immdec.imm24_20\[1\] _04701_ _04706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_167_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05758_ rf_ram.memory\[156\]\[0\] _01614_ _01516_ rf_ram.memory\[157\]\[0\] _01953_
+ rf_ram.memory\[159\]\[0\] _01954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_08546_ _02764_ _02867_ _04037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_148_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_46_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08477_ _01491_ _03989_ net65 _03990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_TAPCELL_ROW_46_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05689_ rf_ram.memory\[394\]\[0\] _01777_ _01778_ rf_ram.memory\[395\]\[0\] _01884_
+ _01885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_49_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09491__A1 cpu.alu.i_rs1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_175_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_148_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07428_ _03326_ _03328_ _03330_ _00291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_64_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05900__B _01707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07359_ rf_ram.memory\[268\]\[0\] _03286_ _03287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_162_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_150_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_21_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_149_Right_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10370_ _00114_ clknet_leaf_276_clk rf_ram.memory\[232\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_66_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_1322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09029_ _04037_ _04339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_40_1305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05568__B1 _01763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_1074 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_142_3031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06780__A2 _02911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_142_3042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_172_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_1159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_103_2303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_1619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_103_2314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06532__A2 _01525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_157_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_139_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08809__A1 net247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_83_1933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05740__B1 _01725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_83_1944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07788__I _03355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06296__A1 _01674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10706_ _00450_ clknet_leaf_88_clk rf_ram.memory\[410\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_113_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_153_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10637_ _00381_ clknet_leaf_91_clk rf_ram.memory\[385\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_102_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_84_1243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10568_ _00312_ clknet_leaf_172_clk rf_ram.memory\[365\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_24_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09785__A2 _04507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_116_Right_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_118_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07796__A1 _02908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_1265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10499_ _00243_ clknet_leaf_200_clk rf_ram.memory\[25\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07548__A1 _03389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_162_3407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09444__S _04593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06771__A2 _02904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06730_ _02873_ _02874_ _02875_ _00048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xinput5 i_dbus_rdt[12] net5 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_127_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_160_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06661_ _02825_ _02826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__07720__A1 _02971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08400_ _03892_ _02761_ _03936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05612_ _01640_ _01808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_09380_ _04562_ _01011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_8_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06592_ _02743_ _02770_ _02771_ _00014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05731__B1 _01925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_177_3672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08331_ _03892_ _02984_ _03893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_74_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_188_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05543_ rf_ram.memory\[272\]\[0\] _01683_ _01615_ _01739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_177_3683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08262_ rf_ram.memory\[205\]\[0\] _03849_ _03850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_6_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05474_ rf_ram.i_raddr\[3\] _01670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_117_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_184_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_138_2955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_138_2966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07213_ _03190_ _03195_ _03196_ _00210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08193_ _03790_ _03805_ _03807_ _00579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_172_775 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_41_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06039__A1 _01351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07144_ rf_ram.memory\[485\]\[1\] _03151_ _03153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_15_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07787__A1 _03524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_18_Left_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_14_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_112_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07075_ rf_ram.memory\[493\]\[1\] _03108_ _03110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05798__B1 _01520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06026_ _02217_ _02218_ _02219_ _02220_ _01495_ _02221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_112_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_1074 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_1085 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_7_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_1062 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08200__A2 _03811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input37_I i_ibus_rdt[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_87_2011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_87_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07977_ _03654_ _03669_ _03671_ _00499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09716_ _04781_ net8 _04788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__06777__I _02908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06928_ _03013_ _03014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XPHY_EDGE_ROW_27_Left_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09700__A2 net3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09647_ _01401_ _04733_ _04734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_179_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06859_ _02822_ _02941_ _02967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_136_1170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09578_ cpu.immdec.imm31 _01419_ _04690_ _04691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_132_1034 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_167_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08529_ rf_ram.memory\[49\]\[1\] _04024_ _04027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_136_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08267__A2 _02795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_61_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11540_ _01272_ clknet_leaf_53_clk rf_ram.memory\[392\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_65_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_92_353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11471_ _01203_ clknet_leaf_169_clk rf_ram.memory\[340\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_52_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_1238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09216__A1 _04431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_36_Left_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_45_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10422_ _00166_ clknet_leaf_185_clk rf_ram.memory\[502\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_116_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07778__A1 _03547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10353_ _00097_ clknet_leaf_137_clk rf_ram.memory\[300\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_103_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_59_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09519__A2 cpu.decode.opcode\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10284_ _00028_ clknet_leaf_142_clk rf_ram.memory\[347\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_45_Left_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05591__I _01514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07702__A1 _03488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_1075 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_150_1123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_155_3266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_155_3277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_54_Left_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07311__I _03013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_181_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_114_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_172_3580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11669_ net121 net193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_71_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_172_3591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_153_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_98_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_116_2549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05190_ cpu.branch_op _01390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_153_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_1036 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07769__A1 _03521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_1182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_133_2863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_133_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06992__A2 _02894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07900_ _02839_ _03547_ _03624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_20_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08880_ rf_ram.memory\[128\]\[1\] _04245_ _04247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08194__A1 _02812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_63_Left_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07831_ _02945_ _03234_ _03581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_138_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06597__I net247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07762_ _02775_ _03481_ _03538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_159_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_179_3712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09501_ _03445_ _02899_ _04635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_179_3723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_155_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06713_ rf_ram.memory\[520\]\[0\] _02862_ _02863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07693_ _03491_ _03493_ _03495_ _00391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_56_1142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_91_1022 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09694__A1 _04740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09432_ _04591_ _01034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06644_ _02773_ _02811_ _02812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_52_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_149_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09363_ _04553_ _01003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_47_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06575_ _01562_ _02717_ _02757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_59_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_164_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_23_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_23_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_72_Left_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05526_ rf_ram.memory\[332\]\[0\] _01709_ _01721_ rf_ram.memory\[333\]\[0\] _01713_
+ rf_ram.memory\[335\]\[0\] _01722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_08314_ rf_ram.memory\[220\]\[0\] _03881_ _03882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09294_ rf_ram.memory\[64\]\[0\] _04511_ _04512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_28_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08245_ _03823_ _03837_ _03839_ _00599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_90_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05457_ _01518_ _01653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_160_701 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09857__B _02690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06680__A1 _02820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_172_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08176_ rf_ram.memory\[542\]\[1\] _03795_ _03797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_43_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_1114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05388_ rf_ram.memory\[560\]\[0\] _01511_ _01552_ _01584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_104_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07127_ rf_ram.memory\[4\]\[0\] _03142_ _03143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_179_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_140_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07058_ rf_ram.memory\[38\]\[1\] _03097_ _03099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput150 net150 o_ext_rs1[20] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput161 net161 o_ext_rs1[30] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_06009_ _02200_ _02201_ _02202_ _02203_ _01494_ _02204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XPHY_EDGE_ROW_81_Left_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xoutput172 net172 o_ext_rs2[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__09592__B _01491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput183 net183 o_ext_rs2[21] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput194 net194 o_ext_rs2[31] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_100_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_54_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07932__A1 _03619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05625__B _01684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05943__B1 _01624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08488__A2 _03496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10971_ _00708_ clknet_leaf_185_clk rf_ram.memory\[499\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_69_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06499__A1 _01375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_845 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_1248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05171__A1 _01368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_183_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06456__B _01562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11408__CLK clknet_5_28__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_282_clk_I clknet_5_19__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11523_ _01255_ clknet_leaf_211_clk rf_ram.memory\[508\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_68_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_163_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06671__A1 _02820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11454_ _01186_ clknet_leaf_298_clk rf_ram.memory\[219\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_68_1079 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_78_1843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_78_1854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_150_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10405_ _00149_ clknet_leaf_118_clk rf_ram.memory\[391\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_151_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_150_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11385_ _01117_ clknet_leaf_219_clk net99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__05586__I _01682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_297_clk_I clknet_5_7__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10336_ _00080_ clknet_leaf_135_clk rf_ram.memory\[303\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_111_2457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06974__A2 _03040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_111_2468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10267_ _00011_ clknet_leaf_37_clk rf_ram.memory\[201\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09912__A2 _02992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_220_clk_I clknet_5_22__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10198_ _05081_ _05086_ _05088_ _01304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06187__B1 _01778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_1321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_159_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_235_clk_I clknet_5_22__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_157_3306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_157_3317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05162__A1 cpu.genblk3.csr.o_new_irq vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_174_3620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_174_3631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10038__A2 _02801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06360_ rf_ram.memory\[224\]\[1\] _01846_ _01956_ _02555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_56_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09979__A2 _04951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08100__A1 _03721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07041__I _03013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05311_ rf_ram.memory\[526\]\[0\] _01502_ _01506_ _01507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_135_2903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06291_ _01909_ _02484_ _02485_ _02486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_72_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08030_ _03668_ _02992_ _03706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_86_1146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_114_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_154_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05242_ cpu.decode.co_mem_word _01442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_86_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_140_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput30 i_dbus_rdt[6] net30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_114_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput41 i_ibus_rdt[16] net41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_142_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput52 i_ibus_rdt[27] net52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput63 i_ibus_rdt[8] net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_4_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_114_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05173_ net138 _01375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__05496__I _01682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05217__A2 cpu.mem_bytecnt\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09981_ _02865_ _02958_ _04955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_08932_ rf_ram.memory\[123\]\[1\] _04277_ _04279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08167__A1 _03790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_36_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08863_ _04234_ _04235_ _04236_ _00820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06178__B1 _01763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07914__A1 _03622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07814_ rf_ram.memory\[434\]\[1\] _03569_ _03571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08794_ _04167_ _04192_ _04193_ _00794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05925__B1 _01793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07390__A2 _03253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_58_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07745_ rf_ram.memory\[396\]\[1\] _03526_ _03528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07676_ _03458_ _03482_ _03484_ _00385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09415_ rf_ram.memory\[299\]\[1\] _04581_ _04583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06627_ _02798_ cpu.immdec.imm11_7\[4\] _02730_ _02799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_164_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_1281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09346_ net227 _03991_ _04540_ net228 _04544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_75_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06558_ rf_ram.memory\[200\]\[0\] _02739_ _02744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_47_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_164_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05509_ _01681_ _01691_ _01700_ _01704_ _01705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_09277_ _01365_ _01392_ _04499_ _04500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_06489_ _01348_ _02678_ _02683_ _02684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__06102__B1 _01625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08642__A2 _02881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_160_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08228_ _03820_ _03828_ _03829_ _00592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_31_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_95_2165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08159_ rf_ram.memory\[545\]\[1\] _03784_ _03786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09442__I1 net72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_981 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11170_ _00906_ clknet_leaf_305_clk rf_ram.memory\[569\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_56_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_56_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_144_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_1096 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_1133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10121_ rf_ram.memory\[438\]\[0\] _05040_ _05041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06956__A2 _02806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_1253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_179_1310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_73_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_max_cap237_I _02903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_73_1762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08158__A1 _03754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10052_ _04985_ _04996_ _04998_ _01248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07905__A1 _02787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05916__B1 _01911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_1073 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_1050 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_39_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10954_ _00692_ clknet_leaf_3_clk rf_ram.memory\[172\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_74_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10885_ _00629_ clknet_leaf_215_clk rf_ram.memory\[242\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06341__B1 _01912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_191_clk clknet_5_28__leaf_clk clknet_leaf_191_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_39_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_128_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05695__A2 _01846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06892__A1 _02970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_152_3214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_152_3225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_170_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06644__A1 _02773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11506_ _01238_ clknet_leaf_212_clk rf_ram.memory\[246\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_124_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05852__C1 _01959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11437_ _01169_ clknet_leaf_239_clk cpu.ctrl.i_jump vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_124_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_130_2811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08397__A1 _03919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_1039 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_120_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11368_ _01100_ clknet_5_20__leaf_clk cpu.decode.opcode\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_22_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_1196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10319_ _00063_ clknet_leaf_211_clk rf_ram.memory\[511\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11299_ _01032_ clknet_leaf_251_clk net94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_167_3490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05860_ rf_ram.memory\[226\]\[0\] _01958_ _01953_ rf_ram.memory\[227\]\[0\] _02055_
+ _02056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XTAP_TAPCELL_ROW_128_2773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09452__S _04593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_174_clk_I clknet_5_31__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05791_ _01351_ _01971_ _01986_ _01362_ _01987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_07530_ _03393_ _03391_ _03394_ _00329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_135_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10259__A2 _03692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_54_clk_I clknet_5_9__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08321__A1 _03884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07461_ _03323_ _03349_ _03350_ _00304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_147_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05712__C net254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_1313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_182_clk clknet_5_29__leaf_clk clknet_leaf_182_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08872__A2 _03945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_186_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_159_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06412_ rf_ram.memory\[112\]\[1\] _01915_ _01916_ _02607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_29_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09200_ rf_ram.memory\[70\]\[0\] _04445_ _04446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06883__A1 _02750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_189_clk_I clknet_5_29__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07392_ _03289_ _03306_ _03307_ _00278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_174_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_72_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06343_ rf_ram.memory\[200\]\[1\] _01915_ _01916_ _02538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09131_ net244 _04005_ _04403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_127_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_69_clk_I clknet_5_8__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09821__A1 _04840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06635__A1 _02773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09062_ _04331_ _04358_ _04359_ _00896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_115_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06274_ _02466_ _02468_ _01564_ _02469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_154_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_112_clk_I clknet_5_15__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_5_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_170_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05225_ _01398_ _01424_ _01425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08013_ rf_ram.memory\[573\]\[1\] _03694_ _03696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_114_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_38_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_38_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05156_ _01337_ _01358_ _01359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_69_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_187_3866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_1258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_90_2062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_127_clk_I clknet_5_13__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07060__A1 _02764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09964_ _03445_ _02829_ _04944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_90_2073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05610__A2 _01804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08915_ _04266_ _04267_ _04268_ _00840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08330__I _02737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09888__A1 _04884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09895_ _04887_ _04899_ _04901_ _01188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_51_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08846_ rf_ram.memory\[133\]\[0\] _04225_ _04226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06020__C1 _01517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08560__A1 _04023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05374__A1 _01351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08777_ _02971_ _04152_ _04183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05989_ net252 _02157_ _02184_ _02185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_95_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07728_ rf_ram.memory\[37\]\[1\] _03515_ _03517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_95_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08312__A1 _03855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07659_ rf_ram.memory\[404\]\[1\] _03472_ _03474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_173_clk clknet_5_31__leaf_clk clknet_leaf_173_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_0_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_149_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_177_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05677__A2 _01666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10670_ _00414_ clknet_leaf_116_clk rf_ram.memory\[395\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_63_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_97_2205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09329_ rf_ram.memory\[309\]\[0\] _04533_ _04534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_11_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_146_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_164_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08615__A2 _04067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09812__A1 _02828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06087__C1 _01715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_75_1802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_161_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08379__A1 _03922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11222_ _00958_ clknet_leaf_176_clk rf_ram.memory\[339\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_31_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09040__A2 _04339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06929__A2 _02801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11153_ _00889_ clknet_leaf_68_clk rf_ram.memory\[104\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10104_ _05017_ _05028_ _05030_ _01268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05601__A2 _01719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11084_ _00821_ clknet_leaf_88_clk rf_ram.memory\[409\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_41_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10035_ _04982_ _04987_ _04988_ _01241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_76_1101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_145_3084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_145_3095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06011__C1 _01554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_19_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_106_2367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08303__A1 _03230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_86_1997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_123_2681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05532__C _01658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10110__A1 net250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10937_ cpu.o_wdata0 clknet_leaf_261_clk rf_ram_if.wdata0_r\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_14_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_164_clk clknet_5_27__leaf_clk clknet_leaf_164_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_129_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_184_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05668__A2 _01863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06865__A1 _02773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10868_ _00612_ clknet_leaf_36_clk rf_ram.memory\[194\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_144_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_26_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_1140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_171_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_5_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_171_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10799_ _00543_ clknet_leaf_333_clk rf_ram.memory\[557\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_147_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_53_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_30_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06617__A1 _02743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_30_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07290__A1 _02836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_169_3530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_169_3541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10177__A1 _03892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07042__A1 _02830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07593__A2 _02822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06250__C1 _01857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09319__C2 cpu.immdec.imm11_7\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_33_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06961_ _02996_ _03035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_182_3774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08700_ rf_ram.memory\[39\]\[0\] _04134_ _04135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05912_ rf_ram.memory\[114\]\[0\] _01856_ _01857_ rf_ram.memory\[115\]\[0\] _02107_
+ _02108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_09680_ _04762_ _01111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06892_ _02970_ _02988_ _02989_ _00096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_94_1223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06002__C1 _01539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08631_ rf_ram.memory\[549\]\[0\] _04091_ _04092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_179_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05843_ _02037_ _02038_ _01860_ _02039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_77_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08562_ _04026_ _04045_ _04047_ _00708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_178_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05774_ _01951_ _01967_ _01969_ _01970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_49_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07513_ _02775_ _03101_ _03383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_18_1051 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_155_clk clknet_5_26__leaf_clk clknet_leaf_155_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08493_ _02829_ _03496_ _04001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_65_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08845__A2 _04195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06856__A1 _02927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05659__A2 _01782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07444_ _02781_ _02815_ _03340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_91_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_1165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_57_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_31_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07375_ _03055_ _02813_ _03297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_146_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_1273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06608__A1 _02743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09114_ _04364_ _04390_ _04391_ _00916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_161_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06326_ rf_ram.memory\[214\]\[1\] _01804_ _02019_ rf_ram.memory\[215\]\[1\] _01968_
+ rf_ram.memory\[213\]\[1\] _02521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_0_72_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06257_ _02448_ _02449_ _02450_ _02451_ _01658_ _02452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XANTENNA__06084__A2 _01706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_92_2102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09045_ _02828_ _04339_ _04349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_32_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_92_2113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05208_ _01399_ _01407_ _01408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_128_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05831__A2 _01515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06188_ _02380_ _02382_ _01790_ _02383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_41_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07033__A1 _03053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05139_ cpu.csr_d_sel _01342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_187_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09156__I _04004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08781__A1 _04170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_70_1710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09947_ rf_ram.memory\[338\]\[1\] _04932_ _04934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_141_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05617__C _01658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_1313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09878_ _04884_ _04890_ _04891_ _01181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08533__A1 _04023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08829_ _04205_ _04213_ _04215_ _00807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05898__A2 _01801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_16_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_68_1661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_68_1672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_146_clk clknet_5_26__leaf_clk clknet_leaf_146_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_67_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_166_921 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10722_ _00466_ clknet_leaf_78_clk rf_ram.memory\[445\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_32_1037 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06847__A1 _02750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_738 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_165_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_101_2275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10653_ _00397_ clknet_leaf_107_clk rf_ram.memory\[381\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_153_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_180_423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10584_ _00328_ clknet_leaf_160_clk rf_ram.memory\[361\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09261__A2 _01385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_1182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_146_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_181_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_161_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06480__C1 _01653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05822__A2 _01523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_1280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10159__A1 _05046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_1058 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07024__A1 _02738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11205_ _00941_ clknet_leaf_49_clk rf_ram.memory\[84\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_147_3124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05594__I _01493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08772__A1 _02953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06232__C1 _01763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11136_ _00872_ clknet_leaf_75_clk rf_ram.memory\[112\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_108_2407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11067_ _00804_ clknet_leaf_12_clk rf_ram.memory\[136\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_125_2710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_125_2721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10018_ _04950_ _04976_ _04977_ _01235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_160_3357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_188_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_160_3368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05543__B _01615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_175_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_137_clk clknet_5_26__leaf_clk clknet_leaf_137_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_47_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_156_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06838__A1 _02930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05490_ _01499_ _01686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_184_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_1071 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07160_ rf_ram.memory\[496\]\[0\] _03163_ _03164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_54_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_172_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06093__C _01658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06111_ _02294_ _02298_ _02302_ _02305_ _02306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_70_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07263__A1 _02738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07091_ _03092_ _03117_ _03119_ _00165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_140_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06042_ rf_ram.memory\[358\]\[1\] _01606_ _01608_ rf_ram.memory\[359\]\[1\] _01610_
+ rf_ram.memory\[357\]\[1\] _02237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_23_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_184_3803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_184_3814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07566__A2 _03390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09801_ _04840_ _04842_ _04844_ _01150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_22_1239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07993_ _03654_ _03679_ _03681_ _00505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_158_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09732_ _04799_ _01126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06944_ rf_ram.memory\[206\]\[1\] _03023_ _03025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07318__A2 _02946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_1065 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09663_ net120 _03975_ _04748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06875_ _02970_ _02977_ _02978_ _00090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_2_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_179_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_2_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_1184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08614_ _04062_ _04079_ _04081_ _00726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05826_ rf_ram.memory\[208\]\[0\] _01537_ _01551_ _02022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_10_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09594_ _04526_ net46 _04705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_55_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08545_ _04026_ _04034_ _04036_ _00702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_89_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05757_ _01695_ _01953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
Xclkbuf_leaf_128_clk clknet_5_13__leaf_clk clknet_leaf_128_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_49_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06829__A1 _02935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08476_ _02695_ _03989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_77_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05688_ rf_ram.memory\[393\]\[0\] _01697_ _01884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_46_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07427_ rf_ram.memory\[333\]\[1\] _03328_ _03330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_63_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_1070 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_45_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_73_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_165_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_163_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07358_ _02788_ _03253_ _03286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_32_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_162_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06057__A2 _01666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_21_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06309_ rf_ram.memory\[172\]\[1\] _01683_ _01516_ rf_ram.memory\[173\]\[1\] _01953_
+ rf_ram.memory\[175\]\[1\] _02504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XTAP_TAPCELL_ROW_21_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_300_clk clknet_5_7__leaf_clk clknet_leaf_300_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07289_ _03225_ _03241_ _03243_ _00239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_115_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05804__A2 _01501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09028_ _04334_ _04336_ _04338_ _00883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_130_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output173_I net173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07006__A1 _03053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05628__B _01746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_1105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08506__A1 cpu.immdec.imm11_7\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_142_3032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_1213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06459__B _01525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_1115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_103_2304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_103_2315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_158_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_119_clk clknet_5_12__leaf_clk clknet_leaf_119_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_83_1934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08809__A2 _04195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_83_1945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_185_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10705_ _00449_ clknet_leaf_99_clk rf_ram.memory\[431\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_113_1171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07493__A1 _02788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05589__I _01686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10636_ _00380_ clknet_leaf_92_clk rf_ram.memory\[385\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_102_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_187_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_64_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_181_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_10_1165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07245__A1 _03193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06048__A2 _01614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10567_ _00311_ clknet_leaf_151_clk rf_ram.memory\[328\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_118_2580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_101_Left_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_118_2591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_1217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07796__A2 _03559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_1108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_1239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10498_ _00242_ clknet_leaf_199_clk rf_ram.memory\[25\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_5_14__f_clk clknet_3_3_0_clk clknet_5_14__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_121_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08745__A1 _01495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06205__C1 _01810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_9_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_1120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_162_3408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_5_11__f_clk_I clknet_3_2_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11119_ _00855_ clknet_leaf_84_clk rf_ram.memory\[121\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_120_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_78_1059 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput6 i_dbus_rdt[13] net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06660_ _02747_ _02825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_188_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06088__C _01717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05611_ rf_ram.memory\[316\]\[0\] _01724_ _01725_ rf_ram.memory\[317\]\[0\] _01726_
+ rf_ram.memory\[319\]\[0\] _01807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_118_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06591_ rf_ram.memory\[233\]\[0\] _02770_ _02771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_176_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_1166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_143_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08330_ _02737_ _03892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_177_3673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05542_ _01675_ _01736_ _01737_ _01738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_177_3684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05473_ rf_ram.memory\[370\]\[0\] _01500_ _01519_ rf_ram.memory\[371\]\[0\] _01668_
+ rf_ram.memory\[369\]\[0\] _01669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_08261_ _03230_ _02844_ _03849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06287__A2 _01662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_1098 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_138_2956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05499__I _01518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_138_2967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07212_ rf_ram.memory\[261\]\[0\] _03195_ _03196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_61_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08192_ rf_ram.memory\[53\]\[1\] _03805_ _03807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_55_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_132_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_41_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07236__A1 _02806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07143_ _03123_ _03151_ _03152_ _00184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_42_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08984__A1 _04298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07074_ _03087_ _03108_ _03109_ _00158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_140_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06025_ rf_ram.memory\[546\]\[1\] _01544_ _01521_ rf_ram.memory\[547\]\[1\] _01517_
+ rf_ram.memory\[545\]\[1\] _02220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_140_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08736__A1 _02713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_7_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_1074 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_1104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06211__A2 _01711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07976_ rf_ram.memory\[46\]\[1\] _03669_ _03671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_87_2012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_87_2023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09715_ _04787_ _01121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06927_ _02742_ _03013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__09161__A1 _04401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09646_ _01409_ _04731_ _04732_ _04733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_06858_ _02930_ _02964_ _02966_ _00085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_182_Right_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_167_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05809_ rf_ram.memory\[190\]\[0\] _01641_ _02004_ _02005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09577_ _01399_ _01469_ cpu.decode.opcode\[1\] _04690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06789_ rf_ram.memory\[510\]\[0\] _02918_ _02919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_78_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08528_ _03689_ _04026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_72_1181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_182_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_1165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_182_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_61_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08459_ net120 net123 _03975_ _03976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_65_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_14_Right_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_18_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11470_ _01202_ clknet_leaf_170_clk rf_ram.memory\[341\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_34_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05202__I cpu.state.stage_two_req vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10421_ _00165_ clknet_leaf_183_clk rf_ram.memory\[490\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_61_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_150_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07778__A2 _03072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output98_I net98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10352_ _00096_ clknet_leaf_137_clk rf_ram.memory\[300\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_61_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06461__C rf_ram.i_raddr\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10283_ _00027_ clknet_leaf_141_clk rf_ram.memory\[346\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_131_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_1272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_178_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_23_Right_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06202__A2 _01804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06968__I _03039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05961__A1 _01599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06189__B _01783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_158_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_32_Right_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_29_738 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06269__A2 _01614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07466__A1 _03323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_166_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_154_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_1249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_155_3267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_155_3278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11668_ net119 net191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_181_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_172_3581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_172_3592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_52_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07218__A1 _03190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10619_ _00363_ clknet_leaf_154_clk rf_ram.memory\[313\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_135_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11599_ _01329_ clknet_leaf_306_clk rf_ram.memory\[574\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_98_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_1003 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_133_2864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_133_2875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_1058 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06441__A2 _01605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_1069 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_41_Right_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08718__A1 _04129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08194__A2 _02846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07830_ _03557_ _03578_ _03580_ _00443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05782__I _01493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07761_ _03524_ _03535_ _03537_ _00417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_155_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09143__A1 _04397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09500_ _04396_ _04634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_06712_ _02728_ _02846_ _02862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_179_3713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_1132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_179_3724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07692_ rf_ram.memory\[401\]\[1\] _03493_ _03495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_155_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_149_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_177_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09431_ net96 net67 _02707_ _04591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06643_ _02719_ _02810_ _02811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_188_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_78_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_50_Right_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09362_ net203 _04549_ _04552_ net204 _04553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06574_ _02720_ _02722_ _02756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XTAP_TAPCELL_ROW_43_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_118_913 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_23_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08313_ _03230_ _02839_ _03881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_23_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05525_ _01714_ _01721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_12
X_09293_ net237 _04507_ _04511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_7_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08244_ rf_ram.memory\[52\]\[1\] _03837_ _03839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_62_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05456_ _01499_ _01652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_133_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09857__C _01391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_160_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_7_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08175_ _03787_ _03795_ _03796_ _00572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_31_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05387_ rf_ram.memory\[564\]\[0\] _01538_ _01555_ rf_ram.memory\[565\]\[0\] _01554_
+ rf_ram.memory\[567\]\[0\] _01583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_15_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_1114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07126_ _02883_ _02997_ _03142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_141_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07057_ _03087_ _03097_ _03098_ _00152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06432__A2 _01785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput140 net140 o_ext_rs1[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_112_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput151 net151 o_ext_rs1[21] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__08709__A1 net235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput162 net162 o_ext_rs1[31] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_06008_ rf_ram.memory\[530\]\[1\] _01501_ _01554_ rf_ram.memory\[531\]\[1\] _01555_
+ rf_ram.memory\[529\]\[1\] _02203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_11_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput173 net173 o_ext_rs2[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput184 net184 o_ext_rs2[22] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput195 net195 o_ext_rs2[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__06196__A1 _02379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_54_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_173_1102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_138_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output136_I net136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07959_ _03651_ _03659_ _03660_ _00492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_74_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10970_ _00707_ clknet_leaf_185_clk rf_ram.memory\[499\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09629_ _04524_ net55 _04723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06499__A2 _02690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05171__A2 _01371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_127_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07448__A1 _03326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_148_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_50_clk clknet_5_12__leaf_clk clknet_leaf_50_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_11522_ _01254_ clknet_leaf_151_clk rf_ram.memory\[307\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_109_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_163_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_163_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_136_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11453_ _01185_ clknet_leaf_298_clk rf_ram.memory\[219\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_123_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_1301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08948__A1 _04269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09339__I _04539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_78_1844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10404_ _00148_ clknet_leaf_118_clk rf_ram.memory\[391\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_184_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_150_3175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_1855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11384_ _01116_ clknet_leaf_218_clk net129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_150_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_150_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_1247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10335_ _00079_ clknet_leaf_175_clk rf_ram.memory\[286\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_131_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_1092 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_111_2458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05631__B1 _01696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10266_ _00010_ clknet_leaf_37_clk rf_ram.memory\[201\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05816__B _01923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10197_ rf_ram.memory\[210\]\[1\] _05086_ _05088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09074__I _04061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_157_3307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_157_3318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05551__B _01746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_115_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_185_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_174_3621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_174_3632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_158_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07439__A1 _02921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_173_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_41_clk clknet_5_13__leaf_clk clknet_leaf_41_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_05310_ _01505_ _01506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_86_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_135_2904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06290_ rf_ram.memory\[140\]\[1\] _01799_ _01931_ rf_ram.memory\[141\]\[1\] _01857_
+ rf_ram.memory\[143\]\[1\] _02485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_140_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_141_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_1109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05241_ _01343_ _01440_ _01441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput20 i_dbus_rdt[26] net20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_25_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput31 i_dbus_rdt[7] net31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_25_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput42 i_ibus_rdt[17] net42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_114_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08939__A1 net245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput53 i_ibus_rdt[28] net53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_130_919 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput64 i_ibus_rdt[9] net64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05172_ _01351_ _01362_ _01374_ _00007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_80_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_969 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_123_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06414__A2 _01856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05217__A3 _01385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09980_ _04953_ _04951_ _04954_ _01220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_40_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08931_ _04266_ _04277_ _04278_ _00846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_58_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08862_ rf_ram.memory\[409\]\[0\] _04235_ _04236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_36_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07813_ _03554_ _03569_ _03570_ _00436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_58_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08793_ rf_ram.memory\[139\]\[0\] _04192_ _04193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09116__A1 _04367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07744_ _03521_ _03526_ _03527_ _00410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_95_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07675_ rf_ram.memory\[384\]\[1\] _03482_ _03484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_95_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05689__B1 _01778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_66_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09414_ _04463_ _04581_ _04582_ _01025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06626_ cpu.immdec.imm11_7\[3\] _02798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__05153__A2 _01343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09345_ _04543_ _00995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_164_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06557_ _02742_ _02743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_48_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_32_clk clknet_5_6__leaf_clk clknet_leaf_32_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_05508_ _01603_ _01701_ _01703_ _01704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09276_ _01364_ cpu.genblk3.csr.mcause3_0\[2\] _04499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06488_ _02679_ _02680_ _02681_ _02682_ rf_ram.i_raddr\[3\] _02683_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_118_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08227_ rf_ram.memory\[532\]\[0\] _03828_ _03829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_117_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07850__A1 _03587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05439_ _01518_ _01635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_172_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06292__B _01923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_95_2155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_880 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_95_2166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08158_ _03754_ _03784_ _03785_ _00566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_30_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07109_ _02728_ _02911_ _03131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07602__A1 _03425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06405__A2 _01652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_1101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08089_ rf_ram.memory\[558\]\[0\] _03742_ _03743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_56_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_113_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_56_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_113_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10120_ _03008_ _03547_ _05040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_179_1322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_73_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_73_1763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_99_clk clknet_5_14__leaf_clk clknet_leaf_99_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10051_ rf_ram.memory\[306\]\[1\] _04996_ _04998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07905__A2 _02832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09107__A1 _02916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05392__A2 _01538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_1040 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10953_ _00691_ clknet_leaf_4_clk rf_ram.memory\[172\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06467__B _01601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_97_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_168_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_167_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10884_ _00628_ clknet_leaf_215_clk rf_ram.memory\[242\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_78_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_182_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_1322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_183_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_600 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_23_clk clknet_5_3__leaf_clk clknet_leaf_23_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_14_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_152_3215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_14_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_152_3226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11505_ _01237_ clknet_leaf_213_clk rf_ram.memory\[246\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_41_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05597__I _01617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05852__B1 _01968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11436_ _01168_ clknet_leaf_242_clk cpu.state.cnt_r\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_110_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_46_1131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_130_2812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09594__A1 _04526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11367_ _01099_ clknet_leaf_235_clk cpu.csr_d_sel vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_104_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10318_ _00062_ clknet_leaf_211_clk rf_ram.memory\[511\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_120_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11298_ _01031_ clknet_leaf_251_clk net93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__09346__A1 net227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_167_3491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10249_ _02838_ _03035_ _05119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05546__B _01620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_128_2774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05790_ _01975_ _01979_ _01982_ _01985_ _01349_ _01986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__05383__A2 _01544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_159_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_88_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07460_ rf_ram.memory\[367\]\[0\] _03349_ _03350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_186_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_174_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_14_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_186_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06411_ _01909_ _02604_ _02605_ _02606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_07391_ rf_ram.memory\[265\]\[0\] _03306_ _03307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_146_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_14_clk clknet_5_2__leaf_clk clknet_leaf_14_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09130_ _04401_ _04398_ _04402_ _00921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_151_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08085__A1 _03721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06342_ _01972_ _02535_ _02536_ _02537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_127_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_154_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09061_ rf_ram.memory\[100\]\[0\] _04358_ _04359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06273_ rf_ram.memory\[154\]\[1\] _01958_ _01959_ rf_ram.memory\[155\]\[1\] _02467_
+ _02468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_127_595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08012_ _03686_ _03694_ _03695_ _00510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05224_ _01412_ _01383_ _01423_ _01424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_130_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_170_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_38_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_1204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05155_ cpu.decode.op26 cpu.decode.co_ebreak _01358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_38_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_187_3867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09963_ _04921_ _04941_ _04943_ _01214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_4_Right_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_110_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07060__A2 _02799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_90_2063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_90_2074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09337__A1 _04466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08914_ rf_ram.memory\[439\]\[0\] _04267_ _04268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_110_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09894_ rf_ram.memory\[18\]\[1\] _04899_ _04901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_40_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_51_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07899__A1 _03622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_51_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08845_ _02794_ _04195_ _04225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_58_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_281_clk_I clknet_5_19__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06020__B1 _01521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08776_ _04170_ _04180_ _04182_ _00787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06571__A1 _02743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05988_ _01349_ _02172_ _02183_ net254 _02184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_169_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input12_I i_dbus_rdt[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07727_ _03488_ _03515_ _03516_ _00404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_149_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07658_ _03455_ _03472_ _03473_ _00378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_0_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06323__A1 _01768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_296_clk_I clknet_5_7__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_0_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_164_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06609_ rf_ram.memory\[235\]\[1\] _02782_ _02784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_76_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07589_ rf_ram.memory\[355\]\[0\] _03430_ _03431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05531__C1 _01726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07897__I _03359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09328_ _03445_ _03072_ _04533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_36_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_97_2206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_11_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09812__A2 _03035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06087__B1 _01654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_1078 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07823__A1 _03554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09259_ cpu.genblk3.csr.mie_mtie _04486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_63_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_146_1321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_1218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11221_ _00957_ clknet_leaf_176_clk rf_ram.memory\[349\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_121_738 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output80_I net80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_1040 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11152_ _00888_ clknet_leaf_68_clk rf_ram.memory\[104\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05598__C1 _01793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09328__A1 _03445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10103_ rf_ram.memory\[311\]\[1\] _05028_ _05030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_101_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11083_ _00820_ clknet_leaf_89_clk rf_ram.memory\[409\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_41_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10034_ rf_ram.memory\[326\]\[0\] _04987_ _04988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_249_clk_I clknet_5_21__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_145_3085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_175_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06011__B1 _01555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_145_3096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_188_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05365__A2 _01544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05813__C _01860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_106_2368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06197__B _01707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08303__A2 _02960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10936_ net259 clknet_leaf_261_clk rf_ram_if.wdata0_r\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_86_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_123_2682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_86_1998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10110__A2 _03088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_1231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10867_ _00611_ clknet_leaf_46_clk rf_ram.memory\[195\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_85_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_183_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_1139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_94_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10798_ _00542_ clknet_leaf_333_clk rf_ram.memory\[557\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_109_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_155_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_1107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06078__B1 _01696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_1196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_1128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07290__A2 _03135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_169_3531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11419_ _01151_ clknet_leaf_24_clk rf_ram.memory\[75\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_112_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10177__A2 _02775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07042__A2 _02939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_1140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09319__A1 _04526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06250__B1 _01931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09319__B2 cpu.immdec.imm11_7\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06960_ _03018_ _03032_ _03034_ _00119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_33_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_3_clk clknet_5_1__leaf_clk clknet_leaf_3_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_33_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07047__I _03017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_129_Left_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_182_3764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_183_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09463__S _04604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input4_I i_dbus_rdt[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05911_ rf_ram.memory\[113\]\[0\] _01787_ _02107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_182_3775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06891_ rf_ram.memory\[300\]\[0\] _02988_ _02989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06002__B1 _01540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08630_ _02794_ _03765_ _04091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_05842_ rf_ram.memory\[202\]\[0\] _01662_ _01636_ rf_ram.memory\[203\]\[0\] _01645_
+ rf_ram.memory\[201\]\[0\] _02038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XANTENNA__06553__A1 _02728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08561_ rf_ram.memory\[499\]\[1\] _04045_ _04047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05773_ rf_ram.memory\[150\]\[0\] _01958_ _01953_ rf_ram.memory\[151\]\[0\] _01968_
+ rf_ram.memory\[149\]\[0\] _01969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_7_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07512_ _03360_ _03380_ _03382_ _00323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_76_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08492_ _03956_ _03998_ _04000_ _00685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_76_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_174_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_146_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07443_ _03326_ _03337_ _03339_ _00297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_169_1310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_146_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_138_Left_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_119_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_175_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_174_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08058__A1 _03721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07374_ _03292_ _03294_ _03296_ _00271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_174_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09113_ rf_ram.memory\[93\]\[0\] _04390_ _04391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_31_1285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06325_ rf_ram.memory\[212\]\[1\] _01510_ _02520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07805__A1 _03557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09044_ _04334_ _04346_ _04348_ _00889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06256_ rf_ram.memory\[424\]\[1\] _01666_ _01810_ rf_ram.memory\[425\]\[1\] _01811_
+ rf_ram.memory\[427\]\[1\] _02451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_60_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_92_2103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_92_2114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05292__A1 cpu.alu.i_rs1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05207_ _01390_ _01382_ _01405_ _01406_ _01407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_25_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06187_ rf_ram.memory\[466\]\[1\] _01777_ _01778_ rf_ram.memory\[467\]\[1\] _02381_
+ _02382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_64_1061 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_1072 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05138_ cpu.state.genblk1.misalign_trap_sync_r cpu.genblk3.csr.o_new_irq _01340_
+ _01341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_40_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08230__A1 _03823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_1102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_147_Left_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_141_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_70_1700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_1213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09946_ _04918_ _04932_ _04933_ _01207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06792__A1 _02876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09877_ rf_ram.memory\[239\]\[0\] _04890_ _04891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09730__A1 _04781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05914__B _01916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08828_ rf_ram.memory\[135\]\[1\] _04213_ _04215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06544__A1 _01347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_79_Right_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08759_ _01363_ _01366_ _04172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_output216_I net216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_68_1662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_16_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_68_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08297__A1 _03855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_156_Left_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_165_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10721_ _00465_ clknet_leaf_120_clk rf_ram.memory\[462\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_32_1027 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_101_2276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08049__A1 _03690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10652_ _00396_ clknet_leaf_107_clk rf_ram.memory\[381\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_165_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_48_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09797__A1 net245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_183_1318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10583_ _00327_ clknet_leaf_163_clk rf_ram.memory\[322\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_8_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09261__A3 cpu.decode.co_ebreak vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_88_Right_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_134_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_173_clk_I clknet_5_31__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_146_1173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06480__B1 _01655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_165_Left_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_clkbuf_leaf_53_clk_I clknet_5_12__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_1292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11204_ _00940_ clknet_leaf_49_clk rf_ram.memory\[84\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08221__A1 _03798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07024__A2 _02813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_147_3125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06232__B1 _01668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11135_ _00871_ clknet_5_10__leaf_clk rf_ram.memory\[113\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08772__A2 _04152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_188_clk_I clknet_5_29__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11066_ _00803_ clknet_leaf_11_clk rf_ram.memory\[137\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_108_2408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_68_clk_I clknet_5_8__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09721__A1 _04781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_97_Right_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10017_ rf_ram.memory\[505\]\[0\] _04976_ _04977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_125_2711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_125_2722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_160_3358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_160_3369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_111_clk_I clknet_5_15__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_188_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_174_Left_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_176_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08288__A1 _03230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_157_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10095__A1 _02814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10919_ _00663_ clknet_leaf_16_clk rf_ram.memory\[177\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_39_460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_126_clk_I clknet_5_13__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_172_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_143_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_41_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_172_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06110_ _01603_ _02303_ _02304_ _02305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_42_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07263__A2 _02883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07090_ rf_ram.memory\[490\]\[1\] _03117_ _03119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_152_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_183_Left_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_70_989 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06041_ rf_ram.memory\[356\]\[1\] _01537_ _02236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_152_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_184_3804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_140_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_112_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_184_3815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09800_ rf_ram.memory\[58\]\[1\] _04842_ _04844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_22_1229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07992_ rf_ram.memory\[477\]\[1\] _03679_ _03681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_5_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_163_Right_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06943_ _03014_ _03023_ _03024_ _00112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09731_ net108 _04790_ _04791_ net110 _04798_ _04799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_09662_ net120 _04747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_94_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06874_ rf_ram.memory\[282\]\[0\] _02977_ _02978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_101_1290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_2_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_2_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08613_ rf_ram.memory\[129\]\[1\] _04079_ _04081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05825_ _01951_ _02018_ _02020_ _02021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09593_ _04477_ cpu.immdec.imm24_20\[2\] _04704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_94_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08544_ rf_ram.memory\[171\]\[1\] _04034_ _04036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05756_ rf_ram.memory\[158\]\[0\] _01501_ _01952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09720__I _04760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_148_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06829__A2 _02946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08475_ _01436_ _03988_ _00680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_77_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05687_ rf_ram.memory\[392\]\[0\] _01782_ _01693_ _01883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_46_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07426_ _03323_ _03328_ _03329_ _00290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_175_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_162_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_63_1570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09779__A1 _04637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07357_ _03260_ _03283_ _03285_ _00265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_33_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_162_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06308_ rf_ram.memory\[174\]\[1\] _01501_ _02503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08451__A1 _02714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_21_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07288_ rf_ram.memory\[471\]\[1\] _03241_ _03243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_61_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09027_ rf_ram.memory\[107\]\[1\] _04336_ _04338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06239_ rf_ram.memory\[438\]\[1\] _01706_ _01911_ rf_ram.memory\[439\]\[1\] _01931_
+ rf_ram.memory\[437\]\[1\] _02434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_130_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08203__A1 _03790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09400__B1 _04564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10010__A1 _04953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09951__A1 _04918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05568__A2 _01500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09929_ _04911_ _03072_ _04923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_130_Right_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08506__A2 cpu.immdec.imm11_7\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09703__A1 _04740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_142_3033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06517__A1 _02703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_172_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_1236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_103_2305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_103_2316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_157_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05740__A2 _01724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_83_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10077__A1 _04985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_83_1946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_120_2630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_166_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10704_ _00448_ clknet_leaf_99_clk rf_ram.memory\[431\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_165_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07493__A2 _03101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_166_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08690__A1 _04126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_165_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_153_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_187_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_37_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_1280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10635_ _00379_ clknet_leaf_114_clk rf_ram.memory\[404\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_153_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_126_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_181_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_1223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10566_ _00310_ clknet_leaf_157_clk rf_ram.memory\[328\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_52_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_118_2581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_118_2592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10497_ _00241_ clknet_leaf_53_clk rf_ram.memory\[468\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_121_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06205__B1 _01811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_9_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_162_3409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11118_ _00854_ clknet_leaf_84_clk rf_ram.memory\[121\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_120_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11049_ _00786_ clknet_leaf_10_clk rf_ram.memory\[143\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput7 i_dbus_rdt[14] net7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07181__A1 _03157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_1050 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05610_ rf_ram.memory\[318\]\[0\] _01804_ _01805_ _01806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_188_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06590_ _02752_ _02766_ _02770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_87_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_176_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05731__A2 _01719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_146_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_87_875 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10068__A1 _02838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05541_ rf_ram.memory\[278\]\[0\] _01687_ _01679_ rf_ram.memory\[279\]\[0\] _01678_
+ rf_ram.memory\[277\]\[0\] _01737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_0_188_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_177_3674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_177_3685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08260_ _03823_ _03846_ _03848_ _00605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_15_1066 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_184_560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08681__A1 _04097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05472_ _01655_ _01668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__06141__C1 _01713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07211_ _02795_ _02941_ _03195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_166_1313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_138_2957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_138_2968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08191_ _03787_ _03805_ _03806_ _00578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_55_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_89_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07142_ rf_ram.memory\[485\]\[0\] _03151_ _03152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07236__A2 _03040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08433__A1 _03956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09481__I0 net89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_294_clk clknet_5_7__leaf_clk clknet_leaf_294_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07073_ rf_ram.memory\[493\]\[0\] _03108_ _03109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_164_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05798__A2 _01958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06024_ rf_ram.memory\[544\]\[1\] _01524_ _01528_ _02219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_11_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_112_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_1162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09933__A1 _04921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07975_ _03651_ _03669_ _03670_ _00498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_87_2013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_87_2024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09714_ net103 _04767_ _04768_ net104 _04786_ _04787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_06926_ _02975_ _03010_ _03012_ _00107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05970__A2 _01514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06857_ rf_ram.memory\[284\]\[1\] _02964_ _02966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09645_ cpu.mem_bytecnt\[1\] _01376_ _01375_ _01385_ _04732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_69_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05808_ _01504_ _02004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_171_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_139_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09576_ _04689_ _01080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_65_1610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06788_ _02915_ _02917_ _02918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_78_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08527_ _04023_ _04024_ _04025_ _00695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_77_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05739_ rf_ram.memory\[430\]\[0\] _01804_ _01805_ _01935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_33_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_78_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_5_20__f_clk clknet_3_5_0_clk clknet_5_20__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_148_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08458_ _03973_ _03974_ _03975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_61_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08672__A1 _02838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_175_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07409_ rf_ram.memory\[372\]\[1\] _03316_ _03318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_136_958 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08389_ _03922_ _03927_ _03929_ _00653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_46_783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10420_ _00164_ clknet_leaf_183_clk rf_ram.memory\[490\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_123_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08424__A1 _03919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05238__A1 net134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_285_clk clknet_5_18__leaf_clk clknet_leaf_285_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__10231__A1 _05078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10351_ _00095_ clknet_leaf_180_clk rf_ram.memory\[281\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_115_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10282_ _00026_ clknet_leaf_141_clk rf_ram.memory\[346\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_130_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_1104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_1284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06738__A1 _02876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_5_3__f_clk_I clknet_3_0_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05946__C1 _01609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09561__S _04678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07163__A1 _03161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06984__I _03013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06371__C1 _01702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_115_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_185_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_96_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_1233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_25_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_1277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_166_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05477__A1 _01600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_155_3268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_155_3279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_127_969 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11667_ net118 net190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_126_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_172_3582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_172_3593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_141_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10618_ _00362_ clknet_leaf_105_clk rf_ram.memory\[313\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_153_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09463__I0 net81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11598_ _00001_ clknet_leaf_281_clk rf_ram.rdata\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_107_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05229__A1 cpu.alu.i_rs1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_109_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_276_clk clknet_5_16__leaf_clk clknet_leaf_276_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_51_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10549_ _00293_ clknet_leaf_149_clk rf_ram.memory\[370\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_24_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_133_2865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_121_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05401__A1 _01369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07760_ rf_ram.memory\[376\]\[1\] _03535_ _03537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09471__S _04604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05952__A2 _01613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06711_ _02826_ _02859_ _02861_ _00043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_2_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_179_3714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07691_ _03488_ _03493_ _03494_ _00390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_179_3725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09430_ _04590_ _01033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_200_clk clknet_5_25__leaf_clk clknet_leaf_200_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_06642_ _02756_ _02724_ _02810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__05165__B1 _01367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06901__A1 _02975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_1128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09361_ _04539_ _04552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_177_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06573_ _02748_ _02753_ _02755_ _00011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_43_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08312_ _03855_ _03878_ _03880_ _00625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05524_ rf_ram.memory\[334\]\[0\] _01719_ _01707_ _01720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_23_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08654__A1 _04094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09292_ _04466_ _04508_ _04510_ _00975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_118_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_878 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08243_ _03820_ _03837_ _03838_ _00598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05455_ rf_ram.memory\[376\]\[0\] _01649_ _01650_ _01651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_7_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08174_ rf_ram.memory\[542\]\[0\] _03795_ _03796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05386_ rf_ram.memory\[566\]\[0\] _01532_ _01505_ _01582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09454__I0 net77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_1240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_127_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_160_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_267_clk clknet_5_17__leaf_clk clknet_leaf_267_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07125_ _03126_ _03139_ _03141_ _00177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10213__A1 _05081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_70_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07056_ rf_ram.memory\[38\]\[0\] _03097_ _03098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_141_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput130 net130 o_dbus_sel[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput141 net141 o_ext_rs1[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__09906__A1 _03445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput152 net152 o_ext_rs1[22] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__08709__A2 _04078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06007_ rf_ram.memory\[528\]\[1\] _01511_ _01552_ _02202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_58_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput163 net163 o_ext_rs1[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput174 net174 o_ext_rs2[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_10_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input42_I i_ibus_rdt[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput185 net185 o_ext_rs2[23] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput196 net196 o_ext_rs2[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__05906__C _01362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05928__C1 _01696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_54_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07958_ rf_ram.memory\[480\]\[0\] _03659_ _03660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05943__A2 _01605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06909_ _02822_ _02997_ _03001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07889_ rf_ram.memory\[445\]\[0\] _03616_ _03617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_output129_I net129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07145__A1 _03126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09628_ _04643_ _01447_ _04663_ _01099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05922__B _02004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09559_ _01491_ _04676_ _04677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_78_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05171__A3 _01372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11521_ _01253_ clknet_leaf_150_clk rf_ram.memory\[307\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_19_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_110_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06120__A2 _01644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_184_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11452_ _01184_ clknet_leaf_281_clk rf_ram.memory\[229\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_135_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_258_clk clknet_5_17__leaf_clk clknet_leaf_258_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__10204__A1 _03892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10403_ _00147_ clknet_leaf_301_clk rf_ram.memory\[215\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_78_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_151_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11383_ _01115_ clknet_5_23__leaf_clk net128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_78_1856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_115_2540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_150_3176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_150_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_81_1237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10334_ _00078_ clknet_leaf_174_clk rf_ram.memory\[286\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_81_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_111_2459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10265_ _00009_ clknet_leaf_33_clk rf_ram.memory\[200\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05919__C1 _01786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10196_ _05078_ _05086_ _05087_ _01303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07384__A1 _03292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06187__A2 _01777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05934__A2 _01530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07136__A1 _02915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08884__A1 _04234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06344__C1 _01645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_157_3308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_157_3319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_174_3622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_146_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_174_3633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08636__A1 _02893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07439__A2 _02883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_135_2905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_182_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_154_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05240_ _01430_ _01431_ _01439_ _01440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
Xinput10 i_dbus_rdt[17] net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput21 i_dbus_rdt[27] net21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_71_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput32 i_dbus_rdt[8] net32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_142_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput43 i_ibus_rdt[18] net43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08939__A2 _04038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_249_clk clknet_5_21__leaf_clk clknet_leaf_249_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xinput54 i_ibus_rdt[29] net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_109_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_24_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05171_ _01368_ _01371_ _01372_ _01373_ _01374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
Xinput65 i_rst net65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_40_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08930_ rf_ram.memory\[123\]\[0\] _04277_ _04278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_149_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_1290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05793__I _01640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_36_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08861_ _02983_ _03559_ _04235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_36_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07375__A1 _03055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06178__A2 _01500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07812_ rf_ram.memory\[434\]\[0\] _03569_ _03570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08792_ net246 _04152_ _04192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_74_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05925__A2 _01863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_1239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07743_ rf_ram.memory\[396\]\[0\] _03526_ _03527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07127__A1 rf_ram.memory\[4\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07674_ _03455_ _03482_ _03483_ _00384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08609__I _04077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06625_ _02796_ _02763_ _02797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_09413_ rf_ram.memory\[299\]\[0\] _04581_ _04582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_149_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_845 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06556_ _02741_ _02742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__08627__A1 _04058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09344_ net224 _03991_ _04540_ net227 _04543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_168_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05507_ rf_ram.memory\[342\]\[0\] _01623_ _01688_ rf_ram.memory\[343\]\[0\] _01702_
+ rf_ram.memory\[341\]\[0\] _01703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_09275_ _04498_ _00970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_8_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06487_ rf_ram.memory\[2\]\[1\] _01661_ _01635_ rf_ram.memory\[3\]\[1\] _01714_ rf_ram.memory\[1\]\[1\]
+ _02682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XANTENNA__06102__A2 _01623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08226_ _03798_ _03135_ _03828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05438_ _01633_ _01634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_160_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09427__I0 net94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_160_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08157_ rf_ram.memory\[545\]\[0\] _03784_ _03785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_95_2156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05369_ _01558_ _01559_ _01560_ _01561_ _01564_ _01565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_TAPCELL_ROW_95_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09052__A1 _04331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07108_ _03126_ _03128_ _03130_ _00171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_114_983 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_1065 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08088_ _02971_ _03729_ _03742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_101_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_56_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07039_ rf_ram.memory\[215\]\[1\] _03084_ _03086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05917__B _01928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_1210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_1232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_73_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_140_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_73_1764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10050_ _04982_ _04996_ _04997_ _01247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07366__A1 _03289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06169__A2 _01631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_1287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05916__A2 _01706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09107__A2 _04005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07118__A1 _03123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_1075 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_27_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08866__A1 _04237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10952_ _00690_ clknet_leaf_259_clk rf_ram_if.wen0_r vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06326__C1 _01968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_1183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10883_ _00627_ clknet_leaf_31_clk rf_ram.memory\[220\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_97_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06341__A2 _01649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_14_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_152_3216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_152_3227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_163_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11504_ _01236_ clknet_leaf_198_clk rf_ram.memory\[505\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_80_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11435_ _01167_ clknet_leaf_242_clk cpu.state.cnt_r\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_123_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_130_2802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_130_2813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09594__A2 net46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11366_ _01098_ clknet_leaf_235_clk cpu.decode.co_mem_word vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_105_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_10_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10317_ _00061_ clknet_leaf_268_clk rf_ram.memory\[512\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11297_ _01030_ clknet_leaf_252_clk net92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__09346__A2 _03991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10248_ _02825_ _05116_ _05118_ _01324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_167_3492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07357__A1 _03260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10179_ _05046_ _05075_ _05076_ _01297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05907__A2 _01510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_128_2775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07109__A1 _02728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08857__A1 _04202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_1234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_1283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06377__C _01860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_1147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_1070 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_1278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06332__A2 _01537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06410_ rf_ram.memory\[118\]\[1\] _01856_ _01911_ rf_ram.memory\[119\]\[1\] _01931_
+ rf_ram.memory\[117\]\[1\] _02605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_18_1289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07390_ _02752_ _03253_ _03306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_85_984 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06341_ rf_ram.memory\[204\]\[1\] _01649_ _01912_ rf_ram.memory\[205\]\[1\] _01925_
+ rf_ram.memory\[207\]\[1\] _02536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_44_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06096__A1 _01368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09060_ net241 _04339_ _04358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_115_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06272_ rf_ram.memory\[153\]\[1\] _01515_ _02467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_72_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08011_ rf_ram.memory\[573\]\[0\] _03694_ _03695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_72_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05223_ _01421_ _01422_ _01383_ _01423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_53_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09034__A1 _04334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_130_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_38_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05154_ _01347_ _01356_ _01357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_38_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_1216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_187_3857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06399__A2 _01683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_187_3868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09962_ rf_ram.memory\[335\]\[1\] _04941_ _04943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_40_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_90_2064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_90_2075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08913_ _03039_ _03083_ _04267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_09893_ _04884_ _04899_ _04900_ _01187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07348__A1 _02813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_51_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08844_ _04205_ _04222_ _04224_ _00813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_51_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08775_ rf_ram.memory\[143\]\[1\] _04180_ _04182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05987_ _01348_ _02177_ _02182_ _02183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_07726_ rf_ram.memory\[37\]\[0\] _03515_ _03516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_178_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_174_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_177_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07657_ rf_ram.memory\[404\]\[0\] _03472_ _03473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_67_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07520__A1 _03356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_177_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06608_ _02743_ _02782_ _02783_ _00018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_94_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07588_ _02889_ _03390_ _03430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05531__B1 _01725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06539_ _02723_ _02724_ _02725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XTAP_TAPCELL_ROW_97_2207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09327_ _04466_ _04530_ _04532_ _00988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_11_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_168_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_11_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_146_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09258_ _04480_ _04482_ _04483_ _04485_ _00966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_TAPCELL_ROW_32_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_91_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08209_ _03798_ _03083_ _03817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_62_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09189_ net242 _04418_ _04439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_121_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_177_Right_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_11220_ _00956_ clknet_leaf_192_clk rf_ram.memory\[349\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_105_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07587__A1 _03425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_max_cap242_I _02865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11151_ _00887_ clknet_leaf_68_clk rf_ram.memory\[105\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05598__B1 _01778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output73_I net73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10102_ _05014_ _05028_ _05029_ _01267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09328__A2 _03072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11082_ _00819_ clknet_leaf_28_clk rf_ram.memory\[131\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10033_ _02805_ _02815_ _04987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_179_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_145_3086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_145_3097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05382__B _01528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_106_2358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08839__A1 _04205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_106_2369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_169_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_98_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10935_ cpu.o_wdata1 clknet_leaf_261_clk rf_ram_if.wdata1_r\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_86_1988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_123_2683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06314__A2 _01989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_86_1999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_151_1061 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_183_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10866_ _00610_ clknet_leaf_46_clk rf_ram.memory\[195\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_67_984 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_995 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10797_ _00541_ clknet_leaf_319_clk rf_ram.memory\[558\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_112_1089 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_186_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_53_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05825__A1 _01951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09016__A1 _04301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_144_Right_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_2_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11418_ _01150_ clknet_leaf_287_clk rf_ram.memory\[58\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_169_3532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11349_ _01081_ clknet_leaf_254_clk cpu.immdec.imm30_25\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_22_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09319__A2 net35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_33_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_33_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_182_3765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05910_ rf_ram.memory\[112\]\[0\] _01915_ _01916_ _02106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_182_3776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06890_ _02788_ _02801_ _02988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_146_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05841_ rf_ram.memory\[200\]\[0\] _01915_ _01916_ _02037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06553__A2 _02738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06388__B _01551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05772_ _01918_ _01968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_08560_ _04023_ _04045_ _04046_ _00707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07511_ rf_ram.memory\[323\]\[1\] _03380_ _03382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_76_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_187_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08491_ rf_ram.memory\[369\]\[1\] _03998_ _04000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_18_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_187_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_1053 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07502__A1 _03360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06305__A2 _01664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_5_1__f_clk clknet_3_0_0_clk clknet_5_1__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_76_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07442_ rf_ram.memory\[36\]\[1\] _03337_ _03339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_18_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_1322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07373_ rf_ram.memory\[267\]\[1\] _03294_ _03296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06324_ net251 _02491_ _02518_ _02519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_73_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09112_ _02959_ _04005_ _04390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_143_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09043_ rf_ram.memory\[104\]\[1\] _04346_ _04348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06255_ rf_ram.memory\[426\]\[1\] _01808_ _01650_ _02450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_115_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09007__A1 _02971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_875 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_92_2104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_309_clk_I clknet_5_5__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_92_2115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05206_ cpu.decode.co_mem_word _01342_ _01406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_111_Right_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06186_ rf_ram.memory\[465\]\[1\] _01697_ _02381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_29_1171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05137_ cpu.decode.op21 _01335_ _01339_ _01340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XANTENNA__05467__B _01504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_70_1701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09945_ rf_ram.memory\[338\]\[0\] _04932_ _04933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09876_ _03309_ _02954_ _04890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08827_ _04202_ _04213_ _04214_ _00806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09730__A2 net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07741__A1 _03524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06544__A2 _01366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08758_ _04170_ _04168_ _04171_ _00780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_174_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_1131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_1180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07709_ _03491_ _03503_ _03505_ _00397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_68_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08689_ rf_ram.memory\[154\]\[0\] _04127_ _04128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10720_ _00464_ clknet_leaf_50_clk rf_ram.memory\[462\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_177_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_83_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_101_2266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_101_2277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10651_ _00395_ clknet_leaf_115_clk rf_ram.memory\[400\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09246__A1 _02714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_81_1896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_180_425 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10582_ _00326_ clknet_leaf_163_clk rf_ram.memory\[322\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09797__A2 _02921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09261__A4 _01460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_134_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_146_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_160_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06480__B2 rf_ram.memory\[13\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_1027 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11203_ _00939_ clknet_leaf_50_clk rf_ram.memory\[85\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05377__B _01528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08221__A2 _03072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_1146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_147_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11134_ _00870_ clknet_leaf_74_clk rf_ram.memory\[113\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_102_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_164_3440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11065_ _00802_ clknet_leaf_11_clk rf_ram.memory\[137\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_108_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10016_ _02910_ _02984_ _04976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09721__A2 net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_125_2712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_125_2723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_160_3359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07732__A1 _03488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06001__B _01528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_1220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_99_884 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_1231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09485__A1 _01411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08288__A2 _02904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_157_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06299__A1 _01552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10095__A2 _02909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_184_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10918_ _00662_ clknet_leaf_16_clk rf_ram.memory\[177\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_74_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_157_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_989 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10849_ _00593_ clknet_leaf_310_clk rf_ram.memory\[532\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_128_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_171_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_109_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_14_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_48_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_280_clk_I clknet_5_19__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06040_ _02211_ _02234_ _02235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_125_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1079 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_184_3805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_184_3816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06223__A1 _01675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_295_clk_I clknet_5_7__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07991_ _03651_ _03679_ _03680_ _00504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_10_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07971__A1 _03654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09730_ _04781_ net12 _04798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_157_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06942_ rf_ram.memory\[206\]\[0\] _03023_ _03024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09661_ _03974_ _04736_ _04745_ _04746_ _01108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_158_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06873_ _02813_ _02941_ _02977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_59_1142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_2_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08612_ _04058_ _04079_ _04080_ _00725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_179_525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05824_ rf_ram.memory\[214\]\[0\] _01940_ _02019_ rf_ram.memory\[215\]\[0\] _01968_
+ rf_ram.memory\[213\]\[0\] _02020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_09592_ _01469_ _04698_ _01491_ _04703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05306__I _01501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_94_1099 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08543_ _04023_ _04034_ _04035_ _00701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05755_ _01693_ _01951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_49_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_233_clk_I clknet_5_23__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_147_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05686_ _01769_ _01880_ _01881_ _01882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_08474_ _01378_ rf_ram_if.rtrig1 rf_ram.rdata\[1\] _03988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_148_956 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_175_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_174_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_163_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07425_ rf_ram.memory\[333\]\[0\] _03328_ _03329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_58_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_148_989 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_147_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09228__A1 _04434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_175_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_63_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_163_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_134_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07356_ rf_ram.memory\[252\]\[1\] _03283_ _03285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_18_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_1102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_248_clk_I clknet_5_21__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_150_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06307_ _02499_ _02501_ _01564_ _02502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_165_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07287_ _03222_ _03241_ _03242_ _00238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_45_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06238_ rf_ram.memory\[436\]\[1\] _01510_ _02433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05265__A2 cpu.decode.co_ebreak vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09026_ _04331_ _04336_ _04337_ _00882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_170_491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06169_ rf_ram.memory\[510\]\[1\] _01631_ _02364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08203__A2 _03811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07962__A1 _02836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09928_ _04921_ _04919_ _04922_ _01200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_102_1066 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09703__A2 net4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_142_3034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09859_ _04878_ _04879_ _04870_ _04880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_99_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07714__A1 _03491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09911__I _02814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_103_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_103_2317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_120_2620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_83_1936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_120_2631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_83_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_166_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10703_ _00447_ clknet_leaf_90_clk rf_ram.memory\[411\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_165_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09219__A1 _03319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_181_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10634_ _00378_ clknet_leaf_102_clk rf_ram.memory\[404\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_183_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10565_ _00309_ clknet_leaf_171_clk rf_ram.memory\[366\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_107_875 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_1235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_118_2582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_162_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_45_1208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06453__A1 _01526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_118_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_161_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10496_ _00240_ clknet_leaf_53_clk rf_ram.memory\[468\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_51_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_121_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10001__A2 _02992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_1100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_1310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11117_ _00853_ clknet_leaf_113_clk rf_ram.memory\[449\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_36_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11048_ _00785_ clknet_leaf_337_clk rf_ram.memory\[144\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07705__A1 _02960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput8 i_dbus_rdt[15] net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05192__A1 _01391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_99_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_1181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10068__A2 _03158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05540_ rf_ram.memory\[276\]\[0\] _01735_ _01736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05570__B _01349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_1023 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_177_3675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_157_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08130__A1 _03757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_1034 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_177_3686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_5_20__f_clk_I clknet_3_5_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_1102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_139_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05471_ rf_ram.memory\[368\]\[0\] _01666_ _01526_ _01667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__06141__B1 _01715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_89_1135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09469__S _04604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07210_ _03193_ _03191_ _03194_ _00209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_138_2958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06692__A1 _02788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08190_ rf_ram.memory\[53\]\[0\] _03805_ _03806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_61_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_171_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07141_ _02795_ _02911_ _03151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_27_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_41_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09630__A1 _04643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07072_ _02844_ _02911_ _03108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_124_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_124_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06023_ rf_ram.memory\[548\]\[1\] _01538_ _01539_ rf_ram.memory\[549\]\[1\] _01540_
+ rf_ram.memory\[551\]\[1\] _02218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XANTENNA__09394__B1 _04564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08736__A3 _03984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07944__A1 _03622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05745__B _01805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07974_ rf_ram.memory\[46\]\[0\] _03669_ _03670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_96_1139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09713_ _04781_ net7 _04786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_87_2014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06925_ rf_ram.memory\[278\]\[1\] _03010_ _03012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09697__A1 _04740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_173_1318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09644_ cpu.mem_bytecnt\[1\] _01376_ _04731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06856_ _02927_ _02964_ _02965_ _00084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_136_1140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_172_clk_I clknet_5_30__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05807_ _01991_ _01995_ _01999_ _02002_ _02003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_09575_ cpu.immdec.imm30_25\[4\] _04688_ _04678_ _04689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_65_1600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06787_ _02916_ _02917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_65_1611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_132_1026 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08526_ rf_ram.memory\[49\]\[0\] _04024_ _04025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_72_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05738_ _01914_ _01921_ _01929_ _01933_ _01934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_38_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08347__I _03902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_52_clk_I clknet_5_9__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_148_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06295__C _01349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_175_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08457_ net109 _03974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_148_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05669_ _01769_ _01862_ _01864_ _01865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__08672__A2 _04078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_187_clk_I clknet_5_28__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07408_ _03289_ _03316_ _03317_ _00284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_19_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06683__A1 _02750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08388_ rf_ram.memory\[189\]\[1\] _03927_ _03929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_61_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05891__C1 _01912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_67_clk_I clknet_5_8__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07339_ rf_ram.memory\[270\]\[0\] _03274_ _03275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09621__A1 _02828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05238__A2 _01436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06435__A1 _01569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_110_clk_I clknet_5_15__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10350_ _00094_ clknet_leaf_180_clk rf_ram.memory\[281\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_61_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_21_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09009_ _04298_ _04325_ _04326_ _00876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10281_ _00025_ clknet_leaf_143_clk rf_ram.memory\[294\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_14_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08188__A1 _03790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_113_2490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07935__A1 _02752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_125_clk_I clknet_5_13__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05655__B _01693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05946__B1 _01607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05374__C _01569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09688__A1 _04740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08360__A1 _03884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_158_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_14_Left_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06371__B1 _01625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06486__B _01525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_159_3350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_154_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11383__CLK clknet_5_23__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_425 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_155_3269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_154_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11666_ net117 net189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_83_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_126_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10617_ _00361_ clknet_leaf_156_clk rf_ram.memory\[353\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_172_3583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_172_3594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09612__A1 _04637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09463__I1 net82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11597_ _00000_ clknet_leaf_282_clk rf_ram.rdata\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_106_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10548_ _00292_ clknet_leaf_149_clk rf_ram.memory\[370\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_150_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_23_Left_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_133_2866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_1196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05634__C1 _01678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10479_ _00223_ clknet_leaf_104_clk rf_ram.memory\[421\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08179__A1 _03798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09679__A1 net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06710_ rf_ram.memory\[521\]\[1\] _02859_ _02861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07690_ rf_ram.memory\[401\]\[0\] _03493_ _03494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_179_3715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_154_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_32_Left_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_179_3726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06641_ _02748_ _02807_ _02809_ _00025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05165__A1 _01353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06362__B1 _01953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09360_ _04551_ _01002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06572_ rf_ram.memory\[201\]\[1\] _02753_ _02755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08103__A1 _02780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_176_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08311_ rf_ram.memory\[243\]\[1\] _03878_ _03880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_75_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05523_ _01686_ _01719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_09291_ rf_ram.memory\[65\]\[1\] _04508_ _04510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09851__A1 _02713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08242_ rf_ram.memory\[52\]\[0\] _03837_ _03838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05454_ _01601_ _01650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_117_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08173_ _02881_ _02917_ _03795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05385_ _01495_ _01575_ _01580_ _01581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_160_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09603__A1 _04643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09454__I1 net78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_41_Left_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_162_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_1252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07124_ rf_ram.memory\[487\]\[1\] _03139_ _03141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_31_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07055_ _02806_ _02869_ _03097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_140_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput120 net120 o_dbus_dat[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_140_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput131 net131 o_dbus_sel[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput142 net142 o_ext_rs1[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_06006_ rf_ram.memory\[532\]\[1\] _01523_ _01516_ rf_ram.memory\[533\]\[1\] _01520_
+ rf_ram.memory\[535\]\[1\] _02201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XTAP_TAPCELL_ROW_58_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_100_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_58_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05640__A2 _01755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09906__A2 _02883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput153 net153 o_ext_rs1[23] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput164 net164 o_ext_rs1[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput175 net175 o_ext_rs2[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__07917__A1 _03619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput186 net186 o_ext_rs2[24] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput197 net197 o_ext_rs2[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__05928__B1 _01848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input35_I i_ibus_rdt[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_1183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07957_ _02903_ _03158_ _03659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_177_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_138_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06908_ _02975_ _02998_ _03000_ _00101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07888_ _02959_ _03234_ _03616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09627_ _04643_ _01400_ _04660_ _01098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_69_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06839_ _02779_ _02786_ _02953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_168_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_167_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09558_ _01469_ _01433_ _02711_ _04676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_183_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05171__A4 _01373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08509_ _01381_ _01469_ _04012_ _01399_ _04013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_136_701 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_182_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09842__A1 _02714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09489_ _02690_ _04622_ _04624_ _04616_ _01058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_38_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_148_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11520_ _01252_ clknet_leaf_199_clk rf_ram.memory\[507\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_136_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09410__B _04539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_163_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1027 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11451_ _01183_ clknet_leaf_281_clk rf_ram.memory\[229\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_163_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06408__A1 _01768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10402_ _00146_ clknet_leaf_301_clk rf_ram.memory\[215\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10204__A2 _02866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_115_2530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05369__C _01564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11382_ _01114_ clknet_leaf_229_clk net127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_78_1846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_1205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_115_2541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_132_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_78_1857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_150_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05616__C1 _01811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_150_3188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07081__A1 _03092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10333_ _00077_ clknet_leaf_146_clk rf_ram.memory\[304\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_132_984 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05631__A2 _01777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10264_ _00008_ clknet_leaf_33_clk rf_ram.memory\[200\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10195_ rf_ram.memory\[210\]\[0\] _05086_ _05087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05919__B1 _01931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07156__I _03017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09572__S _04678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_156_1313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_89_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08333__A1 _03884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07136__A2 _02923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06344__B1 _01636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_194_clk clknet_5_28__leaf_clk clknet_leaf_194_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08884__A2 _04248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_157_3309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06895__A1 _02716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_97_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05404__I _01599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_174_3623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_174_3634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_1173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_173_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08636__A2 _04067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_135_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11649_ net99 net171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput11 i_dbus_rdt[18] net11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_114_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09436__I1 net69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput22 i_dbus_rdt[28] net22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_154_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_140_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput33 i_dbus_rdt[9] net33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_114_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput44 i_ibus_rdt[19] net44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05170_ _01353_ cpu.immdec.imm19_12_20\[8\] _01367_ cpu.immdec.imm24_20\[4\] _01373_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
Xinput55 i_ibus_rdt[2] net55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_3_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput66 i_timer_irq net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_13_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07072__A1 _02844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06280__C1 _01968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05622__A2 _01543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_876 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_1144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08860_ _04057_ _04234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_36_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_36_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08572__A1 _04026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07375__A2 _02813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07811_ net236 _03234_ _03569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08791_ _04170_ _04189_ _04191_ _00793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_97_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_1109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07742_ _02788_ _03481_ _03526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08324__A1 _03887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05138__A1 cpu.state.genblk1.misalign_trap_sync_r vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07673_ rf_ram.memory\[384\]\[0\] _03482_ _03483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10131__A1 _02805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_185_clk clknet_5_28__leaf_clk clknet_leaf_185_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_88_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09412_ net246 _02801_ _04581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05689__A2 _01777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06624_ cpu.immdec.imm11_7\[2\] _02730_ _02796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_94_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05314__I _01509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09343_ _04542_ _00994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_87_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06555_ _01353_ rf_ram_if.wdata1_r\[0\] _02740_ _02741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_176_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_158_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09824__A1 _04837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_158_Right_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_164_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05506_ _01609_ _01702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_12
XFILLER_0_114_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_118_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09274_ cpu.genblk3.csr.mcause3_0\[0\] _04496_ _04497_ _04498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_145_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06486_ rf_ram.memory\[0\]\[1\] _01613_ _01525_ _02681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_106_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08225_ _03823_ _03825_ _03827_ _00591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05437_ _01508_ _01633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_145_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08156_ net238 _03765_ _03784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_43_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05368_ _01563_ _01564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_95_2157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10198__A1 _05081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_95_2168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07107_ rf_ram.memory\[501\]\[1\] _03128_ _03130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_30_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05299_ _01494_ _01495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_08087_ _03724_ _03739_ _03741_ _00539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_141_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09456__I _01411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05613__A2 _01808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06810__A1 _02927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07038_ _03050_ _03084_ _03085_ _00146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_11_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_73_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_73_1765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_41_1255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08563__A1 _02915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06023__C1 _01540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08989_ _04298_ _04313_ _04314_ _00868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05933__B net251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08315__A1 _03852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_1140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_27_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10951_ _00689_ clknet_leaf_18_clk rf_ram.memory\[79\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_176_clk clknet_5_30__leaf_clk clknet_leaf_176_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_138_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10122__A1 _05014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_27_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06326__B1 _02019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06877__A1 _02975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10130__I _02742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10882_ _00626_ clknet_leaf_32_clk rf_ram.memory\[220\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_79_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_38_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_183_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_183_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_149_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_125_Right_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_65_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_93_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_38_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_152_3217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06483__C _01562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11503_ _01235_ clknet_leaf_199_clk rf_ram.memory\[505\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_164_884 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_53_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11434_ _01166_ clknet_leaf_242_clk cpu.state.cnt_r\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05852__A2 _01614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07054__A1 _03092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_130_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_130_2814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_100_clk clknet_5_14__leaf_clk clknet_leaf_100_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_132_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11365_ _01097_ clknet_leaf_235_clk cpu.bne_or_bge vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__05604__A2 _01799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10316_ _00060_ clknet_leaf_271_clk rf_ram.memory\[512\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11296_ _01029_ clknet_leaf_253_clk net91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_10247_ rf_ram.memory\[264\]\[1\] _05116_ _05118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_167_3493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10178_ rf_ram.memory\[202\]\[0\] _05075_ _05076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_128_2765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05843__B _01860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_128_2776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07109__A2 _02911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_167_clk clknet_5_30__leaf_clk clknet_leaf_167_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_44_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_187_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_146_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09806__A1 _04840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06340_ rf_ram.memory\[206\]\[1\] _01531_ _02535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_173_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_121_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06271_ rf_ram.memory\[152\]\[1\] _01735_ _01956_ _02466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_44_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05222_ _01385_ cpu.state.o_cnt\[2\] cpu.mem_bytecnt\[1\] _01422_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08010_ _02959_ _03693_ _03694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_25_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_170_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_167_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_114_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_7_Left_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_52_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05153_ cpu.decode.op21 _01343_ _01336_ _01356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_170_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_38_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_38_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_187_3858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_187_3869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09961_ _04918_ _04941_ _04942_ _01213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_110_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_90_2065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08912_ _04057_ _04266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_90_2076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09892_ rf_ram.memory\[18\]\[0\] _04899_ _04900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08545__A1 _04026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05309__I _01504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07348__A2 _02997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08843_ rf_ram.memory\[134\]\[1\] _04222_ _04224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_51_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06020__A2 _01532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08774_ _04167_ _04180_ _04181_ _00786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05986_ _02178_ _02179_ _02180_ _02181_ _01493_ _02182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__07524__I _03100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_79_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07725_ _02795_ _02869_ _03515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10104__A1 _05017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_158_clk clknet_5_27__leaf_clk clknet_leaf_158_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__06859__A1 _02822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07656_ _03088_ _03135_ _03472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_178_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_138_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_0_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_0_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06607_ rf_ram.memory\[235\]\[0\] _02782_ _02783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07587_ _03425_ _03427_ _03429_ _00351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_47_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09326_ rf_ram.memory\[109\]\[1\] _04530_ _04532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06538_ rf_ram.i_raddr\[3\] _02717_ _02724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XTAP_TAPCELL_ROW_97_2208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_152_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_11_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06087__A2 _01652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07284__A1 _03225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09257_ _04484_ _01484_ _04485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xclkbuf_leaf_330_clk clknet_5_1__leaf_clk clknet_leaf_330_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_06469_ rf_ram.memory\[18\]\[1\] _01605_ _01624_ rf_ram.memory\[19\]\[1\] _02663_
+ _02664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_145_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08208_ _03790_ _03814_ _03816_ _00585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_16_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05834__A2 _01501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09188_ _04434_ _04436_ _04438_ _00943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_160_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output189_I net189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07036__A1 _02738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08139_ rf_ram.memory\[54\]\[1\] _03772_ _03774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08784__A1 _04167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11150_ _00886_ clknet_leaf_67_clk rf_ram.memory\[105\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_144_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05647__C _01670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10101_ rf_ram.memory\[311\]\[0\] _05028_ _05029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_max_cap235_I _03082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11081_ _00818_ clknet_leaf_27_clk rf_ram.memory\[131\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_41_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08536__A1 _02865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10032_ _04985_ _04983_ _04986_ _01240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06011__A2 _01538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_145_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_187_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_149_clk clknet_5_26__leaf_clk clknet_leaf_149_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_59_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_106_2359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_169_954 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10934_ net258 clknet_leaf_261_clk rf_ram_if.wdata1_r\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_169_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_123_2673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_86_1989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_123_2684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_1233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_39_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10865_ _00609_ clknet_leaf_42_clk rf_ram.memory\[197\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_155_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_1181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_1200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10796_ _00540_ clknet_leaf_320_clk rf_ram.memory\[558\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_38_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_1079 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07275__A1 _02899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06078__A2 _01687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_321_clk clknet_5_5__leaf_clk clknet_leaf_321_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_81_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_843 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11417_ _01149_ clknet_leaf_287_clk rf_ram.memory\[58\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_50_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_169_3533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11348_ _01080_ clknet_leaf_254_clk cpu.immdec.imm30_25\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_22_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06250__A2 _01799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11279_ _01014_ clknet_leaf_244_clk net215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_33_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08527__A1 _04023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_33_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_182_3766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_158_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_182_3777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06002__A2 _01544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05840_ _01972_ _02034_ _02035_ _02036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_55_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_169_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05771_ rf_ram.memory\[148\]\[0\] _01523_ _01967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07510_ _03356_ _03380_ _03381_ _00322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_18_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08490_ _03953_ _03998_ _03999_ _00684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_18_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_162_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_159_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_1076 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07441_ _03323_ _03337_ _03338_ _00296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_147_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_1270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07372_ _03289_ _03294_ _03295_ _00270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_130_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09255__A2 _01356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_1292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_1254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09111_ _04367_ _04387_ _04389_ _00915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06069__A2 _01543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06323_ _01768_ _02506_ _02517_ _01569_ _02518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
Xclkbuf_leaf_312_clk clknet_5_5__leaf_clk clknet_leaf_312_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_73_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05816__A2 _01922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09042_ _04331_ _04346_ _04347_ _00888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06254_ rf_ram.memory\[428\]\[1\] _01724_ _01725_ rf_ram.memory\[429\]\[1\] _01726_
+ rf_ram.memory\[431\]\[1\] _02449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_170_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_60_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09007__A2 _04303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_92_2105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05205_ cpu.decode.co_mem_word cpu.bne_or_bge _01405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_92_2116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06185_ rf_ram.memory\[464\]\[1\] _01782_ _01693_ _02380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_142_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08766__A1 _04170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06226__C1 _01608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_1183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_1063 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05136_ cpu.decode.opcode\[2\] cpu.branch_op _01339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_111_740 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_180_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09944_ _04911_ _02923_ _04932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06241__A2 _01782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_70_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08518__A1 _03956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09875_ _02713_ _04889_ _01180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09191__A1 _04431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08826_ rf_ram.memory\[135\]\[0\] _04213_ _04214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_174_1051 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_169_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08757_ rf_ram.memory\[146\]\[1\] _04168_ _04171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05752__A1 net252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05969_ rf_ram.memory\[24\]\[0\] _01682_ _01550_ _02165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_68_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07708_ rf_ram.memory\[381\]\[1\] _03503_ _03505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_68_1664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08688_ _02812_ _04078_ _04127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_75_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_71_1034 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_166_913 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07639_ rf_ram.memory\[406\]\[1\] _03460_ _03462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_output104_I net104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_101_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10650_ _00394_ clknet_leaf_115_clk rf_ram.memory\[400\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_101_2278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_635 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07257__A1 _02894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09309_ _04477_ _01491_ _04013_ _04521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_0_119_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_81_1897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10581_ _00325_ clknet_leaf_162_clk rf_ram.memory\[362\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_303_clk clknet_5_6__leaf_clk clknet_leaf_303_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_63_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06465__C1 _01617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_1174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_133_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07009__A1 _03050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_16_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06480__A2 _01643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05658__B _01790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11202_ _00938_ clknet_leaf_49_clk rf_ram.memory\[85\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_47_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06232__A2 _01509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_147_3127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11133_ _00869_ clknet_leaf_74_clk rf_ram.memory\[114\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_43_1158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_164_3441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_79_Left_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_11064_ _00801_ clknet_leaf_11_clk rf_ram.memory\[138\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05991__A1 _02017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10015_ _04953_ _04973_ _04975_ _01234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05393__B _01528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_125_2713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_125_2724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09485__A2 _03989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_169_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10917_ _00661_ clknet_leaf_16_clk rf_ram.memory\[178\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_184_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_1074 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_88_Left_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_128_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_132_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10848_ _00592_ clknet_leaf_311_clk rf_ram.memory\[532\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_26_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05412__I _01607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07248__A1 _03190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_171_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_172_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_171_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10779_ _00523_ clknet_leaf_328_clk rf_ram.memory\[567\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_27_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_87_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08996__A1 _04301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_152_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06471__A2 _01682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_140_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_164_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_50_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_184_3806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_184_3817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_97_Left_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07420__A1 _03323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07990_ rf_ram.memory\[477\]\[0\] _03679_ _03680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06941_ _02738_ _02972_ _03023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06399__B _01684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09660_ net1 net13 _04736_ _04746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06872_ _02975_ _02973_ _02976_ _00089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_94_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08611_ rf_ram.memory\[129\]\[0\] _04079_ _04080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_94_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_2_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05823_ _01695_ _02019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_09591_ _04702_ _01082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_94_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_55_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_179_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_173_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08542_ rf_ram.memory\[171\]\[0\] _04034_ _04035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05754_ _01373_ _01817_ _01949_ _01950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_166_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07487__A1 _03360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08473_ _03987_ _00679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05685_ rf_ram.memory\[396\]\[0\] _01711_ _01772_ rf_ram.memory\[397\]\[0\] _01773_
+ rf_ram.memory\[399\]\[0\] _01881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_147_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07424_ _03319_ _02844_ _03328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_92_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_1040 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_63_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_175_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_135_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07355_ _03257_ _03283_ _03284_ _00264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_169_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08987__A1 net236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06306_ rf_ram.memory\[170\]\[1\] _01989_ _01520_ rf_ram.memory\[171\]\[1\] _02500_
+ _02501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_33_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07286_ rf_ram.memory\[471\]\[0\] _03241_ _03242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_5_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_171_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09025_ rf_ram.memory\[107\]\[0\] _04336_ _04337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_170_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06237_ _01768_ _02419_ _02431_ net254 _02432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_32_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input65_I i_rst vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06168_ _02351_ _02355_ _02359_ _02362_ _02363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_13_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06214__A2 _01697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_1170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06099_ _01675_ _02292_ _02293_ _02294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__07962__A2 _03009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09927_ rf_ram.memory\[342\]\[1\] _04919_ _04922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_102_1078 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09164__A1 _04397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09858_ _01399_ _01381_ _02710_ _04879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_176_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_142_3024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_142_3035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_1243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08911__A1 _04237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08809_ net247 _04195_ _04203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_38_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09789_ _04637_ _04834_ _04836_ _01146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_96_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_103_2307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05941__B _01550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_103_2318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08808__I _04057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_157_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_83_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_120_2621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07478__A1 _02728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_166_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_83_1948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_120_2632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_80_clk clknet_5_11__leaf_clk clknet_leaf_80_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_113_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10702_ _00446_ clknet_leaf_89_clk rf_ram.memory\[411\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_55_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06150__A1 _01600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_1225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09219__A2 _02960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10633_ _00377_ clknet_leaf_80_clk rf_ram.memory\[386\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_119_670 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10564_ _00308_ clknet_leaf_171_clk rf_ram.memory\[366\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_10_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_162_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_1247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_118_2583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07650__A1 _03458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05388__B _01552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_20_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_118_2594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_1269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10495_ _00239_ clknet_leaf_54_clk rf_ram.memory\[471\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_20_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09575__S _04678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06205__A2 _01801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_9_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11116_ _00852_ clknet_leaf_113_clk rf_ram.memory\[449\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_120_1134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_1322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05964__A1 _01903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09155__A1 _04401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11047_ _00784_ clknet_leaf_337_clk rf_ram.memory\[144\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06012__B _01552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07705__A2 _03496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05407__I _01602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08902__A1 _02916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput9 i_dbus_rdt[16] net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_308_clk_I clknet_5_5__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05192__A2 net134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_71_clk clknet_5_8__leaf_clk clknet_leaf_71_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_188_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_177_3676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_911 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_177_3687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_157_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05470_ _01643_ _01666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_129_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_28_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06692__A2 _02846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_171_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_138_2959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07140_ _03126_ _03148_ _03150_ _00183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_109_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09630__A2 _01382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07641__A1 _02889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07071_ _03092_ _03105_ _03107_ _00157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06444__A2 _01513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06022_ rf_ram.memory\[550\]\[1\] _01502_ _01506_ _02217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_113_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_1164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_61_1066 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07973_ _03668_ _02972_ _03669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09146__A1 net250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09712_ _04785_ _01120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_87_2015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06924_ _02970_ _03010_ _03011_ _00106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09697__A2 net33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09643_ _04637_ _04728_ _04730_ _01106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06855_ rf_ram.memory\[284\]\[0\] _02964_ _02965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_78_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05761__B _01956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05806_ _01552_ _02000_ _02001_ _02002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_136_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09574_ cpu.immdec.imm30_25\[5\] net54 _03967_ _04688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06786_ _02773_ _02837_ _02916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__06380__A1 _01368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_65_1601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_65_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08525_ net248 _02869_ _04024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05737_ _01909_ _01930_ _01932_ _01933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_33_1102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_888 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_62_clk clknet_5_8__leaf_clk clknet_leaf_62_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_92_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_136_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08456_ net98 _03973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05668_ rf_ram.memory\[476\]\[0\] _01863_ _01848_ rf_ram.memory\[477\]\[0\] _01778_
+ rf_ram.memory\[479\]\[0\] _01864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_0_175_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_93_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07407_ rf_ram.memory\[372\]\[0\] _03316_ _03317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_92_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07880__A1 _03587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08387_ _03919_ _03927_ _03928_ _00652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05599_ _01675_ _01792_ _01794_ _01795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_107_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05891__B1 _01925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07338_ _02958_ _02972_ _03274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_34_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09621__A2 _04507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07632__A1 _03455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05238__A3 _01437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06435__A2 _02618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07269_ _03230_ _02899_ _03231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_103_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_1112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_143_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09008_ rf_ram.memory\[110\]\[0\] _04325_ _04326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10280_ _00024_ clknet_leaf_145_clk rf_ram.memory\[294\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_991 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output171_I net171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_113_2491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07935__A2 _02832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09688__A2 net30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07699__A1 _03491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05671__B _01707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05390__C _01495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_159_3340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_159_3351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_53_clk clknet_5_12__leaf_clk clknet_leaf_53_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_95_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_1246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_294_clk_I clknet_5_7__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_25_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_25_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_126_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11665_ net116 net188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_36_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10616_ _00360_ clknet_leaf_156_clk rf_ram.memory\[353\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_181_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_172_3584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_135_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11596_ _01328_ clknet_leaf_38_clk rf_ram.memory\[9\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_172_3595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_91_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06426__A2 _01989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07623__A1 _03425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10547_ _00291_ clknet_leaf_167_clk rf_ram.memory\[333\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06007__B _01552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05634__B1 _01688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_133_2867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10478_ _00222_ clknet_leaf_104_clk rf_ram.memory\[421\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_121_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_161_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08179__A2 _02960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05846__B _01650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_232_clk_I clknet_5_23__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_10_Right_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_21_1072 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_247_clk_I clknet_5_21__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_139_Right_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_179_3716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_1184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06640_ rf_ram.memory\[294\]\[1\] _02807_ _02809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_56_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_151_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_63_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06571_ _02743_ _02753_ _02754_ _00010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_leaf_44_clk clknet_5_12__leaf_clk clknet_leaf_44_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08103__A2 _03729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08310_ _03852_ _03878_ _03879_ _00624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09300__A1 _04463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05522_ _01708_ _01710_ _01712_ _01716_ _01717_ _01718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XTAP_TAPCELL_ROW_43_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09290_ _04463_ _04508_ _04509_ _00974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06114__A1 _01527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_185_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_170_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08241_ _03668_ _03135_ _03837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_6_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_60_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05453_ _01613_ _01649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__07862__A1 _03590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_184_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_172_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_133_919 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08172_ _03790_ _03792_ _03794_ _00571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_28_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05384_ _01576_ _01577_ _01578_ _01579_ _01495_ _01580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_55_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_172_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07123_ _03123_ _03139_ _03140_ _00176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_126_993 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07614__A1 _03445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06417__A2 _01918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_1106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_113_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07054_ _03092_ _03094_ _03096_ _00151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xoutput110 net110 o_dbus_dat[20] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_113_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput121 net121 o_dbus_dat[30] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput132 net132 o_dbus_sel[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_06005_ rf_ram.memory\[534\]\[1\] _01532_ _01505_ _02200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_140_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput143 net143 o_ext_rs1[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_58_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput154 net154 o_ext_rs1[24] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_58_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput165 net165 o_ext_rs1[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_56_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xoutput176 net176 o_ext_rs2[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput187 net187 o_ext_rs2[25] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__05475__C _01670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05389__C1 _01555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput198 net198 o_ext_rs2[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__09119__A1 _04364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06050__B1 _01608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07956_ _03654_ _03656_ _03658_ _00491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input28_I i_dbus_rdt[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06907_ rf_ram.memory\[2\]\[1\] _02998_ _03000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07887_ _03590_ _03613_ _03615_ _00465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_98_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_106_Right_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06838_ _02930_ _02950_ _02952_ _00079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09626_ _04643_ _01452_ _04658_ _01097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_69_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_179_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09557_ cpu.immdec.imm30_25\[1\] net50 _03967_ _04675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06769_ _02716_ _02887_ _02903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_38_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_35_clk clknet_5_6__leaf_clk clknet_leaf_35_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08508_ _01469_ net134 _04012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_38_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09488_ net87 _03989_ _04622_ _04624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_109_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_176_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_1111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08439_ _02953_ _03949_ _03961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_114_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07853__A1 _02971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_1310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_92_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11450_ _01182_ clknet_leaf_284_clk rf_ram.memory\[239\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_68_1039 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05510__I _01686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_530 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_117_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_163_598 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10401_ _00145_ clknet_leaf_300_clk rf_ram.memory\[216\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07605__A1 _03422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11381_ _01113_ clknet_leaf_229_clk net126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_116_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_1847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_115_2531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_115_2542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05616__B1 _01810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_150_3178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_78_1858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_1217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_150_3189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10332_ _00076_ clknet_leaf_146_clk rf_ram.memory\[304\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10263_ _02825_ _05125_ _05127_ _01330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08030__A1 _03668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10194_ _03892_ _02923_ _05086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_121_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_79_1146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06592__A1 _02743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09652__I net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_950 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_26_clk clknet_5_3__leaf_clk clknet_leaf_26_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08097__A1 _03724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_174_3624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_1077 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_68_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07844__A1 _03587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_166_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_154_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_135_2907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11648_ net129 net201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput12 i_dbus_rdt[19] net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput23 i_dbus_rdt[29] net23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09597__A1 _03992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput34 i_ibus_ack net34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_163_1318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput45 i_ibus_rdt[20] net45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_11579_ _01311_ clknet_leaf_34_clk rf_ram.memory\[207\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput56 i_ibus_rdt[30] net56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_107_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07072__A2 _02911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_171_clk_I clknet_5_30__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06280__B1 _01959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_51_clk_I clknet_5_12__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_36_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07810_ _03557_ _03566_ _03568_ _00435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_36_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08790_ rf_ram.memory\[149\]\[1\] _04189_ _04191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05386__A2 _01532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06583__A1 _02731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_186_clk_I clknet_5_28__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07741_ _03524_ _03522_ _03525_ _00409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_leaf_66_clk_I clknet_5_8__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09521__A1 _03967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07672_ _02904_ _03481_ _03482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08178__I _02845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05138__A2 cpu.genblk3.csr.o_new_irq vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10131__A2 _02832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09411_ _04576_ _04580_ _01024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_176_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06623_ _02794_ _02795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_48_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_983 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_17_clk clknet_5_2__leaf_clk clknet_leaf_17_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_181_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09342_ net213 _03991_ _04540_ net224 _04542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06554_ _01369_ rf_ram_if.wdata0_r\[0\] _02740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__08088__A1 _02971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_1188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05505_ rf_ram.memory\[340\]\[0\] _01537_ _01701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07835__A1 _03557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09273_ _01387_ _01465_ _04481_ _04497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_75_666 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_173_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06485_ rf_ram.memory\[4\]\[1\] _01643_ _01714_ rf_ram.memory\[5\]\[1\] _01635_ rf_ram.memory\[7\]\[1\]
+ _02680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_117_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_47_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_124_clk_I clknet_5_13__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08224_ rf_ram.memory\[533\]\[1\] _03825_ _03827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05436_ rf_ram.memory\[366\]\[0\] _01631_ _01632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_16_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05330__I _01525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09588__A1 _02709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08155_ _03757_ _03781_ _03783_ _00565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_28_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05367_ _01562_ _01563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_31_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_95_2158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_95_2169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07106_ _03123_ _03128_ _03129_ _00170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_leaf_139_clk_I clknet_5_27__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08260__A1 _03823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08086_ rf_ram.memory\[55\]\[1\] _03739_ _03741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05298_ _01493_ _01494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_07037_ rf_ram.memory\[215\]\[0\] _03084_ _03085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_28_1089 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_19_clk_I clknet_5_2__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08012__A1 _03686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_73_1755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_110_2450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06023__B1 _01539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08563__A2 _02960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08988_ rf_ram.memory\[114\]\[0\] _04313_ _04314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05377__A2 _01524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_1000 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output134_I net134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07939_ _03622_ _03645_ _03647_ _00485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_39_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10950_ _00688_ clknet_leaf_18_clk rf_ram.memory\[79\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_27_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_168_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_1016 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09609_ rf_ram.memory\[73\]\[0\] _04714_ _04715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_39_1196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10881_ _00625_ clknet_leaf_282_clk rf_ram.memory\[243\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_74_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_109_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07826__A1 _02839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_152_3218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11502_ _01234_ clknet_leaf_191_clk rf_ram.memory\[348\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_1183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_81_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09579__A1 _01391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11433_ _01165_ clknet_leaf_238_clk cpu.state.cnt_r\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_145_1015 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10189__A2 _02972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_130_2804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08251__A1 _02845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_85_1183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11364_ _01096_ clknet_leaf_63_clk rf_ram.memory\[71\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_130_2815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10315_ _00059_ clknet_leaf_267_clk rf_ram.memory\[513\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05396__B _01351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11295_ _01028_ clknet_leaf_250_clk net90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_120_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_60_Left_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10246_ _02819_ _05116_ _05117_ _01323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08003__A1 _03686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_167_3494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10177_ _03892_ _02775_ _05075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_128_2766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05773__C1 _01968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_128_2777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_1230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09503__A1 _04634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_158_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_1072 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05540__A2 _01735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05828__B1 _02019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_13_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06270_ _01951_ _02463_ _02464_ _02465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__08490__A1 _03953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_170_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_167_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_154_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05221_ _01416_ _01420_ _01421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_71_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_738 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_53_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_170_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05152_ cpu.immdec.imm24_20\[1\] _01338_ _01344_ _01355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_123_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_38_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_38_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_187_3859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09990__A1 _04953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09960_ rf_ram.memory\[335\]\[0\] _04941_ _04942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_6_clk clknet_5_2__leaf_clk clknet_leaf_6_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_40_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_55_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_90_2066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_111_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08911_ _04237_ _04263_ _04265_ _00839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_90_2077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09891_ _02922_ _03035_ _04899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08842_ _04202_ _04222_ _04223_ _00812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_51_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_1005 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_97_1054 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08773_ rf_ram.memory\[143\]\[0\] _04180_ _04181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_100_1165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05985_ rf_ram.memory\[2\]\[0\] _01661_ _01635_ rf_ram.memory\[3\]\[0\] _01714_ rf_ram.memory\[1\]\[0\]
+ _02181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_97_1098 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07724_ _03491_ _03512_ _03514_ _00403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_79_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05325__I _01520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_108_Left_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_19_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07655_ _03458_ _03469_ _03471_ _00377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06859__A2 _02941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06606_ _02766_ _02781_ _02782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_0_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07586_ rf_ram.memory\[316\]\[1\] _03427_ _03429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05531__A2 _01724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09325_ _04463_ _04530_ _04531_ _00987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07808__A1 _03554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06537_ _02720_ _02722_ _02723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_0_91_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_97_2209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_11_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_146_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09256_ _01356_ _04484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_90_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06468_ rf_ram.memory\[17\]\[1\] _01514_ _02663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_91_956 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08207_ rf_ram.memory\[536\]\[1\] _03814_ _03816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_32_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_146_1313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05419_ _01550_ _01615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_106_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09187_ rf_ram.memory\[179\]\[1\] _04436_ _04438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_161_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06399_ rf_ram.memory\[88\]\[1\] _01683_ _01684_ _02594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_90_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08138_ _03754_ _03772_ _03773_ _00558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08233__A1 _03820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07036__A2 _03083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10040__A1 _04982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09981__A1 _02865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08069_ rf_ram.memory\[562\]\[0\] _03730_ _03731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_102_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05598__A2 _01777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10100_ _02800_ _03083_ _05028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11080_ _00817_ clknet_leaf_15_clk rf_ram.memory\[132\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_179_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_80_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10031_ rf_ram.memory\[327\]\[1\] _04983_ _04986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08536__A2 _03945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09733__A1 _04781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05944__B _01493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_5_26__f_clk clknet_3_6_0_clk clknet_5_26__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_145_3088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_169_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05507__C1 _01702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10933_ rf_ram_if.wdata1_r\[1\] clknet_leaf_261_clk rf_ram_if.wdata1_r\[0\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_58_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_85_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_123_2674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_169_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_1223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_123_2685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_151_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10864_ _00608_ clknet_leaf_42_clk rf_ram.memory\[197\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_184_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_13_1111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_67_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_1096 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10795_ _00539_ clknet_leaf_298_clk rf_ram.memory\[55\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_183_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_171_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07275__A2 _03234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08472__A1 _01369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_170_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_152_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_87_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11416_ _01148_ clknet_leaf_48_clk rf_ram.memory\[80\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_1_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_169_3534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11347_ _01079_ clknet_leaf_264_clk cpu.immdec.imm30_25\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_22_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06786__A1 _02773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06015__B _01351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_1143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11278_ _01013_ clknet_leaf_243_clk net214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09724__A1 _04781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05854__B _01956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10229_ _02765_ _02844_ _05107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_33_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_1115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_182_3767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06538__A1 rf_ram.i_raddr\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_1137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_182_3778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_5_14__f_clk_I clknet_3_3_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold1 rf_ram_if.wdata1_r\[2\] net258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__05746__C1 _01646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_179_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05770_ _01963_ _01965_ _01494_ _01966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05761__A2 _01735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_1071 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_18_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_18_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07440_ rf_ram.memory\[36\]\[0\] _03337_ _03338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08456__I net98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_8_Right_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_57_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_92_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07371_ rf_ram.memory\[267\]\[0\] _03294_ _03295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_174_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_174_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09110_ rf_ram.memory\[94\]\[1\] _04387_ _04389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_174_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06322_ _01600_ _02511_ _02516_ _02517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_31_1277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09041_ rf_ram.memory\[104\]\[0\] _04346_ _04347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06253_ rf_ram.memory\[430\]\[1\] _01804_ _01805_ _02448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_72_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11610__I net90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09287__I _04004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05204_ cpu.state.init_done _01390_ _01341_ _01404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XTAP_TAPCELL_ROW_92_2106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08215__A1 _03798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_92_2117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06184_ _01769_ _02377_ _02378_ _02379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_170_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_142_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06226__B1 _01702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09963__A1 _04921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05135_ _01334_ _01337_ _01338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_0_1_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09943_ _04921_ _04929_ _04931_ _01206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_70_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_39_Right_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05985__C1 _01714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_110_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06529__A1 _02714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09874_ cpu.state.init_done _01418_ _04471_ _04889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08825_ _02828_ _04195_ _04213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_116_Left_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08756_ _04061_ _04170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_05968_ _02161_ _02163_ _01493_ _02164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_139_1183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input10_I i_dbus_rdt[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10089__A1 _05017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07707_ _03488_ _03503_ _03504_ _00396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08687_ _04057_ _04126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_68_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05899_ _02093_ _02094_ _01746_ _02095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_178_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07638_ _03455_ _03460_ _03461_ _00370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_165_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06701__A1 _02826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_48_Right_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_64_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07569_ rf_ram.memory\[357\]\[1\] _03416_ _03418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_165_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_101_2268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_181_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_101_2279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_165_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09308_ cpu.immdec.imm11_7\[1\] _04520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_63_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_75_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10580_ _00324_ clknet_leaf_162_clk rf_ram.memory\[362\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07257__A2 _03040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_81_1898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_125_Left_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_35_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10261__A1 _02819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06465__B1 _01624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09239_ rf_ram.memory\[319\]\[1\] _04468_ _04470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_185_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_16_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08206__A1 _03787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06614__I _02787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_1165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_1240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10013__A1 _04950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11201_ _00937_ clknet_leaf_45_clk rf_ram.memory\[86\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09954__A1 _04911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06768__A1 _02876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_57_Right_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_11132_ _00868_ clknet_leaf_74_clk rf_ram.memory\[114\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_147_3117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_147_3128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_164_3431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09557__I1 net50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11063_ _00800_ clknet_leaf_11_clk rf_ram.memory\[138\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_164_3442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_134_Left_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10014_ rf_ram.memory\[348\]\[1\] _04973_ _04975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07193__A1 _03161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_125_2714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_125_2725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_153_1114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06940__A1 _03018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_99_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_66_Right_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10916_ _00660_ clknet_leaf_16_clk rf_ram.memory\[178\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_157_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08693__A1 _04129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_157_958 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10847_ _00591_ clknet_leaf_310_clk rf_ram.memory\[533\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_156_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_143_Left_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_183_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10778_ _00522_ clknet_leaf_329_clk rf_ram.memory\[567\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_81_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_775 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05849__B _01350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_188_3910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_151_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1059 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_124_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_75_Right_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_23_875 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_184_3807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06759__A1 _02873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_184_3818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_152_Left_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06940_ _03018_ _03020_ _03022_ _00111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_158_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input2_I i_dbus_rdt[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05982__A2 _01640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_181_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06871_ rf_ram.memory\[302\]\[1\] _02973_ _02976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_59_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07184__A1 _02738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05822_ rf_ram.memory\[212\]\[0\] _01523_ _02018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08610_ net238 _04078_ _04079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_230_clk clknet_5_23__leaf_clk clknet_leaf_230_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_101_1293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09590_ _04697_ cpu.immdec.imm24_20\[0\] _04701_ _04702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__05734__A2 _01531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06931__A1 _03014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_84_Right_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_82_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08541_ net246 _03949_ _04034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05753_ _01372_ _01879_ _01948_ _01949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_49_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08472_ _01369_ _01378_ rf_ram.rdata\[1\] _03987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_05684_ rf_ram.memory\[398\]\[0\] _01770_ _01880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08684__A1 _04094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_161_Left_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_159_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05603__I _01613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07423_ _03326_ _03324_ _03327_ _00289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_46_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_46_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_175_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_63_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07354_ rf_ram.memory\[252\]\[0\] _03283_ _03284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_134_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08436__A1 _03953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10243__A1 _02825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06305_ rf_ram.memory\[169\]\[1\] _01664_ _02500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_128_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08987__A2 _04303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_297_clk clknet_5_7__leaf_clk clknet_leaf_297_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07285_ _02836_ _03083_ _03241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_73_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_182_1321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_93_Right_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_116_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09024_ net246 _04303_ _04336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06236_ _02422_ _02425_ _01660_ _02430_ _02431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_26_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_170_493 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05670__A1 _01850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09936__A1 _04918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08739__A2 _04158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06167_ _01603_ _02360_ _02361_ _02362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_130_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input58_I i_ibus_rdt[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06098_ rf_ram.memory\[278\]\[1\] _01687_ _01679_ rf_ram.memory\[279\]\[1\] _01678_
+ rf_ram.memory\[277\]\[1\] _02293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__05958__C1 _01655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09926_ _04400_ _04921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_141_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05973__A2 _01530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09857_ _01382_ _04871_ _02690_ _01391_ _04878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_77_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_142_3025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_142_3036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_1109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_221_clk clknet_5_22__leaf_clk clknet_leaf_221_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08808_ _04057_ _04202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_77_1255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09788_ rf_ram.memory\[76\]\[1\] _04834_ _04836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06922__A1 _02958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_103_2308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08739_ _01497_ _04158_ _04159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_103_2319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_120_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07478__A2 _02815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_83_1938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_120_2633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_83_1949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05513__I _01508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10701_ _00445_ clknet_leaf_81_clk rf_ram.memory\[432\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_138_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_165_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_153_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_181_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_154_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10632_ _00376_ clknet_leaf_93_clk rf_ram.memory\[386\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09475__I0 net88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_148_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10234__A1 _02737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_288_clk clknet_5_18__leaf_clk clknet_leaf_288_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_118_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_181_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10563_ _00307_ clknet_leaf_203_clk rf_ram.memory\[32\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_107_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_118_2584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_20_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_118_2595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10494_ _00238_ clknet_leaf_54_clk rf_ram.memory\[471\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_20_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_31_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11115_ _00851_ clknet_leaf_86_clk rf_ram.memory\[122\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_9_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11046_ _00783_ clknet_leaf_336_clk rf_ram.memory\[145\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07166__A1 _03157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_212_clk clknet_5_19__leaf_clk clknet_leaf_212_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08902__A2 _04038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06374__C1 _01625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06913__A1 _02975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06126__C1 _01773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08666__A1 _04097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_1063 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_878 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_177_3677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_177_3688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06141__A2 _01709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_89_1137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08418__A1 _03919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_172_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_279_clk clknet_5_17__leaf_clk clknet_leaf_279_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_15_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09091__A1 _04367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_41_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07070_ rf_ram.memory\[494\]\[1\] _03105_ _03107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_124_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07641__A2 _03089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_1182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06021_ _02212_ _02213_ _02214_ _02215_ _02216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_140_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_168_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_1034 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_1089 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07972_ _02868_ _03668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__05955__A2 _01661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09711_ net102 _04767_ _04768_ net103 _04784_ _04785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__09146__A2 _03035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06923_ rf_ram.memory\[278\]\[0\] _03010_ _03011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_87_2016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_203_clk clknet_5_24__leaf_clk clknet_leaf_203_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09642_ rf_ram.memory\[78\]\[1\] _04728_ _04730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06854_ _02839_ _02941_ _02964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06365__C1 _01968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06904__A1 _02894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_171_1022 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05805_ rf_ram.memory\[172\]\[0\] _01692_ _01516_ rf_ram.memory\[173\]\[0\] _01953_
+ rf_ram.memory\[175\]\[0\] _02001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_179_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09573_ _04687_ _01079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_78_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06785_ _02910_ _02915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__05183__A3 _01382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06380__A2 _02547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_65_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_65_1613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05736_ rf_ram.memory\[444\]\[0\] _01799_ _01931_ rf_ram.memory\[445\]\[0\] _01857_
+ rf_ram.memory\[447\]\[0\] _01932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_08524_ _03685_ _04023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__08657__A1 _02953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_1114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_1185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08455_ _01408_ _02694_ _01401_ _03972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05667_ _01633_ _01863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_92_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06132__A2 _01782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_1169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07406_ _03100_ _03135_ _03316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_148_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_956 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09457__I0 net78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08386_ rf_ram.memory\[189\]\[0\] _03927_ _03928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08409__A1 _03922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05598_ rf_ram.memory\[294\]\[0\] _01777_ _01778_ rf_ram.memory\[295\]\[0\] _01793_
+ rf_ram.memory\[293\]\[0\] _01794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_0_45_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10216__A1 _05078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07337_ _03260_ _03271_ _03273_ _00257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_163_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05489__B _01684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09082__A1 net239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07268_ _02737_ _03230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_131_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06219_ rf_ram.memory\[386\]\[1\] _01785_ _01786_ rf_ram.memory\[387\]\[1\] _02413_
+ _02414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_09007_ _02971_ _04303_ _04325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07199_ _02761_ _02941_ _03187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_131_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07396__A1 _03309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06199__A2 _01706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_113_2492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_1287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_6_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05946__A2 _01661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09909_ rf_ram.memory\[292\]\[1\] _04908_ _04910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07148__A1 _03123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05952__B _01601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08896__A1 _04237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05254__S0 _01376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06371__A2 _01606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_159_3341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_154_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_96_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_159_3352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07320__A1 _03257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_25_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_1034 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09448__I0 net74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11664_ net115 net187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_148_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10615_ _00359_ clknet_leaf_105_clk rf_ram.memory\[314\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_148_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_1110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09073__A1 _04364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_181_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_172_3585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_425 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11595_ _01327_ clknet_leaf_38_clk rf_ram.memory\[9\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_172_3596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10546_ _00290_ clknet_leaf_142_clk rf_ram.memory\[333\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_135_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08820__A1 net250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_133_2868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10477_ _00221_ clknet_leaf_101_clk rf_ram.memory\[422\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07387__A1 _03289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05418__I _01613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05937__A2 _01682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_159_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11029_ _00766_ clknet_leaf_2_clk rf_ram.memory\[150\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08887__A1 _03672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08729__I _04077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06347__C1 _01713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07633__I _03359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_1039 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_179_3717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06362__A2 _01958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06570_ rf_ram.memory\[201\]\[0\] _02753_ _02754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_144_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_176_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05521_ _01493_ _01717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_43_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_129_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08240_ _03823_ _03834_ _03836_ _00597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05452_ _01527_ _01642_ _01647_ _01648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XTAP_TAPCELL_ROW_60_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_60_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_117_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_117_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08171_ rf_ram.memory\[543\]\[1\] _03792_ _03794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_145_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05383_ rf_ram.memory\[546\]\[0\] _01544_ _01521_ rf_ram.memory\[547\]\[0\] _01517_
+ rf_ram.memory\[545\]\[0\] _01579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XANTENNA__09064__A1 _04334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07122_ rf_ram.memory\[487\]\[0\] _03139_ _03140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_125_460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07614__A2 _02984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08811__A1 _04202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_970 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_43_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07053_ rf_ram.memory\[390\]\[1\] _03094_ _03096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_63_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_179_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput100 net100 o_dbus_dat[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_141_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput111 net111 o_dbus_dat[21] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_06004_ _01495_ _02193_ _02198_ _02199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xoutput122 net122 o_dbus_dat[31] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_101_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput133 net133 o_dbus_sel[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_58_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput144 net144 o_ext_rs1[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput155 net155 o_ext_rs1[25] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_58_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput166 net166 o_ext_rs1[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput177 net177 o_ext_rs2[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput188 net188 o_ext_rs2[26] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__05389__B1 _01554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_5_7__f_clk clknet_3_1_0_clk clknet_5_7__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__05928__A2 _01863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput199 net199 o_ext_rs2[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__05328__I _01523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11002__CLK clknet_5_0__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07955_ rf_ram.memory\[481\]\[1\] _03656_ _03658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06906_ _02970_ _02998_ _02999_ _00100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08639__I _04061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07886_ rf_ram.memory\[462\]\[1\] _03613_ _03615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09625_ _04637_ _04720_ _04722_ _01096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06837_ rf_ram.memory\[286\]\[1\] _02950_ _02952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06353__A2 _01501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07550__A1 _03393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09556_ _04673_ _04674_ _04523_ _01075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06768_ _02876_ _02900_ _02902_ _00059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_78_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08507_ cpu.immdec.imm11_7\[0\] cpu.immdec.imm11_7\[1\] cpu.immdec.imm11_7\[4\] _04011_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_05719_ _01536_ _01915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__06105__A2 _01626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09487_ _02690_ _04622_ _04623_ _01057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06699_ _02820_ _02853_ _02854_ _00038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07302__A1 _03222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_175_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_22_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08438_ _03956_ _03958_ _03960_ _00671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07853__A2 _03234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_22_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_149_1322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_701 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05864__A1 _01951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_154_3260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09055__A1 _02794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08369_ rf_ram.memory\[185\]\[0\] _03916_ _03917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_135_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xwire249 _02751_ net249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_10400_ _00144_ clknet_leaf_300_clk rf_ram.memory\[216\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11380_ _01112_ clknet_leaf_232_clk cpu.bufreg2.o_sh_done_r vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__08802__A1 _04170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_115_2532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05616__A1 rf_ram.memory\[312\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_78_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10331_ _00075_ clknet_leaf_174_clk rf_ram.memory\[287\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_150_3179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_307_clk_I clknet_5_4__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output89_I net89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10262_ rf_ram.memory\[574\]\[1\] _05125_ _05127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07369__A1 _03292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_1096 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_178_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10193_ _05081_ _05083_ _05085_ _01302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08030__A2 _02992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05919__A2 _01799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08869__A1 _04234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07541__A1 _03319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06344__A2 _01662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_1000 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_1022 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_139_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_174_3625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_173_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_127_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_135_2908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_182_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11647_ net128 net200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_181_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_71_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput13 i_dbus_rdt[1] net13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_108_983 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09597__A2 net47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput24 i_dbus_rdt[2] net24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_25_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput35 i_ibus_rdt[10] net35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput46 i_ibus_rdt[21] net46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11578_ _01310_ clknet_leaf_56_clk rf_ram.memory\[442\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput57 i_ibus_rdt[31] net57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_123_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05857__B _01564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10529_ _00273_ clknet_leaf_217_clk rf_ram.memory\[250\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_172_Right_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_24_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_58_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_1282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_1184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_23_1146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05148__I _01350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_36_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_36_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07780__A1 _03521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06583__A2 _02764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_53_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07740_ rf_ram.memory\[378\]\[1\] _03522_ _03525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07363__I _03013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07671_ _03088_ _03481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_149_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09410_ _04578_ _04579_ _04539_ _04580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_88_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_1112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06622_ _02750_ _02793_ _02794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_34_1231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09341_ _04541_ _00993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06553_ _02728_ _02738_ _02739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08088__A2 _03729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06099__A1 _01675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05504_ _01694_ _01699_ _01620_ _01700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_47_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09272_ _01365_ _04495_ _04496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06484_ rf_ram.memory\[6\]\[1\] _01640_ _01503_ _02679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_7_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_99_2240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08223_ _03820_ _03825_ _03826_ _00590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_62_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05435_ _01530_ _01631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__09037__A1 _04331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_173_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_117_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08154_ rf_ram.memory\[546\]\[1\] _03781_ _03783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05366_ rf_ram.i_raddr\[3\] _01562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_0_132_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_95_2159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_884 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07105_ rf_ram.memory\[501\]\[0\] _03128_ _03129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05767__B _01956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08085_ _03721_ _03739_ _03740_ _00538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_30_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05297_ rf_ram.i_raddr\[3\] _01493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_141_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07036_ _02738_ _03083_ _03084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_101_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_2_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_1149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_73_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_110_2440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input40_I i_ibus_rdt[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_293_clk_I clknet_5_7__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_1279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08987_ net236 _04303_ _04313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07771__A1 _03524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07938_ rf_ram.memory\[457\]\[1\] _03645_ _03647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_98_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07869_ rf_ram.memory\[408\]\[0\] _03604_ _03605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_138_1078 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_27_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06326__A2 _01804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_27_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09608_ net249 _04507_ _04714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_74_1066 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10880_ _00624_ clknet_leaf_282_clk rf_ram.memory\[243\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_168_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_156_3300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_151_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_149_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09539_ _04648_ _04659_ _04662_ _04663_ _01069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_112_1207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09276__A1 _01364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_183_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_231_clk_I clknet_5_23__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07826__A2 _03559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05521__I _01493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_108_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_152_3219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11501_ _01233_ clknet_leaf_177_clk rf_ram.memory\[348\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_109_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09028__A1 _04334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_163_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_840 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11432_ _01164_ clknet_leaf_293_clk rf_ram.memory\[61\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_105_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_163_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_151_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_246_clk_I clknet_5_21__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_184_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_132_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_130_2805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_1135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11363_ _01095_ clknet_leaf_64_clk rf_ram.memory\[71\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_130_2816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08251__A2 _02954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10314_ _00058_ clknet_leaf_268_clk rf_ram.memory\[513\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11294_ _01027_ clknet_leaf_250_clk net87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_104_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10245_ rf_ram.memory\[264\]\[0\] _05116_ _05117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_167_3495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10176_ _05049_ _05072_ _05074_ _01296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06565__A2 _02748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07762__A1 _02775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05773__B1 _01953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_128_2767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_128_2778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06317__A2 _01631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_1133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_187_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_159_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_53_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_159_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_97_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_146_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06527__I _02713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_13_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_72_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_13_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_170_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_142_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05220_ cpu.immdec.imm31 _01418_ _01419_ _01420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_182_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_163_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05151_ cpu.immdec.imm19_12_20\[5\] _01354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_64_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_170_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_38_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_38_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_150_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_55_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05461__C1 _01656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08910_ rf_ram.memory\[125\]\[1\] _04263_ _04265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_55_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_90_2067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09890_ _04887_ _04896_ _04898_ _01186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_90_2078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_176_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08841_ rf_ram.memory\[134\]\[0\] _04222_ _04223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_104_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_139_1310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08772_ _02953_ _04152_ _04180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05984_ rf_ram.memory\[0\]\[0\] _01613_ _01525_ _02180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07723_ rf_ram.memory\[398\]\[1\] _03512_ _03514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07505__A1 _03356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06308__A2 _01501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07654_ rf_ram.memory\[386\]\[1\] _03469_ _03471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_177_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06605_ _02780_ _02781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_0_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07585_ _03422_ _03427_ _03428_ _00350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_76_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_1050 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09324_ rf_ram.memory\[109\]\[0\] _04530_ _04531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06536_ _01352_ _02721_ _01341_ _02722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_48_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05341__I _01536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05819__A1 _01600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09255_ cpu.genblk3.csr.mstatus_mpie _01356_ _04482_ _01341_ _04483_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_111_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06467_ rf_ram.memory\[16\]\[1\] _01682_ _01601_ _02662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_16_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_173_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08206_ _03787_ _03814_ _03815_ _00584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_32_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06492__A1 _02603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_172_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05418_ _01613_ _01614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_16_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09186_ _04431_ _04436_ _04437_ _00942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06398_ _01769_ _02591_ _02592_ _02593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_05349_ rf_ram.memory\[514\]\[0\] _01544_ _01540_ rf_ram.memory\[515\]\[0\] _01539_
+ rf_ram.memory\[513\]\[0\] _01545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_16_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08137_ rf_ram.memory\[54\]\[0\] _03772_ _03773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07268__I _02737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08068_ net236 _03729_ _03730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09981__A2 _02958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07019_ _03055_ _03072_ _03073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_149_3170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10030_ _04400_ _04985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__09733__A2 net14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_1099 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07744__A1 _03521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_145_3089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_169_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_1318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10932_ _00676_ clknet_leaf_254_clk rf_ram_if.rreq_r vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05960__B _01599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05507__B1 _01688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_123_2675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_170_clk_I clknet_5_31__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_123_2686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10863_ _00607_ clknet_leaf_31_clk rf_ram.memory\[205\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_79_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_1195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_137_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_50_clk_I clknet_5_12__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10794_ _00538_ clknet_leaf_297_clk rf_ram.memory\[55\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_39_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_185_clk_I clknet_5_28__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_81_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_65_clk_I clknet_5_8__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11415_ _01147_ clknet_leaf_48_clk rf_ram.memory\[80\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_152_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_169_3524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_169_3535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11346_ _01078_ clknet_leaf_260_clk cpu.immdec.imm30_25\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_22_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07983__A1 _03654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11277_ _01012_ clknet_leaf_245_clk net212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08511__B _01366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_33_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10228_ _05081_ _05104_ _05106_ _01316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09724__A2 net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_33_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_182_3768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_182_3779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_123_clk_I clknet_5_13__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05746__B1 _01810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_146_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xhold2 rf_ram_if.wdata0_r\[1\] net259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_10159_ _05046_ _05063_ _05064_ _01289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05210__A2 _01409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09488__A1 net87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08160__A1 _03757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_138_clk_I clknet_5_25__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_18_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_186_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_76_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_18_clk_I clknet_5_2__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_175_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07370_ _02781_ _03253_ _03294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_48_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_146_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05161__I cpu.state.genblk1.misalign_trap_sync_r vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06321_ _02512_ _02513_ _02514_ _02515_ _01978_ _02516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__09660__A1 net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_1289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06252_ _02435_ _02439_ _02443_ _02446_ _02447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_09040_ net250 _04339_ _04346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_155_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_3_5_0_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_142_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05203_ _01342_ cpu.bufreg2.o_sh_done_r cpu.state.init_done _01402_ _01403_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_111_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_170_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_92_2107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06183_ rf_ram.memory\[470\]\[1\] _01785_ _01786_ rf_ram.memory\[471\]\[1\] _01848_
+ rf_ram.memory\[469\]\[1\] _02378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__08215__A2 _03009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09412__A1 net246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05134_ _01335_ _01336_ _01337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_29_1174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_1005 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_1076 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_187_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09942_ rf_ram.memory\[33\]\[1\] _04929_ _04931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05985__B1 _01635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_70_1704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09873_ _02713_ _01413_ _03989_ _01179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_08824_ _04205_ _04210_ _04212_ _00805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_31_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05336__I _01531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08755_ _04167_ _04168_ _04169_ _00779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09479__A1 cpu.bufreg.i_sh_signed vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05967_ rf_ram.memory\[18\]\[0\] _01605_ _01624_ rf_ram.memory\[19\]\[0\] _02162_
+ _02163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_07706_ rf_ram.memory\[381\]\[0\] _03503_ _03504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05780__B _01923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_1123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08686_ _04097_ _04123_ _04125_ _00754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_68_1655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_1003 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_1059 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08151__A1 _02893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_105_2350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05898_ rf_ram.memory\[90\]\[0\] _01801_ _01646_ rf_ram.memory\[91\]\[0\] _01645_
+ rf_ram.memory\[89\]\[0\] _02094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_36_1145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_68_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07637_ rf_ram.memory\[406\]\[0\] _03460_ _03461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_178_775 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_85_1980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_165_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07568_ _03389_ _03416_ _03417_ _00344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_0_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_101_2269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09307_ _04466_ _04517_ _04519_ _00981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_118_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06519_ _02707_ _02708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_64_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07499_ rf_ram.memory\[324\]\[0\] _03374_ _03375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_36_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09651__A1 net98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_81_1899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09238_ _04463_ _04468_ _04469_ _00962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_output194_I net194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_146_1144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09169_ _04397_ _04425_ _04426_ _00936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_181_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11200_ _00936_ clknet_leaf_45_clk rf_ram.memory\[86\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09954__A2 _02946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_max_cap240_I _02888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11131_ _00867_ clknet_leaf_74_clk rf_ram.memory\[115\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_43_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_147_3118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05955__B _01503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_147_3129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output71_I net71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_164_3432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11062_ _00799_ clknet_leaf_31_clk rf_ram.memory\[13\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_164_3443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07717__A1 _03488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10013_ _04950_ _04973_ _04974_ _01233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_5_6__f_clk_I clknet_3_1_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08390__A1 _03892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_125_2715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_125_2726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_157_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_4_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05690__B _01746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_169_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10915_ _00659_ clknet_leaf_29_clk rf_ram.memory\[209\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09890__A1 _04887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_184_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_1065 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10846_ _00590_ clknet_leaf_299_clk rf_ram.memory\[533\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_27_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10777_ _00521_ clknet_leaf_307_clk rf_ram.memory\[568\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_109_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05259__A2 _01382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_137_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06805__I _02825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_1076 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_188_3900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_152_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_188_3911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_140_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06208__A1 _01674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_112_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_184_3808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07956__A1 _03654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_184_3819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11329_ _01061_ clknet_leaf_123_clk rf_ram.memory\[289\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05967__B1 _01624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05431__A2 _01626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_1071 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_1101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06870_ _02825_ _02975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_158_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07184__A2 _02806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05821_ net251 _01987_ _02016_ _02017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_08540_ _04026_ _04031_ _04033_ _00700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05752_ net252 _01908_ _01947_ _01948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__08133__A1 _03754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_386 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08471_ _02714_ _03986_ _00678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05683_ _01368_ _01845_ _01878_ _01879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__09881__A1 _03309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07422_ rf_ram.memory\[371\]\[1\] _03324_ _03327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05498__A2 _01692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_46_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_773 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_135_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_63_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_63_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07353_ _03055_ _02839_ _03283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09633__A1 _04524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11621__I net71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06304_ rf_ram.memory\[168\]\[1\] _01510_ _01956_ _02499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_122_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07284_ _03225_ _03238_ _03240_ _00237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_33_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09023_ _04334_ _04332_ _04335_ _00881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_170_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06235_ _02426_ _02427_ _02428_ _02429_ _01670_ _02430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_171_984 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_170_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_170_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_170_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06166_ rf_ram.memory\[486\]\[1\] _01623_ _01688_ rf_ram.memory\[487\]\[1\] _01702_
+ rf_ram.memory\[485\]\[1\] _02361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_40_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06097_ rf_ram.memory\[276\]\[1\] _01735_ _02292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_141_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05958__B1 _01653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05422__A2 _01617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09925_ _04918_ _04919_ _04920_ _01199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_102_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09856_ cpu.state.genblk1.misalign_trap_sync_r _01413_ _04877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_142_3026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08372__A1 _03887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_142_3037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08807_ _04170_ _04199_ _04201_ _00799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05186__A1 cpu.mem_bytecnt\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09787_ _04634_ _04834_ _04835_ _01145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_99_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06999_ _03050_ _03059_ _03060_ _00132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06922__A2 _03009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_1_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08738_ _01369_ _01496_ _04158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_103_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08124__A1 _03757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09321__C2 cpu.immdec.imm11_7\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08669_ _04094_ _04114_ _04115_ _00747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_83_1939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_120_2623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09872__A1 _04887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_120_2634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10700_ _00444_ clknet_leaf_81_clk rf_ram.memory\[432\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05489__A2 _01683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_166_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_166_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06150__A3 _02344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10631_ _00375_ clknet_leaf_115_clk rf_ram.memory\[405\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_119_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_181_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09475__I1 net89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_1284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06438__A1 _01903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10234__A2 _02946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_1314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10562_ _00306_ clknet_leaf_205_clk rf_ram.memory\[32\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_180_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_24_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_52_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05646__C1 _01668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_118_2585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10493_ _00237_ clknet_leaf_126_clk rf_ram.memory\[472\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_20_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_118_2596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09388__B1 _04564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_121_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11114_ _00850_ clknet_leaf_86_clk rf_ram.memory\[122\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_9_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06610__A1 _02748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11045_ _00782_ clknet_leaf_336_clk rf_ram.memory\[145\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_60_1293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08363__A1 _02991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06374__B1 _01678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08115__A1 _02751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_98_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06126__B1 _01848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09863__A1 _04837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_188_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_188_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_177_3678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_177_3689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_156_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_1127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10829_ _00573_ clknet_leaf_274_clk rf_ram.memory\[542\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_39_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09615__A1 _04634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_184_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_138_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_116_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_156_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_41_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_41_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_153_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_140_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_112_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06020_ rf_ram.memory\[554\]\[1\] _01532_ _01521_ rf_ram.memory\[555\]\[1\] _01517_
+ rf_ram.memory\[553\]\[1\] _02215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_26_1111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07929__A1 _03622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05595__B _01790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07971_ _03654_ _03665_ _03667_ _00497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09710_ _04781_ net6 _04784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_06922_ _02958_ _03009_ _03010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_184_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_87_2017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09641_ _04634_ _04728_ _04729_ _01105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06853_ _02930_ _02961_ _02963_ _00083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05168__A1 _01369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06365__B1 _01959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10161__A1 _05049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06904__A2 _02997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05804_ rf_ram.memory\[174\]\[0\] _01501_ _02000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_171_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09572_ cpu.immdec.imm30_25\[3\] _04686_ _04678_ _04687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_78_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_175_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06784_ _02876_ _02912_ _02914_ _00063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_136_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05614__I _01714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_65_1603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08523_ _03956_ _04020_ _04022_ _00694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05735_ _01626_ _01931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_37_1251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_65_1614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_701 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09854__A1 _01385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08657__A2 _03945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08454_ _01401_ _03970_ net126 _03971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_93_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05666_ rf_ram.memory\[478\]\[0\] _01543_ _01862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_175_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_148_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_1305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_148_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07405_ _03292_ _03313_ _03315_ _00283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_186_Right_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_135_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08385_ _02959_ _03903_ _03927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_92_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09457__I1 net79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05597_ _01617_ _01793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_73_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07336_ rf_ram.memory\[254\]\[1\] _03271_ _03273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05891__A2 _01719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09082__A2 _04339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07267_ _03225_ _03227_ _03229_ _00231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_131_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_116_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09006_ _04301_ _04322_ _04324_ _00875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06218_ rf_ram.memory\[385\]\[1\] _01787_ _02413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_131_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05643__A2 _01662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_147_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_44_1211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07198_ _03161_ _03184_ _03186_ _00205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_103_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06149_ _02340_ _02341_ _02342_ _02343_ _01658_ _02344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_130_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_112_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06053__C1 _01636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08593__A1 _02805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07396__A2 _02992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_113_2493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_6_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09908_ _04884_ _04908_ _04909_ _01193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08345__A1 _03887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09839_ rf_ram_if.rgnt _03984_ _02709_ _04868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_154_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05254__S1 _01375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_186_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09845__A1 _01413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_159_3342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_159_3353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06659__A1 _02820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_1237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_25_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05867__C1 _01636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_25_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11663_ net114 net186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_181_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_153_Right_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09448__I1 net75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_166_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10614_ _00358_ clknet_leaf_105_clk rf_ram.memory\[314\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_148_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05882__A2 _01922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11594_ _01326_ clknet_leaf_204_clk rf_ram.memory\[28\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_180_Left_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_172_3586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_141_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_172_3597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07084__A1 _03087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10545_ _00289_ clknet_leaf_153_clk rf_ram.memory\[371\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_106_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_130_clk clknet_5_24__leaf_clk clknet_leaf_130_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08820__A2 _04195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_106_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06831__A1 _02927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05634__A2 _01623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_133_2858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10476_ _00220_ clknet_leaf_101_clk rf_ram.memory\[422\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_133_2869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06304__B _01956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_159_1110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08336__A1 _03309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11028_ _00765_ clknet_leaf_327_clk rf_ram.memory\[150\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_95_1142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06347__B1 _01721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_197_clk clknet_5_28__leaf_clk clknet_leaf_197_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08887__A2 _02909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_172_1321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_179_3718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_154_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_87_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_176_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09836__A1 _04840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05520_ rf_ram.memory\[322\]\[0\] _01652_ _01713_ rf_ram.memory\[323\]\[0\] _01715_
+ rf_ram.memory\[321\]\[0\] _01716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_129_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05451_ rf_ram.memory\[380\]\[0\] _01644_ _01645_ rf_ram.memory\[381\]\[0\] _01646_
+ rf_ram.memory\[383\]\[0\] _01647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_118_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_60_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_172_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_60_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_120_Right_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_172_534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_1181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08170_ _03787_ _03792_ _03793_ _00570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_55_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05873__A2 _01989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05382_ rf_ram.memory\[544\]\[0\] _01524_ _01528_ _01578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_15_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_160_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07121_ _02829_ _02911_ _03139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_126_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_1109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_121_clk clknet_5_13__leaf_clk clknet_leaf_121_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_28_1206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06822__A1 _02909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07052_ _03087_ _03094_ _03095_ _00150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05625__A2 _01683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput101 net101 o_dbus_dat[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_88_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06003_ _02194_ _02195_ _02196_ _02197_ _01495_ _02198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_51_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput112 net112 o_dbus_dat[22] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_23_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput123 net123 o_dbus_dat[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput134 net134 o_dbus_we vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput145 net145 o_ext_rs1[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_58_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput156 net156 o_ext_rs1[26] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_58_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08575__A1 _04023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05609__I _01503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput167 net167 o_ext_rs1[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput178 net178 o_ext_rs2[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput189 net189 o_ext_rs2[27] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_11_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06050__A2 _01606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07954_ _03651_ _03656_ _03657_ _00490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08327__A1 _03884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06905_ rf_ram.memory\[2\]\[0\] _02998_ _02999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_138_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_188_clk clknet_5_29__leaf_clk clknet_leaf_188_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07885_ _03587_ _03613_ _03614_ _00464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_173_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06889__A1 _02975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09624_ rf_ram.memory\[71\]\[1\] _04720_ _04722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06836_ _02927_ _02950_ _02951_ _00078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_168_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05344__I _01520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09555_ cpu.immdec.imm7 _02709_ _04526_ _04674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06767_ rf_ram.memory\[513\]\[1\] _02900_ _02902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09827__A1 _03668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08506_ cpu.immdec.imm11_7\[2\] cpu.immdec.imm11_7\[3\] _04010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_77_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05718_ _01909_ _01910_ _01913_ _01914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_38_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09486_ _01375_ _04622_ _04623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_38_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06698_ rf_ram.memory\[523\]\[0\] _02853_ _02854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_66_849 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08437_ rf_ram.memory\[174\]\[1\] _03958_ _03960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_176_884 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_22_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05649_ _01600_ _01832_ _01844_ net253 _01845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_148_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_22_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_154_3250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08368_ _02983_ _03903_ _03916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_154_3261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09055__A2 _04339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwire239 _02893_ net239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__07066__A1 _03092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07319_ rf_ram.memory\[272\]\[0\] _03262_ _03263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_112_clk clknet_5_15__leaf_clk clknet_leaf_112_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08299_ rf_ram.memory\[244\]\[0\] _03872_ _03873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_61_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_115_2533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05616__A2 _01666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10330_ _00074_ clknet_leaf_174_clk rf_ram.memory\[287\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_132_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_1849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10261_ _02819_ _05125_ _05126_ _01329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_103_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05519__I _01714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10192_ rf_ram.memory\[238\]\[1\] _05083_ _05085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_160_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06041__A2 _01537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_179_clk clknet_5_29__leaf_clk clknet_leaf_179_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__10125__A1 net244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05682__C _01362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07541__A2 _02904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_185_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_174_3626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_1034 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_16_1165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_135_2909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05855__A2 _01515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11646_ net127 net199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_108_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput14 i_dbus_rdt[20] net14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07057__A1 _03087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput25 i_dbus_rdt[30] net25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_24_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_103_clk clknet_5_15__leaf_clk clknet_leaf_103_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xinput36 i_ibus_rdt[11] net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_52_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11577_ _01309_ clknet_leaf_56_clk rf_ram.memory\[442\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput47 i_ibus_rdt[22] net47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__06804__A1 _02927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput58 i_ibus_rdt[3] net58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06813__I _02800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10528_ _00272_ clknet_leaf_217_clk rf_ram.memory\[250\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_122_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_123_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06280__A2 _01940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10459_ _00203_ clknet_leaf_43_clk rf_ram.memory\[473\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_62_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05429__I _01624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08557__A1 _04026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_36_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05873__B _01783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_36_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05791__A1 _01351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07670_ _03458_ _03478_ _03480_ _00383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06621_ _02785_ _02792_ _02793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_172_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_149_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09809__A1 _04837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09340_ cpu.ctrl.pc _03991_ _04540_ net213 _04541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06552_ _02737_ _02738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_74_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05503_ rf_ram.memory\[338\]\[0\] _01687_ _01696_ rf_ram.memory\[339\]\[0\] _01698_
+ _01699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_34_1265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09271_ _01364_ cpu.genblk3.csr.mcause3_0\[1\] _04495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_157_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06483_ _02674_ _02675_ _02676_ _02677_ _01562_ _02678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_185_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_99_2230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_16_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08222_ rf_ram.memory\[533\]\[0\] _03825_ _03826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05434_ _01622_ _01628_ _01629_ _01630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_99_2241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05846__A2 _01649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_173_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_55_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_160_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08153_ _03754_ _03781_ _03782_ _00564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05365_ rf_ram.memory\[538\]\[0\] _01544_ _01540_ rf_ram.memory\[539\]\[0\] _01539_
+ rf_ram.memory\[537\]\[0\] _01561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_7_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06256__C1 _01811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08796__A1 _04170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07104_ _02915_ _03072_ _03128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_70_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_1220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08084_ rf_ram.memory\[55\]\[0\] _03739_ _03740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_67_1074 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05296_ _01492_ _00003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07035_ net235 _03083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_140_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06271__A2 _01735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06008__C1 _01555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08548__A1 net235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_105_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_110_2441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_73_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_1236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06023__A2 _01538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07220__A1 _03193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05783__B _01978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08986_ _04301_ _04310_ _04312_ _00867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input33_I i_dbus_rdt[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07937_ _03619_ _03645_ _03646_ _00484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10107__A1 _05014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_1170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07868_ _02991_ _03559_ _03604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_27_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09607_ _04643_ _01331_ _04681_ _01087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06819_ _02796_ _02735_ _02939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__05534__A1 _01674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07799_ rf_ram.memory\[415\]\[1\] _03560_ _03562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_39_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09538_ _04526_ net39 _04663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_156_3301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_183_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07287__A1 _03222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09469_ net84 net85 _04604_ _04611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_164_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_333_clk clknet_5_4__leaf_clk clknet_leaf_333_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_93_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11500_ _01232_ clknet_leaf_179_clk rf_ram.memory\[277\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_152_3209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_184_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_1040 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_163_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11431_ _01163_ clknet_leaf_291_clk rf_ram.memory\[61\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_7_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_149_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08787__A1 _03071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11362_ _01094_ clknet_leaf_257_clk cpu.decode.co_ebreak vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_104_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_130_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_130_2817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_1147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10313_ _00057_ clknet_leaf_267_clk rf_ram.memory\[514\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_81_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11293_ _01026_ clknet_leaf_133_clk rf_ram.memory\[299\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_131_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10244_ _02727_ _02958_ _05116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07211__A1 _02795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_167_3496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10175_ rf_ram.memory\[20\]\[1\] _05072_ _05074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_128_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_1210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_128_2779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_156_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08711__A1 _04126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_18_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_324_clk clknet_5_5__leaf_clk clknet_leaf_324_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_84_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05828__A2 _01804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_13_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_13_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11629_ net79 net152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05868__B _01684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_13_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05150_ _01352_ _01353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__06543__I cpu.immdec.imm11_7\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_1214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_38_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06253__A2 _01804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_38_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05159__I _01361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05461__B1 _01654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_55_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_55_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_90_2068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_90_2079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06005__A2 _01532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08840_ _02805_ _04195_ _04222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_85_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06410__C1 _01931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08771_ _04170_ _04177_ _04179_ _00785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_139_1322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05983_ rf_ram.memory\[4\]\[0\] _01643_ _01714_ rf_ram.memory\[5\]\[0\] _01635_ rf_ram.memory\[7\]\[0\]
+ _02179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XANTENNA_clkbuf_3_1_0_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07722_ _03488_ _03512_ _03513_ _00402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07653_ _03455_ _03469_ _03470_ _00376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_79_248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11624__I net74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06604_ _02779_ _02726_ _02780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA_clkbuf_leaf_306_clk_I clknet_5_5__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07584_ rf_ram.memory\[316\]\[0\] _03427_ _03428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_149_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06718__I _02865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09323_ net243 _04037_ _04530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06535_ cpu.immdec.imm11_7\[0\] _02721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07269__A1 _03230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_315_clk clknet_5_5__leaf_clk clknet_leaf_315_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_75_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_111_1241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09254_ _01356_ _01462_ _04481_ _04482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_06466_ _01903_ _02659_ _02660_ _02661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_146_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08205_ rf_ram.memory\[536\]\[0\] _03814_ _03815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_28_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05417_ _01508_ _01613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_160_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_526 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_32_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09185_ rf_ram.memory\[179\]\[0\] _04436_ _04437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06492__A2 _02630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06397_ rf_ram.memory\[92\]\[1\] _01711_ _01772_ rf_ram.memory\[93\]\[1\] _01773_
+ rf_ram.memory\[95\]\[1\] _02592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_44_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06229__C1 _01721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08769__A1 _04167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08136_ _03668_ _03009_ _03772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05348_ _01543_ _01544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_160_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_913 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07441__A1 _03323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08067_ _03692_ _03729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_31_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05279_ _01366_ _01475_ _01477_ cpu.o_wdata0 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_3_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_109_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07018_ _03071_ _03072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_102_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_149_3160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09194__A1 net236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_149_3171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06402__B _01707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_1077 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08941__A1 _04266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08969_ rf_ram.memory\[118\]\[1\] _04299_ _04302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_169_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10931_ _00675_ clknet_leaf_12_clk rf_ram.memory\[176\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_3_Left_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_123_2676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_169_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10862_ _00606_ clknet_leaf_30_clk rf_ram.memory\[205\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_123_2687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_184_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_1065 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_1076 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_140_2990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10793_ _00537_ clknet_leaf_325_clk rf_ram.memory\[560\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_306_clk clknet_5_5__leaf_clk clknet_leaf_306_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_82_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_1173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_183_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_137_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_137_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_10_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11414_ _01146_ clknet_leaf_21_clk rf_ram.memory\[76\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_169_3525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_169_3536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11345_ _01077_ clknet_leaf_260_clk cpu.immdec.imm30_25\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_120_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_186_3850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11276_ _01011_ clknet_leaf_246_clk net211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_24_1231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10227_ rf_ram.memory\[212\]\[1\] _05104_ _05106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_123_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_33_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06312__B _02004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05707__I _01525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_182_3769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10158_ rf_ram.memory\[44\]\[0\] _05063_ _05064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_94_1207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_50_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10089_ _05017_ _05019_ _05021_ _01262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09488__A2 _03989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05870__C _01620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_18_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_18_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_162_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06171__A1 _01527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_48_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_1149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08999__A1 _04298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06320_ rf_ram.memory\[178\]\[1\] _01856_ _01911_ rf_ram.memory\[179\]\[1\] _01931_
+ rf_ram.memory\[177\]\[1\] _02515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_127_320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_5_23__f_clk_I clknet_3_5_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_292_clk_I clknet_5_24__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_183_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06251_ _01909_ _02444_ _02445_ _02446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__10935__D cpu.o_wdata1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05202_ cpu.state.stage_two_req _01402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_115_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06182_ rf_ram.memory\[468\]\[1\] _01846_ _02377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_92_2108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_40_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09412__A2 _02801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06206__C _01717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07423__A1 _03326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06226__A2 _01634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05133_ cpu.decode.opcode\[2\] cpu.branch_op _01336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_0_40_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09941_ _04918_ _04929_ _04930_ _01205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_64_1099 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11619__I net69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_70_1705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09176__A1 _04401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_230_clk_I clknet_5_23__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09872_ _04887_ _04885_ _04888_ _01178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08923__A1 _04269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08823_ rf_ram.memory\[136\]\[1\] _04210_ _04212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05737__A1 _01909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08754_ rf_ram.memory\[146\]\[0\] _04168_ _04169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05966_ rf_ram.memory\[17\]\[0\] _01514_ _02162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__09479__A2 net89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07705_ _02960_ _03496_ _03503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_36_1102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_245_clk_I clknet_5_21__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08685_ rf_ram.memory\[155\]\[1\] _04123_ _04125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_174_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_105_2340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05897_ rf_ram.memory\[88\]\[0\] _01683_ _01684_ _02093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xclkbuf_leaf_92_clk clknet_5_11__leaf_clk clknet_leaf_92_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_135_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_68_1656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_1135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08151__A2 _03765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_68_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_1184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_105_2351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07636_ _03008_ _03089_ _03460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_85_1970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_85_1981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07567_ rf_ram.memory\[357\]\[0\] _03416_ _03417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_36_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09306_ rf_ram.memory\[63\]\[1\] _04517_ _04519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06518_ _01411_ _02707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_64_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07498_ _03319_ _02883_ _03374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_36_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09237_ rf_ram.memory\[319\]\[0\] _04468_ _04469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_145_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06465__A2 _01605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06449_ _01903_ _02642_ _02643_ _02644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_161_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_173_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09168_ rf_ram.memory\[86\]\[0\] _04425_ _04426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_16_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output187_I net187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_39_Left_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07414__A1 _03289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_146_1167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06217__A2 _01782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08119_ _03757_ _03759_ _03761_ _00551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_32_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_146_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09099_ _04364_ _04381_ _04382_ _00910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_11130_ _00866_ clknet_leaf_73_clk rf_ram.memory\[115\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_47_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_147_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09167__A1 _03008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11061_ _00798_ clknet_leaf_31_clk rf_ram.memory\[13\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_164_3433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06132__B _01783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_164_3444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10012_ rf_ram.memory\[348\]\[0\] _04973_ _04974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08390__A2 _02829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_125_2716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_125_2727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_48_Left_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_98_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_93_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_54_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_83_clk clknet_5_11__leaf_clk clknet_leaf_83_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_54_1235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_1246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10914_ _00658_ clknet_leaf_28_clk rf_ram.memory\[209\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_98_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06153__A1 _01597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_184_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10845_ _00589_ clknet_leaf_308_clk rf_ram.memory\[534\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_183_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_156_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10776_ _00520_ clknet_leaf_324_clk rf_ram.memory\[568\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_82_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07653__A1 _03455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_1310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06307__B _01564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_57_Left_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_70_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_188_3901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_188_3912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06026__C _01495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07405__A1 _03292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_849 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_184_3809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11328_ _01060_ clknet_leaf_123_clk rf_ram.memory\[289\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_22_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11259_ _00994_ clknet_leaf_250_clk net213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__05437__I _01508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_66_Left_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05820_ _01768_ _02003_ _02015_ _01569_ _02016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_94_1037 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_167_Right_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_167_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05751_ _01674_ _01934_ _01946_ _01569_ _01947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_82_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_74_clk clknet_5_10__leaf_clk clknet_leaf_74_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09330__A1 _04463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08470_ rf_ram_if.rreq_r _03986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_49_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05682_ _01674_ _01866_ _01877_ _01362_ _01878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_187_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_148_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09881__A2 _02795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_58_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07421_ _03017_ _03326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__07892__A1 _03590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_175_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_163_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_175_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_1032 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07352_ _03260_ _03280_ _03282_ _00263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_46_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_63_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_63_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_162_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09633__A2 net59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06303_ _02495_ _02497_ _01494_ _02498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XPHY_EDGE_ROW_75_Left_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_61_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06447__A2 _01536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07283_ rf_ram.memory\[472\]\[1\] _03238_ _03240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_73_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_155_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06217__B _01783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09022_ rf_ram.memory\[108\]\[1\] _04332_ _04335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06234_ rf_ram.memory\[402\]\[1\] _01500_ _01763_ rf_ram.memory\[403\]\[1\] _01656_
+ rf_ram.memory\[401\]\[1\] _02429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_143_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_116_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_1318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06165_ rf_ram.memory\[484\]\[1\] _01735_ _02360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_14_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06731__I _02825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06096_ _01368_ _02263_ _02290_ _02291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_09924_ rf_ram.memory\[342\]\[0\] _04919_ _04920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05347__I _01530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_84_Left_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09855_ _02713_ _01418_ _04876_ _01172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_TAPCELL_ROW_142_3027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08806_ rf_ram.memory\[13\]\[1\] _04199_ _04201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_142_3038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_184_clk_I clknet_5_29__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06998_ rf_ram.memory\[225\]\[0\] _03059_ _03060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05186__A2 _01385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09786_ rf_ram.memory\[76\]\[0\] _04834_ _04835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06383__A1 _01972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_1_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_134_Right_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_1_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08737_ _01369_ _04157_ _00773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05949_ rf_ram.memory\[62\]\[0\] _01530_ _02145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_68_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_64_clk_I clknet_5_8__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_65_clk clknet_5_8__leaf_clk clknet_leaf_65_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09321__A1 _04526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09321__B2 cpu.immdec.imm30_25\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_139_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08668_ rf_ram.memory\[157\]\[0\] _04114_ _04115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_68_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_120_2624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_96_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_120_2635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_113_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07619_ _02904_ _03390_ _03449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_199_clk_I clknet_5_25__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07883__A1 _02836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08599_ rf_ram.memory\[165\]\[0\] _04071_ _04072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10630_ _00374_ clknet_leaf_102_clk rf_ram.memory\[405\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_165_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_93_Left_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_49_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_76_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_79_clk_I clknet_5_11__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_147_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_91_530 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10561_ _00305_ clknet_leaf_163_clk rf_ram.memory\[367\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07635__A1 _03458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_122_clk_I clknet_5_15__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_162_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05646__B1 _01763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10492_ _00236_ clknet_leaf_126_clk rf_ram.memory\[472\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_106_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_118_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_20_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09388__A1 net216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_118_2597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_137_clk_I clknet_5_26__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11113_ _00849_ clknet_leaf_93_clk rf_ram.memory\[399\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_120_1104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_9_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_17_clk_I clknet_5_2__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11044_ _00781_ clknet_leaf_259_clk rf_ram_if.wen1_r vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08363__A2 _03903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_101_Right_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_157_1093 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_56_clk clknet_5_9__leaf_clk clknet_leaf_56_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08115__A2 _03729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_98_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_169_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_19_1196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_177_3679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_157_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10828_ _00572_ clknet_leaf_274_clk rf_ram.memory\[542\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_28_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_156_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05720__I _01550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07626__A1 _03422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06429__A2 _01641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10759_ _00503_ clknet_leaf_125_clk rf_ram.memory\[467\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_125_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_42_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_991 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_41_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_1145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07970_ rf_ram.memory\[47\]\[1\] _03665_ _03667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06921_ _03008_ _03009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_87_2007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_87_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09551__A1 _01391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06852_ rf_ram.memory\[285\]\[1\] _02961_ _02963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09640_ rf_ram.memory\[78\]\[0\] _04728_ _04729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_93_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05803_ _01996_ _01998_ _01564_ _01999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_117_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09571_ cpu.immdec.imm30_25\[4\] net53 _03967_ _04686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06783_ rf_ram.memory\[511\]\[1\] _02912_ _02914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_136_1144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09303__A1 _03668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_47_clk clknet_5_12__leaf_clk clknet_leaf_47_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08522_ rf_ram.memory\[188\]\[1\] _04020_ _04022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05734_ rf_ram.memory\[446\]\[0\] _01531_ _01930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_65_1604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_65_1615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_148_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08453_ _01418_ _02695_ _03970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_147_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_77_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05665_ _01855_ _01859_ _01860_ _01861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07865__A1 _03587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11632__I net82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07404_ rf_ram.memory\[247\]\[1\] _03313_ _03315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_93_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_175_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08384_ _03922_ _03924_ _03926_ _00651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_163_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05596_ rf_ram.memory\[292\]\[0\] _01735_ _01792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_46_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07335_ _03257_ _03271_ _03272_ _00256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_116_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_144_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08290__A1 _03852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07266_ rf_ram.memory\[196\]\[1\] _03227_ _03229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_143_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09005_ rf_ram.memory\[111\]\[1\] _04322_ _04324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_147_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06217_ rf_ram.memory\[384\]\[1\] _01782_ _01783_ _02412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_130_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07197_ rf_ram.memory\[474\]\[1\] _03184_ _03186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input63_I i_ibus_rdt[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_1223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06148_ rf_ram.memory\[312\]\[1\] _01666_ _01810_ rf_ram.memory\[313\]\[1\] _01811_
+ rf_ram.memory\[315\]\[1\] _02343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XANTENNA__08042__A1 _03686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_1159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06053__B1 _01610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_1267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08593__A2 _04067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_113_2494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06079_ _02271_ _02273_ _01620_ _02274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_111_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_6_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09907_ rf_ram.memory\[292\]\[0\] _04908_ _04909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09542__A1 _04478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09838_ cpu.state.cnt_r\[3\] _04866_ _04867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10152__A2 _02894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09769_ _04824_ _01138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_77_1098 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_38_clk clknet_5_7__leaf_clk clknet_leaf_38_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_150_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09845__A2 _03989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_159_3343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_159_3354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_178_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05867__B1 _01610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06636__I _02805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_25_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11662_ net113 net185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_126_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10613_ _00357_ clknet_leaf_156_clk rf_ram.memory\[354\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07608__A1 _02898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11593_ _01325_ clknet_leaf_210_clk rf_ram.memory\[28\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_137_2940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_172_3587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10544_ _00288_ clknet_leaf_153_clk rf_ram.memory\[371\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_36_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_991 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_107_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10475_ _00219_ clknet_leaf_103_clk rf_ram.memory\[423\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_150_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_133_2859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_150_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_159_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08336__A2 _02946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11027_ _00764_ clknet_leaf_2_clk rf_ram.memory\[151\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09533__A1 _04478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05715__I _01695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_179_3719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_1176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_29_clk clknet_5_1__leaf_clk clknet_leaf_29_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_91_1018 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07847__A1 _03590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_131_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_75_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_157_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_43_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_170_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_68_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05450_ _01635_ _01646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__05450__I _01635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_60_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_60_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05381_ rf_ram.memory\[548\]\[0\] _01538_ _01539_ rf_ram.memory\[549\]\[0\] _01540_
+ rf_ram.memory\[551\]\[0\] _01577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_28_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_172_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07120_ _03126_ _03136_ _03138_ _00175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_55_596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08272__A1 _03855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07051_ rf_ram.memory\[390\]\[0\] _03094_ _03095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_112_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06822__A2 _02941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06002_ rf_ram.memory\[514\]\[1\] _01544_ _01540_ rf_ram.memory\[515\]\[1\] _01539_
+ rf_ram.memory\[513\]\[1\] _02197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
Xoutput102 net102 o_dbus_dat[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput113 net113 o_dbus_dat[23] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput124 net124 o_dbus_dat[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__08024__A1 _03690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput135 net135 o_ext_funct3[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_2_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput146 net146 o_ext_rs1[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_58_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09772__A1 _04634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput157 net157 o_ext_rs1[27] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_58_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput168 net168 o_ext_rs1[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput179 net179 o_ext_rs2[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__05389__A2 _01544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07953_ rf_ram.memory\[481\]\[0\] _03656_ _03657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05794__C1 _01516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11627__I net77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06904_ _02894_ _02997_ _02998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_128_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06338__A1 _01972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07884_ rf_ram.memory\[462\]\[0\] _03613_ _03614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06230__B _01629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09623_ _04634_ _04720_ _04721_ _01095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06835_ rf_ram.memory\[286\]\[0\] _02950_ _02951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06766_ _02873_ _02900_ _02901_ _00058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09554_ cpu.immdec.imm31 _01491_ _01419_ _04673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_167_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05561__A2 _01755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09827__A2 _02917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05717_ rf_ram.memory\[438\]\[0\] _01706_ _01911_ rf_ram.memory\[439\]\[0\] _01912_
+ rf_ram.memory\[437\]\[0\] _01913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_08505_ _01369_ _01491_ _04009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07838__A1 _03554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09485_ _01411_ _03989_ _04621_ _04622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_06697_ _02781_ _02846_ _02853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_93_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_176_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_919 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08436_ _03953_ _03958_ _03959_ _00670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05648_ _01835_ _01838_ _01660_ _01843_ _01844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_110_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06510__A1 _01382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_22_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_163_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_50_1271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08367_ _03887_ _03913_ _03915_ _00645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_154_3251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05579_ _01769_ _01771_ _01774_ _01775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_46_563 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_154_3262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07318_ _02958_ _02946_ _03262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_61_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08263__A1 _03820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08298_ _03309_ _03135_ _03872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_150_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_1288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10070__A1 _04982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07249_ rf_ram.memory\[420\]\[1\] _03216_ _03218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_115_2534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10260_ rf_ram.memory\[574\]\[0\] _05125_ _05126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08015__A1 _02839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06124__C _01361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10191_ _05078_ _05083_ _05084_ _01301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_100_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05785__C1 _01857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06140__B _01707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10125__A2 _02832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_1172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05552__A2 _01543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_1160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_96_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_90_1062 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_1073 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_174_3616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_174_3627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06501__A1 cpu.ctrl.pc vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_166_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_166_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11645_ net126 net198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_83_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_126_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput15 i_dbus_rdt[21] net15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11576_ _01308_ clknet_leaf_29_clk rf_ram.memory\[211\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput26 i_dbus_rdt[31] net26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_25_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput37 i_ibus_rdt[12] net37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_91_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput48 i_ibus_rdt[23] net48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput59 i_ibus_rdt[4] net59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10527_ _00271_ clknet_leaf_140_clk rf_ram.memory\[267\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_52_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_165_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_21_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10458_ _00202_ clknet_leaf_44_clk rf_ram.memory\[473\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_122_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_161_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_1165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10389_ _00133_ clknet_leaf_273_clk rf_ram.memory\[225\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_58_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_36_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_36_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09506__A1 _04637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05791__A2 _01971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05445__I _01640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06620_ _02723_ _02757_ _02792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_177_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08756__I _04061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06740__A1 _02716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05543__A2 _01683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_137_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06551_ _02731_ _02736_ _02737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_90_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_1233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05502_ rf_ram.memory\[337\]\[0\] _01697_ _01698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_09270_ _04492_ _04493_ _04494_ _01485_ _00969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_87_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08493__A1 _02829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06482_ rf_ram.memory\[8\]\[1\] _01643_ _01714_ rf_ram.memory\[9\]\[1\] _01653_ rf_ram.memory\[11\]\[1\]
+ _02677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_158_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08221_ _03798_ _03072_ _03825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_185_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_16_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_99_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05433_ _01563_ _01629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_56_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_99_2242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05700__C1 _01608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08152_ rf_ram.memory\[546\]\[0\] _03781_ _03782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05364_ rf_ram.memory\[536\]\[0\] _01511_ _01552_ _01560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08245__A1 _03823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_911 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10052__A1 _04985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07103_ _03126_ _03124_ _03127_ _00169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06256__B1 _01810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09993__A1 _04950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08083_ _03668_ _03083_ _03739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_67_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_9_clk clknet_5_0__leaf_clk clknet_leaf_9_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_05295_ _01486_ _01490_ _01491_ _01492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_30_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_1037 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_5_15__f_clk clknet_3_3_0_clk clknet_5_15__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07034_ _02779_ _03007_ _03082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_3_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06008__B1 _01554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08548__A2 _04038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_110_2442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_73_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08985_ rf_ram.memory\[115\]\[1\] _04310_ _04312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09255__C _01341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05231__A1 cpu.bufreg.i_sh_signed vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07936_ rf_ram.memory\[457\]\[0\] _03645_ _03646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05355__I _01550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input26_I i_dbus_rdt[31] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07867_ _03590_ _03601_ _03603_ _00457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_138_1069 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_27_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09606_ _04712_ _04713_ _01086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_97_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06818_ _02930_ _02936_ _02938_ _00073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_35_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07798_ _03554_ _03560_ _03561_ _00430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_79_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09537_ cpu.csr_imm _04654_ _04662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06749_ _02888_ _02889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_93_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09468_ _04610_ _01051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_66_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_148_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06495__B1 _02462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08419_ rf_ram.memory\[29\]\[1\] _03946_ _03948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09399_ _04572_ _01020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_65_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_188_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_11_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08236__A1 _03798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11430_ _01162_ clknet_leaf_289_clk rf_ram.memory\[62\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_20_Left_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_11_1085 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10043__A1 _02812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06247__B1 _01925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11361_ _01093_ clknet_leaf_258_clk cpu.decode.op21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__08787__A2 _04152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06798__A1 _02873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_1321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06135__B _01790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_130_2807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10312_ _00056_ clknet_leaf_262_clk rf_ram.memory\[514\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_output94_I net94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_130_2818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11292_ _01025_ clknet_leaf_133_clk rf_ram.memory\[299\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_120_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09736__A1 _04781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10243_ _02825_ _05113_ _05115_ _01322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_30_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10174_ _05046_ _05072_ _05073_ _01295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07211__A2 _02941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_167_3497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05758__C1 _01953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05222__A1 _01385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05773__A2 _01958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_128_2769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_1109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_159_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06183__C1 _01848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06722__A1 _02866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_1075 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05930__C1 _01772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_186_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08475__A1 _01436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_127_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_13_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_13_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11628_ net78 net151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_53_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_154_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_128_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09975__A1 _02922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11559_ _01291_ clknet_leaf_112_clk rf_ram.memory\[448\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_25_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_94_2150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_38_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05997__C1 _01517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09727__A1 _04781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_55_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_90_2069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06410__B1 _01911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_260_clk clknet_5_17__leaf_clk clknet_leaf_260_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08770_ rf_ram.memory\[144\]\[1\] _04177_ _04179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05982_ rf_ram.memory\[6\]\[0\] _01640_ _01503_ _02178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_97_1057 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05764__A2 _01515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07721_ rf_ram.memory\[398\]\[0\] _03512_ _03513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_178_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07652_ rf_ram.memory\[386\]\[0\] _03469_ _03470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_177_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05516__A2 _01711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_137_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06603_ _01496_ _01498_ _02779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_76_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07583_ _02935_ _02839_ _03427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_149_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_177_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06534_ _01332_ _01366_ _01347_ _02720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_09322_ _04529_ _00986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_75_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_158_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07269__A2 _02899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_168_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09253_ _01366_ _01418_ _04481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_06465_ rf_ram.memory\[22\]\[1\] _01605_ _01624_ rf_ram.memory\[23\]\[1\] _01617_
+ rf_ram.memory\[21\]\[1\] _02660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_90_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_185_1310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_948 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_146_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05416_ _01603_ _01604_ _01611_ _01612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_08204_ _03798_ _02992_ _03814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_91_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_141_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09184_ net242 _04067_ _04436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_133_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06396_ rf_ram.memory\[94\]\[1\] _01770_ _02591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_32_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10025__A1 _04953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06229__B1 _01726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09966__A1 _04918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08135_ _03757_ _03769_ _03771_ _00557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_43_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05347_ _01530_ _01543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_160_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_44_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08066_ _03724_ _03726_ _03728_ _00531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05278_ _01381_ _01412_ _01476_ _01366_ _01477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_102_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_1051 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05452__A1 _01527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07017_ _02750_ _03007_ _03071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_105_1024 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_149_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_105_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09194__A2 _04418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_251_clk clknet_5_20__leaf_clk clknet_leaf_251_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08968_ _04061_ _04301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA_output132_I net132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07919_ _03622_ _03633_ _03635_ _00477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08899_ _04234_ _04257_ _04258_ _00834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_162_3394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10930_ _00674_ clknet_leaf_6_clk rf_ram.memory\[176\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05507__A2 _01623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06704__A1 _02820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_1131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_169_969 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_168_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10861_ _00605_ clknet_leaf_315_clk rf_ram.memory\[526\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_79_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_85_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_123_2677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_168_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_123_2688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_184_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_183_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_140_2991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_1088 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10792_ _00536_ clknet_leaf_323_clk rf_ram.memory\[560\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_148_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_1204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05969__B _01550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_93_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08209__A1 _03798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11413_ _01145_ clknet_leaf_21_clk rf_ram.memory\[76\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_151_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_90_981 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_169_3526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11344_ _01076_ clknet_leaf_260_clk cpu.immdec.imm30_25\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_169_3537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_162_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_104_Left_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_132_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_186_3840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_186_3851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11275_ _01010_ clknet_leaf_246_clk net210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07475__I _03359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05994__A2 _01502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_148_Right_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10226_ _05078_ _05104_ _05105_ _01315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_123_1179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07196__A1 _03157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_33_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_242_clk clknet_5_21__leaf_clk clknet_leaf_242_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10157_ _02787_ _02921_ _05063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__05746__A2 _01666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_50_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06943__A1 _03014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10088_ rf_ram.memory\[30\]\[1\] _05019_ _05021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_89_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08696__A1 _04126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_134_1220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_18_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_18_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05903__C1 _01715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_146_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08448__A1 _03956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_48_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07120__A1 _03126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_1258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06250_ rf_ram.memory\[444\]\[1\] _01799_ _01931_ rf_ram.memory\[445\]\[1\] _01857_
+ rf_ram.memory\[447\]\[1\] _02445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_26_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_182_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05201_ _01399_ _01400_ _01401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__09948__A1 _04921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05682__A1 _01674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06181_ _01600_ _02363_ _02375_ net253 _02376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_41_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_92_2109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05132_ cpu.decode.co_mem_word cpu.bne_or_bge cpu.csr_d_sel _01335_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__or3_2
XANTENNA__08620__A1 _02760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_1176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_744 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09940_ rf_ram.memory\[33\]\[0\] _04929_ _04930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05985__A2 _01661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_70_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_115_Right_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09871_ rf_ram.memory\[60\]\[1\] _04885_ _04888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_233_clk clknet_5_23__leaf_clk clknet_leaf_233_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08822_ _04202_ _04210_ _04211_ _00804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08753_ net236 _04152_ _04168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05965_ rf_ram.memory\[16\]\[0\] _01682_ _01601_ _02161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09479__A3 _03989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07704_ _03491_ _03500_ _03502_ _00395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_178_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_178_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08684_ _04094_ _04123_ _04124_ _00753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05896_ _01769_ _02090_ _02091_ _02092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_17_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_105_2341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_68_1657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_105_2352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07635_ _03458_ _03456_ _03459_ _00369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_68_1668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06162__A2 _01697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_85_1971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08439__A1 _02953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_85_1982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07566_ _02795_ _03390_ _03416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_177_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_165_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10246__A1 _02819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09305_ _04463_ _04517_ _04518_ _00980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_118_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06517_ _02703_ _02705_ _02706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05789__B _01928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07497_ _03360_ _03371_ _03373_ _00317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07111__A1 _03123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_180_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09236_ _03445_ _02909_ _04468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_17_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_145_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06448_ rf_ram.memory\[38\]\[1\] _01661_ _01607_ rf_ram.memory\[39\]\[1\] _01609_
+ rf_ram.memory\[37\]\[1\] _02643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XPHY_EDGE_ROW_17_Right_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_118_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06379_ _01768_ _02562_ _02573_ _01569_ _02574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_09167_ _03008_ _04418_ _04425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_31_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08118_ rf_ram.memory\[553\]\[1\] _03759_ _03761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_31_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09098_ rf_ram.memory\[96\]\[0\] _04381_ _04382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_47_1276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_744 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08049_ _03690_ _03715_ _03717_ _00525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05808__I _01504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11060_ _00797_ clknet_leaf_10_clk rf_ram.memory\[140\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09167__A2 _04418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_164_3434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07178__A1 _03161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_164_3445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10011_ _04911_ _02839_ _04973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_224_clk clknet_5_22__leaf_clk clknet_leaf_224_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_EDGE_ROW_26_Right_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05728__A2 _01922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_125_2717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_4_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10913_ _00657_ clknet_leaf_288_clk rf_ram.memory\[17\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_58_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07350__A1 _03257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_184_703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_156_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10844_ _00588_ clknet_leaf_312_clk rf_ram.memory\[534\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_67_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05900__A2 _01785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10775_ _00519_ clknet_leaf_294_clk rf_ram.memory\[56\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07102__A1 rf_ram.memory\[48\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_35_Right_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_94_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_171_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08850__A1 net241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_188_3902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_1089 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_112_Left_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_22_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08602__A1 _04062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05416__A1 _01603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11327_ _01059_ clknet_leaf_233_clk cpu.alu.cmp_r vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_127_1090 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_305_clk_I clknet_5_4__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05967__A2 _01605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11258_ _00993_ clknet_leaf_248_clk cpu.ctrl.pc vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XPHY_EDGE_ROW_44_Right_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07169__A1 _02915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_215_clk clknet_5_19__leaf_clk clknet_leaf_215_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10209_ net245 _03547_ _05095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_158_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11189_ _00925_ clknet_leaf_8_clk rf_ram.memory\[169\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_66_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06916__A1 _02970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_89_2060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_121_Left_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05195__A3 cpu.decode.opcode\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06392__A2 _01510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05750_ _01350_ _01939_ _01945_ _01946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__08669__A1 _04094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05453__I _01613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_530 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05681_ _01350_ _01871_ _01876_ _01877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_77_528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07420_ _03323_ _03324_ _03325_ _00288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_159_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_147_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09469__I0 net84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_53_Right_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10228__A1 _05081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07351_ rf_ram.memory\[26\]\[1\] _03280_ _03282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_63_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09094__A1 _04364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_63_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_1093 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_100_2260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06302_ rf_ram.memory\[162\]\[1\] _01958_ _01953_ rf_ram.memory\[163\]\[1\] _02496_
+ _02497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_31_1066 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07282_ _03222_ _03238_ _03239_ _00236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_155_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_80_1890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06233_ rf_ram.memory\[400\]\[1\] _01634_ _01903_ _02428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_31_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09021_ _04061_ _04334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_182_1313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_171_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06164_ _02356_ _02358_ _01620_ _02359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_06095_ _01350_ _02278_ _02289_ _01361_ _02290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_40_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_180_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06233__B _01903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_62_Right_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05958__A2 _01499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09923_ _04911_ _03009_ _04919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08004__I _02747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_206_clk clknet_5_24__leaf_clk clknet_leaf_206_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09854_ _01385_ _04487_ cpu.mem_bytecnt\[1\] _04876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08805_ _04167_ _04199_ _04200_ _00798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_142_3028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05791__C _01362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_142_3039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_1247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09785_ _02787_ _04507_ _04834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06997_ _03055_ _02899_ _03059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08736_ _02713_ _04156_ _03984_ _04157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XTAP_TAPCELL_ROW_1_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05948_ _02132_ _02136_ _02140_ _02143_ _02144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_1_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09321__A2 net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08667_ _02959_ _04078_ _04114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05879_ rf_ram.memory\[78\]\[0\] _01531_ _02075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07332__A1 _03260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_71_Right_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_120_2625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_166_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07618_ _03425_ _03446_ _03448_ _00363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08598_ _02794_ _04067_ _04071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07883__A2 _02972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_701 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07549_ rf_ram.memory\[35\]\[1\] _03404_ _03406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_113_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_165_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10560_ _00304_ clknet_leaf_162_clk rf_ram.memory\[367\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_118_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08832__A1 _04202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_1305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_1316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_162_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09219_ _03319_ _02960_ _04457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10491_ _00235_ clknet_leaf_98_clk rf_ram.memory\[417\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_134_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_20_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_118_2587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_118_2598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_20_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_80_Right_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_130_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05949__A2 _01530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06071__A1 _01675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11112_ _00848_ clknet_leaf_93_clk rf_ram.memory\[399\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_9_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_9_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11043_ _00780_ clknet_leaf_336_clk rf_ram.memory\[146\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05982__B _01503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08899__A1 _04234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_291_clk_I clknet_5_18__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07571__A1 _02935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06374__A2 _01677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_1061 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06126__A2 _01863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07323__A1 _03055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_1175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08584__I _04061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_157_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_45_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_157_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10827_ _00571_ clknet_leaf_312_clk rf_ram.memory\[543\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09076__A1 _04367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05222__B cpu.mem_bytecnt\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07626__A2 _03452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10758_ _00502_ clknet_leaf_125_clk rf_ram.memory\[467\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_27_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06037__C _01564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_41_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_666 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10689_ _00433_ clknet_leaf_82_clk rf_ram.memory\[435\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_113_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_1174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_164_1065 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_140_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_244_clk_I clknet_5_21__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_125_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_168_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05448__I _01643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06920_ _02773_ _03007_ _03008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA_clkbuf_leaf_259_clk_I clknet_5_17__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_87_2008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_87_2019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06851_ _02927_ _02961_ _02962_ _00082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06365__A2 _01940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05802_ rf_ram.memory\[170\]\[0\] _01989_ _01520_ rf_ram.memory\[171\]\[0\] _01997_
+ _01998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_09570_ _04680_ _04678_ _04685_ _01078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06782_ _02873_ _02912_ _02913_ _00062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_78_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_1231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08521_ _03953_ _04020_ _04021_ _00693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09303__A2 _02909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05733_ _01924_ _01927_ _01928_ _01929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_171_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_65_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_102_2300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_65_1616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07314__A1 _03257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_1106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_148_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08452_ _01369_ _01496_ _03969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_147_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05664_ _01563_ _01860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_93_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_82_1930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07403_ _03289_ _03313_ _03314_ _00282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05876__A1 _01600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_92_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05595_ _01784_ _01789_ _01790_ _01791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08383_ rf_ram.memory\[180\]\[1\] _03924_ _03926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_92_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09067__A1 _04331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_175_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_948 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06228__B _01615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07334_ rf_ram.memory\[254\]\[0\] _03271_ _03272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07617__A2 _03446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08814__A1 _04205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07265_ _03222_ _03227_ _03228_ _00230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_5_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_84_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_104_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09004_ _04298_ _04322_ _04323_ _00874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06216_ _02408_ _02410_ _01746_ _02411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_42_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07196_ _03157_ _03184_ _03185_ _00204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_14_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_1251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06147_ rf_ram.memory\[314\]\[1\] _01808_ _01650_ _02342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_42_995 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05358__I _01520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input56_I i_ibus_rdt[30] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06078_ rf_ram.memory\[338\]\[1\] _01687_ _01696_ rf_ram.memory\[339\]\[1\] _02272_
+ _02273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_TAPCELL_ROW_113_2495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09906_ _03445_ _02883_ _04908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_6_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09837_ cpu.mem_bytecnt\[1\] _01385_ cpu.state.o_cnt\[2\] _04866_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__09542__A2 net41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06356__A2 _01735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07553__A1 _03389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09768_ net122 _04766_ _04760_ _01439_ _04823_ _04824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_0_96_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08719_ _02983_ _04005_ _04146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_68_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06108__A2 _01543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09699_ _04776_ _01116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_95_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_166_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_159_3344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_159_3355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_25_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11661_ net112 net184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_25_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10612_ _00356_ clknet_leaf_160_clk rf_ram.memory\[354\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07608__A2 _03390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_166_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08805__A1 _04167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_181_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11592_ _01324_ clknet_leaf_139_clk rf_ram.memory\[264\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_37_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_137_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_1102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05619__A1 _01768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_172_3588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10543_ _00287_ clknet_leaf_143_clk rf_ram.memory\[334\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_135_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05977__B _01503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_1135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_1026 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10474_ _00218_ clknet_leaf_103_clk rf_ram.memory\[423\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_33_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09230__A1 net249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08579__I _04057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11026_ _00763_ clknet_leaf_328_clk rf_ram.memory\[151\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06347__A2 _01709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_1144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_179_3709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_1188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09297__A1 _04466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09049__A1 _04334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06048__B _01615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_60_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_172_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05380_ rf_ram.memory\[550\]\[0\] _01502_ _01506_ _01576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_60_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_144_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_153_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07050_ _02806_ _03089_ _03094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_183_clk_I clknet_5_29__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_1219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_97_2192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06001_ rf_ram.memory\[512\]\[1\] _01524_ _01528_ _02196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_140_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput103 net103 o_dbus_dat[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA_clkbuf_leaf_63_clk_I clknet_5_8__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09221__A1 _04431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput114 net114 o_dbus_dat[24] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput125 net125 o_dbus_dat[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput136 net136 o_ext_funct3[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput147 net147 o_ext_rs1[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_58_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_58_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_1100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput158 net158 o_ext_rs1[28] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput169 net169 o_ext_rs1[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__07783__A1 net237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_198_clk_I clknet_5_28__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07952_ _02898_ _03158_ _03656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05794__B1 _01520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_78_clk_I clknet_5_11__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06903_ _02996_ _02997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_177_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07883_ _02836_ _02972_ _03613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07535__A1 _03393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_1218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_121_clk_I clknet_5_13__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09622_ rf_ram.memory\[71\]\[0\] _04720_ _04721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_128_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06834_ _02917_ _02941_ _02950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_97_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09553_ _04654_ _04671_ _04672_ _01074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06765_ rf_ram.memory\[513\]\[0\] _02900_ _02901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09288__A1 net238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08504_ _03956_ _04006_ _04008_ _00689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05716_ _01626_ _01912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_66_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09484_ _04620_ _01384_ _01387_ _03989_ _04621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_77_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06696_ _02826_ _02850_ _02852_ _00037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_leaf_136_clk_I clknet_5_26__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08435_ rf_ram.memory\[174\]\[0\] _03958_ _03959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_109_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_175_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05647_ _01839_ _01840_ _01841_ _01842_ _01670_ _01843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_19_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06510__A2 cpu.decode.opcode\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_1115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_16_clk_I clknet_5_2__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08366_ rf_ram.memory\[184\]\[1\] _03913_ _03915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05578_ rf_ram.memory\[300\]\[0\] _01711_ _01772_ rf_ram.memory\[301\]\[0\] _01773_
+ rf_ram.memory\[303\]\[0\] _01774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_0_92_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_154_3252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_1283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_184_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_154_3263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_135_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_1245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07317_ _03260_ _03258_ _03261_ _00249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_46_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08297_ _03855_ _03869_ _03871_ _00619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_117_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07248_ _03190_ _03216_ _03217_ _00224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_115_2535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_131_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_61_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08015__A2 _03693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_42_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07179_ _02899_ _02997_ _03175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_output162_I net162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10190_ rf_ram.memory\[238\]\[0\] _05083_ _05084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07774__A1 _03521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05785__B1 _01931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06329__A2 _01515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_1140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_69_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_139_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06647__I _02814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_174_3617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_174_3628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_96_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_182_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11644_ cpu.bufreg2.o_sh_done_r net197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_126_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11575_ _01307_ clknet_leaf_29_clk rf_ram.memory\[211\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_64_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput16 i_dbus_rdt[22] net16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput27 i_dbus_rdt[3] net27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_123_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_25_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06265__A1 net252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput38 i_ibus_rdt[13] net38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_107_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10526_ _00270_ clknet_leaf_140_clk rf_ram.memory\[267\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput49 i_ibus_rdt[24] net49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_107_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05473__C1 _01668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09203__A1 _04434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10457_ _00201_ clknet_leaf_45_clk rf_ram.memory\[198\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_32_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_62_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10388_ _00132_ clknet_leaf_274_clk rf_ram.memory\[225\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_62_1165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_1296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_1176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_36_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06331__B _01978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05726__I _01536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07517__A1 _03360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11009_ _00746_ clknet_leaf_1_clk rf_ram.memory\[158\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_5_17__f_clk_I clknet_3_4_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_133_1115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06557__I _02742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06550_ cpu.immdec.imm11_7\[2\] _02730_ _02735_ _02736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_34_1223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_987 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_142_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_59_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05501_ _01514_ _01697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_06481_ rf_ram.memory\[10\]\[1\] _01686_ _01525_ _02676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08493__A2 _03496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_1109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08220_ _03823_ _03821_ _03824_ _00589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05432_ rf_ram.memory\[362\]\[0\] _01623_ _01625_ rf_ram.memory\[363\]\[0\] _01627_
+ _01628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_90_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_184_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05700__B1 _01702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_16_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_99_2232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_99_2243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_145_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_458 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05363_ rf_ram.memory\[540\]\[0\] _01538_ _01555_ rf_ram.memory\[541\]\[0\] _01554_
+ rf_ram.memory\[543\]\[0\] _01559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_08151_ _02893_ _03765_ _03781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_172_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07102_ rf_ram.memory\[48\]\[1\] _03124_ _03127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_160_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05294_ _01409_ _01491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_08082_ _03724_ _03736_ _03738_ _00537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_28_1005 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07033_ _03053_ _03079_ _03081_ _00145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_114_989 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_110_2432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07756__A1 _03524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_73_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06559__A2 _02743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_1318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11638__I net89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_73_1759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_110_2443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_1287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08984_ _04298_ _04310_ _04311_ _00866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06241__B _01916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05231__A2 net134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07935_ _02752_ _02832_ _03645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07508__A1 _03319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07866_ rf_ram.memory\[42\]\[1\] _03601_ _03603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08181__A1 _03787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09605_ _04524_ net49 _04701_ cpu.immdec.imm24_20\[4\] _04713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_78_1194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06817_ rf_ram.memory\[288\]\[1\] _02936_ _02938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_921 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input19_I i_dbus_rdt[25] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_27_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07797_ rf_ram.memory\[415\]\[0\] _03560_ _03561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_39_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09536_ _04653_ _04659_ _04660_ _04661_ _01068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06748_ _02779_ _02887_ _02888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_79_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_149_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09467_ net83 net84 _04604_ _04610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_164_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06679_ rf_ram.memory\[476\]\[0\] _02840_ _02841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_65_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_164_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_159_Left_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06495__A1 _01371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08418_ _03919_ _03946_ _03947_ _00664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_93_456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09398_ net221 _04561_ _04564_ net222 _04572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_93_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_163_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08349_ rf_ram.memory\[181\]\[0\] _03904_ _03905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_163_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08236__A2 _02923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_123_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06416__B _01916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_129_Right_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_73_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10043__A2 _03158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11360_ _01092_ clknet_leaf_257_clk cpu.decode.op22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_130_2808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10311_ _00055_ clknet_leaf_271_clk rf_ram.memory\[515\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_85_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_130_2819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11291_ _00006_ clknet_leaf_239_clk cpu.ctrl.pc_plus_offset_cy_r vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_131_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output87_I net87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10242_ rf_ram.memory\[213\]\[1\] _05113_ _05115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07747__A1 _02983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_168_Left_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05758__B1 _01516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10173_ rf_ram.memory\[20\]\[0\] _05072_ _05073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_100_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_167_3487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_167_3498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05990__B _01372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08172__A1 _03790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06183__B1 _01786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06722__A2 _02869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05930__B1 _01857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_177_Left_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_84_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_5_21__f_clk clknet_3_5_0_clk clknet_5_21__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_85_946 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_840 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06486__A1 rf_ram.memory\[0\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_166_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08592__I _03902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_182_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_170_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11627_ net77 net150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_53_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11558_ _01290_ clknet_leaf_127_clk rf_ram.memory\[44\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09975__A2 _03253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_94_2140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07986__A1 _03651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_94_2151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10509_ _00253_ clknet_leaf_217_clk rf_ram.memory\[255\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_111_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_38_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05997__B1 _01521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11489_ _01221_ clknet_leaf_189_clk rf_ram.memory\[275\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_186_Left_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05461__A2 _01652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06840__I _02953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09727__A2 net11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_55_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07738__A1 _03521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06061__B _01658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05456__I _01499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05213__A2 cpu.mem_bytecnt\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05981_ _02173_ _02174_ _02175_ _02176_ _01562_ _02177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_07720_ _02971_ _03481_ _03512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_100_1169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07671__I _03088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07651_ net239 _03089_ _03469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07910__A1 _02822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06602_ _02748_ _02776_ _02778_ _00017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07582_ _03425_ _03423_ _03426_ _00349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_48_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09321_ _04526_ net36 _04521_ cpu.immdec.imm30_25\[0\] _04522_ cpu.immdec.imm11_7\[4\]
+ _04529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_76_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06533_ _02717_ _02718_ _02719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_4
XANTENNA__08466__A2 _01364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09663__A1 net120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06477__A1 _01903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09252_ cpu.genblk3.csr.mstatus_mie _04480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_91_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_47_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06464_ rf_ram.memory\[20\]\[1\] _01536_ _02659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_157_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_185_1322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05685__C1 _01773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08203_ _03790_ _03811_ _03813_ _00583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05415_ rf_ram.memory\[358\]\[0\] _01606_ _01608_ rf_ram.memory\[359\]\[0\] _01610_
+ rf_ram.memory\[357\]\[0\] _01611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XTAP_TAPCELL_ROW_151_3200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_16_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09183_ _04434_ _04432_ _04435_ _00941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06395_ _02578_ _02582_ _02586_ _02589_ _02590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__06236__B _01660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_141_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08134_ rf_ram.memory\[550\]\[1\] _03769_ _03771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_161_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05346_ rf_ram.memory\[512\]\[0\] _01524_ _01528_ _01542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_71_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07977__A1 _03654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08065_ rf_ram.memory\[563\]\[1\] _03726_ _03728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05277_ _01381_ _01426_ _01476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_113_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07016_ _03053_ _03068_ _03070_ _00139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07729__A1 _03491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_149_3162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05366__I rf_ram.i_raddr\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08967_ _04298_ _04299_ _04300_ _00860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07918_ rf_ram.memory\[45\]\[1\] _03633_ _03635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08898_ rf_ram.memory\[429\]\[0\] _04257_ _04258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_162_3395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07849_ rf_ram.memory\[410\]\[0\] _03592_ _03593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_169_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10860_ _00604_ clknet_leaf_315_clk rf_ram.memory\[526\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_155_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05912__B1 _01857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_123_2678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_151_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_123_2689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_156_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09519_ _01399_ cpu.decode.opcode\[1\] _01450_ _04647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_17_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_1142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_140_2992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10791_ _00535_ clknet_leaf_332_clk rf_ram.memory\[561\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_52_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_93_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_164_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08209__A2 _03083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11412_ _01144_ clknet_leaf_18_clk rf_ram.memory\[187\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10016__A2 _02984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05691__A2 _01782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11343_ _01075_ clknet_leaf_236_clk cpu.immdec.imm7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_169_3527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_169_3538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06660__I _02747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_186_3841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11274_ _01009_ clknet_leaf_246_clk net209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_120_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_186_3852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_1147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10225_ rf_ram.memory\[212\]\[0\] _05104_ _05105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10182__I _02742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10156_ _05049_ _05060_ _05062_ _01288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_50_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10087_ _05014_ _05019_ _05020_ _01261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08145__A1 _03757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1020 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09893__A1 _04884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_187_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_18_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_18_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05903__B1 _01654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_1107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_70_1231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_174_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09645__A1 cpu.mem_bytecnt\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_1242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10989_ _00726_ clknet_leaf_28_clk rf_ram.memory\[129\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_29_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_48_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06459__A1 rf_ram.memory\[48\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_183_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_142_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05200_ cpu.decode.co_mem_word _01400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
X_06180_ _02366_ _02369_ _01660_ _02374_ _02375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_128_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_170_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07959__A1 _03651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05131_ _01333_ cpu.decode.op26 cpu.decode.co_ebreak _01334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_41_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08620__A2 _02881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_1057 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06092__C1 _01713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09870_ _04400_ _04887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_70_1707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08384__A1 _03922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08821_ rf_ram.memory\[136\]\[0\] _04210_ _04211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_110_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10191__A1 _05078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08752_ _04057_ _04167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_05964_ _01903_ _02158_ _02159_ _02160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__08136__A1 _03668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_144_3070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07703_ rf_ram.memory\[400\]\[1\] _03500_ _03502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08683_ rf_ram.memory\[155\]\[0\] _04123_ _04124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_139_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05895_ rf_ram.memory\[92\]\[0\] _01711_ _01772_ rf_ram.memory\[93\]\[0\] _01773_
+ rf_ram.memory\[95\]\[0\] _02091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_07634_ rf_ram.memory\[388\]\[1\] _03456_ _03459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_152_1321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_68_1658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_105_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_68_1669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_105_2353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_85_1972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07565_ _03393_ _03413_ _03415_ _00343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_85_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09636__A1 _04524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08439__A2 _03949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11651__I net101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09304_ rf_ram.memory\[63\]\[0\] _04517_ _04518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06516_ cpu.bufreg.c_r _02704_ _02705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_07496_ rf_ram.memory\[364\]\[1\] _03371_ _03373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_146_631 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09235_ _04466_ _04464_ _04467_ _00961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_134_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06447_ rf_ram.memory\[36\]\[1\] _01536_ _02642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_118_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_173_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_12_1181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09939__A2 _02899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09166_ _04401_ _04422_ _04424_ _00935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05673__A2 _01719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06378_ _01600_ _02567_ _02572_ _02573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_43_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08117_ _03754_ _03759_ _03760_ _00550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_121_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05329_ rf_ram.i_raddr\[2\] _01525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_142_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_701 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09097_ net237 _04339_ _04381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_160_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_142_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07576__I _03355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06622__A1 _02750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08048_ rf_ram.memory\[566\]\[1\] _03715_ _03717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_47_1288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_164_3435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10010_ _04953_ _04970_ _04972_ _01232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_164_3446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06386__B1 _01925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09999_ rf_ram.memory\[276\]\[1\] _04964_ _04966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_181_3760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_125_2718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_153_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09875__A1 _02713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06689__A1 _02820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10912_ _00656_ clknet_leaf_288_clk rf_ram.memory\[17\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_39_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_157_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10843_ _00587_ clknet_leaf_299_clk rf_ram.memory\[535\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09627__A1 _04643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_184_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10774_ _00518_ clknet_leaf_294_clk rf_ram.memory\[56\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_82_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_181_Right_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_leaf_160_clk clknet_5_27__leaf_clk clknet_leaf_160_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_137_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08850__A2 _04195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_180_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06861__A1 _02927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_1292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_188_3903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_152_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_1322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_152_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11326_ _00004_ clknet_leaf_255_clk cpu.bufreg.c_r vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06613__A1 _02716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06323__C _01569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11257_ _00992_ clknet_leaf_77_clk rf_ram.memory\[99\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_63_1090 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07169__A2 _02954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10208_ _05081_ _05092_ _05094_ _01308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_66_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11188_ _00924_ clknet_leaf_9_clk rf_ram.memory\[169\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_140_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_1310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10139_ _05046_ _05051_ _05052_ _01281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_59_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_89_2050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_89_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_101_1286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_1305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05680_ _01872_ _01873_ _01874_ _01875_ _01717_ _01876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_49_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_187_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09618__A1 _04643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_159_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_1181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_1061 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07350_ _03257_ _03280_ _03281_ _00262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_175_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_174_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_100_2250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_63_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_100_2261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06301_ rf_ram.memory\[161\]\[1\] _01664_ _02496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_46_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_63_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07281_ rf_ram.memory\[472\]\[0\] _03238_ _03239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_151_clk clknet_5_26__leaf_clk clknet_leaf_151_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_72_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_80_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_80_1891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09020_ _04331_ _04332_ _04333_ _00880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06232_ rf_ram.memory\[404\]\[1\] _01509_ _01668_ rf_ram.memory\[405\]\[1\] _01763_
+ rf_ram.memory\[407\]\[1\] _02427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XANTENNA__05655__A2 _01782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_170_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06163_ rf_ram.memory\[482\]\[1\] _01687_ _01696_ rf_ram.memory\[483\]\[1\] _02357_
+ _02358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_142_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06065__C1 _01664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06604__A1 _02779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06094_ _01349_ _02283_ _02288_ _02289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_111_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_141_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05812__C1 _01773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06080__A2 _01537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09922_ _04396_ _04918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_146_3110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08357__A1 _03887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09853_ _02713_ _04875_ _01171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10164__A1 _05046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_1099 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08804_ rf_ram.memory\[13\]\[0\] _04199_ _04200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_147_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09784_ _04637_ _04831_ _04833_ _01144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_142_3029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06996_ _03053_ _03056_ _03058_ _00131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08109__A1 net247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08735_ _03968_ _04156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05947_ _01903_ _02141_ _02142_ _02143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_1_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09857__A1 _01382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_1_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_178_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_178_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08666_ _04097_ _04111_ _04113_ _00746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05878_ _01368_ _02046_ _02073_ _01597_ _02074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_139_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07617_ rf_ram.memory\[313\]\[1\] _03446_ _03448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_120_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08597_ _04062_ _04068_ _04070_ _00720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_72_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_166_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_178_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10219__A2 _03082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07548_ _03389_ _03404_ _03405_ _00336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05894__A2 _01770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_1243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_36_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06408__C _01362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07096__A1 _03092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07479_ rf_ram.memory\[328\]\[0\] _03362_ _03363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_142_clk clknet_5_27__leaf_clk clknet_leaf_142_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_118_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_174_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09218_ _04434_ _04454_ _04456_ _00955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_118_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06843__A1 _02927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05646__A2 _01500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10490_ _00234_ clknet_leaf_95_clk rf_ram.memory\[417\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_84_1219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output192_I net192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_20_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09149_ rf_ram.memory\[8\]\[1\] _04412_ _04414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_118_2588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06424__B _02004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_114_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_183_3800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11111_ _00847_ clknet_leaf_86_clk rf_ram.memory\[123\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_31_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_9_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08348__A1 _03071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11042_ _00779_ clknet_leaf_336_clk rf_ram.memory\[146\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08899__A2 _04257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07571__A2 _02960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_169_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07323__A2 _02909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10826_ _00570_ clknet_leaf_312_clk rf_ram.memory\[543\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_45_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_45_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_184_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_172_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07087__A1 _02775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_171_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10757_ _00501_ clknet_leaf_123_clk rf_ram.memory\[478\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_133_clk clknet_5_24__leaf_clk clknet_leaf_133_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_109_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06834__A1 _02917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05637__A2 _01631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10688_ _00432_ clknet_leaf_81_clk rf_ram.memory\[435\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_129_1142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_125_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_164_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_35_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_125_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08587__A1 _02828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05729__I _01695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_1125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_1039 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06062__A2 _01662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11309_ _01042_ clknet_leaf_266_clk net74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_61_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09645__B _01375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10146__A1 _05049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07011__A1 _03053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_87_2009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_184_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06850_ rf_ram.memory\[285\]\[0\] _02961_ _02962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05464__I _01599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_172_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05801_ rf_ram.memory\[169\]\[0\] _01664_ _01997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06781_ rf_ram.memory\[511\]\[0\] _02912_ _02913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08520_ rf_ram.memory\[188\]\[0\] _04020_ _04021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05732_ _01563_ _01928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_136_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_78_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_65_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08511__A1 _03989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_102_2301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_65_1617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08451_ _02714_ _03968_ _00676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05663_ rf_ram.memory\[474\]\[0\] _01856_ _01857_ rf_ram.memory\[475\]\[0\] _01858_
+ _01859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_33_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_82_1920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_82_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07402_ rf_ram.memory\[247\]\[0\] _03313_ _03314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_19_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08382_ _03919_ _03924_ _03925_ _00650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_9_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05594_ _01493_ _01790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_58_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07333_ _03055_ _02917_ _03271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_116_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_124_clk clknet_5_13__leaf_clk clknet_leaf_124_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_27_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_144_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_740 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07264_ rf_ram.memory\[196\]\[0\] _03227_ _03228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_27_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_14_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_738 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_147_1242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09003_ rf_ram.memory\[111\]\[0\] _04322_ _04323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06215_ rf_ram.memory\[394\]\[1\] _01777_ _01778_ rf_ram.memory\[395\]\[1\] _02409_
+ _02410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_131_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07195_ rf_ram.memory\[474\]\[0\] _03184_ _03185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_115_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06244__B _01790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_41_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_77_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06146_ rf_ram.memory\[316\]\[1\] _01724_ _01725_ rf_ram.memory\[317\]\[1\] _01726_
+ rf_ram.memory\[319\]\[1\] _02341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_14_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07250__A1 _03193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06053__A2 _01644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_884 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06077_ rf_ram.memory\[337\]\[1\] _01697_ _02272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__09555__B _04526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_113_2496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09905_ _04887_ _04905_ _04907_ _01192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_6_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input49_I i_ibus_rdt[24] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05800__A2 _01510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10137__A1 _02794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07002__A1 _03055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09836_ _04840_ _04863_ _04865_ _01164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06979_ _02775_ _03040_ _03047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09767_ _04804_ net26 _04823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_38_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08718_ _04129_ _04143_ _04145_ _00766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09698_ net129 _04767_ _04768_ net99 _04775_ _04776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
Xclkbuf_5_2__f_clk clknet_3_0_0_clk clknet_5_2__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08502__A1 _03953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08649_ _04094_ _04102_ _04103_ _00739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_179_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_159_3345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_159_3356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_140_Left_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06419__B _01928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_1090 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_304_clk_I clknet_5_4__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05867__A2 _01634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11660_ net111 net183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_138_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_176_3670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_25_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_25_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10611_ _00355_ clknet_leaf_105_clk rf_ram.memory\[315\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_181_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07069__A1 _03087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_166_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_115_clk clknet_5_15__leaf_clk clknet_leaf_115_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_11591_ _01323_ clknet_leaf_139_clk rf_ram.memory\[264\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_36_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_137_2942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10542_ _00286_ clknet_leaf_143_clk rf_ram.memory\[334\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_146_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06816__A1 _02927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_1114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06933__I _03017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_172_3589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_148_1039 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_319_clk_I clknet_5_5__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_1147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_107_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06292__A2 _01922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10473_ _00217_ clknet_leaf_104_clk rf_ram.memory\[424\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_106_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06029__C1 _01554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09230__A2 _02815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07241__A1 _02795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06044__A2 _01614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11025_ _00762_ clknet_leaf_328_clk rf_ram.memory\[152\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_172_1313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_99_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_185_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05858__A2 _01846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_60_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_106_clk clknet_5_15__leaf_clk clknet_leaf_106_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10809_ _00553_ clknet_leaf_320_clk rf_ram.memory\[552\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_60_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_921 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_144_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06807__A1 _02930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07480__A1 _03356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06283__A2 _01531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06064__B _01526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_97_2193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06000_ rf_ram.memory\[516\]\[1\] _01538_ _01539_ rf_ram.memory\[517\]\[1\] _01540_
+ rf_ram.memory\[519\]\[1\] _02195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XANTENNA__05459__I _01513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput104 net104 o_dbus_dat[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_51_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput115 net115 o_dbus_dat[25] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_10_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput126 net126 o_dbus_dat[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__06035__A2 _01524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput137 net137 o_ext_funct3[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput148 net148 o_ext_rs1[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_58_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput159 net159 o_ext_rs1[29] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_58_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_1112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07783__A2 _03234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_75_1790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07951_ _03654_ _03652_ _03655_ _00489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10119__A1 _05017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_1167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06902_ _02867_ _02939_ _02996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_07882_ _03590_ _03610_ _03612_ _00463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_128_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08732__A1 _04126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06833_ _02930_ _02947_ _02949_ _00077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_37_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09621_ _02828_ _04507_ _04720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09552_ _04478_ net44 _04650_ cpu.immdec.imm19_12_20\[8\] _04672_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_179_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06764_ _02881_ _02899_ _02900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__09288__A2 _04507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08503_ rf_ram.memory\[79\]\[1\] _04006_ _04008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_77_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05715_ _01695_ _01911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__07299__A1 _03225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09483_ cpu.state.cnt_r\[1\] _04620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06695_ rf_ram.memory\[524\]\[1\] _02850_ _02852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_148_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05143__B _01341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08434_ _02971_ _03949_ _03958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_176_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05646_ rf_ram.memory\[498\]\[0\] _01500_ _01763_ rf_ram.memory\[499\]\[0\] _01668_
+ rf_ram.memory\[497\]\[0\] _01842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_58_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08365_ _03884_ _03913_ _03914_ _00644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_46_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05577_ _01695_ _01773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_154_3253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08454__B net126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06259__C1 _01646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07316_ rf_ram.memory\[256\]\[1\] _03258_ _03261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_154_3264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_290_clk_I clknet_5_24__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08296_ rf_ram.memory\[203\]\[1\] _03869_ _03871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_61_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07247_ rf_ram.memory\[420\]\[0\] _03216_ _03217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07471__A1 _02972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_115_2525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_171_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_147_1061 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_115_2536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07178_ _03161_ _03172_ _03174_ _00197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_132_2850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07223__A1 _03190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06129_ rf_ram.memory\[297\]\[1\] _01697_ _02324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA_output155_I net155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08723__A1 _04129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09819_ _04837_ _04854_ _04855_ _01157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06928__I _03013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_243_clk_I clknet_5_21__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_336_clk clknet_5_0__leaf_clk clknet_leaf_336_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_51_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_179_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_1184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_1026 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_174_3618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_174_3629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_876 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11643_ net124 net196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_clkbuf_leaf_258_clk_I clknet_5_17__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_182_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_65_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11574_ _01306_ clknet_leaf_27_clk rf_ram.memory\[191\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_119_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_135_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput17 i_dbus_rdt[23] net17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_123_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput28 i_dbus_rdt[4] net28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput39 i_ibus_rdt[14] net39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10525_ _00269_ clknet_leaf_215_clk rf_ram.memory\[251\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05473__B1 _01519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10456_ _00200_ clknet_leaf_44_clk rf_ram.memory\[198\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_20_421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06017__A2 _01502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_1144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10387_ _00131_ clknet_leaf_272_clk rf_ram.memory\[226\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_53_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08714__A1 _03008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11008_ _00745_ clknet_leaf_1_clk rf_ram.memory\[158\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_53_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_149_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_1240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_177_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_327_clk clknet_5_4__leaf_clk clknet_leaf_327_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__06059__B _01650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05500_ _01695_ _01696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_06480_ rf_ram.memory\[12\]\[1\] _01643_ _01655_ rf_ram.memory\[13\]\[1\] _01653_
+ rf_ram.memory\[15\]\[1\] _02675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_87_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_114_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05431_ rf_ram.memory\[361\]\[0\] _01626_ _01627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_99_2233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_16_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_99_2244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08150_ _03757_ _03778_ _03780_ _00563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05362_ rf_ram.memory\[542\]\[0\] _01532_ _01505_ _01558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_28_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_1000 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_160_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07101_ _03017_ _03126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__06256__A2 _01666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07453__A1 _03326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08081_ rf_ram.memory\[560\]\[1\] _03736_ _03738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_43_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05293_ _01430_ _01487_ _01488_ _01489_ _01490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_126_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05189__I cpu.ctrl.pc vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_67_1066 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07032_ rf_ram.memory\[216\]\[1\] _03079_ _03081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_77_1830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_28_1039 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_183_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_141_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06008__A2 _01501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07205__A1 _02806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_110_2433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08953__A1 _04269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_73_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_110_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08983_ rf_ram.memory\[115\]\[0\] _04310_ _04311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_177_1032 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07934_ _03622_ _03642_ _03644_ _00483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07508__A2 _02889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07865_ _03587_ _03601_ _03602_ _00456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11654__I net104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09604_ _04478_ cpu.immdec.imm30_25\[0\] _04700_ _04712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_155_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06816_ _02927_ _02936_ _02937_ _00072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07796_ _02908_ _03559_ _03560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_27_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05652__I _01617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_108_2395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06747_ _02719_ _02792_ _02887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_09535_ cpu.immdec.imm19_12_20\[2\] _04649_ _04661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_78_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_318_clk clknet_5_5__leaf_clk clknet_leaf_318_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09130__A1 _04401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09466_ _04609_ _01050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06678_ _02836_ _02839_ _02840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_94_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_148_353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06495__A2 _02235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08417_ rf_ram.memory\[29\]\[0\] _03946_ _03947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05629_ rf_ram.memory\[480\]\[0\] _01692_ _01693_ _01825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_114_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09397_ _04571_ _01019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_108_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_1093 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_164_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_74_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05601__B _01707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_1032 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08348_ _03071_ _03903_ _03904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_46_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07444__A1 _02781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_1178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06247__A2 _01719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08279_ rf_ram.memory\[194\]\[0\] _03860_ _03861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_131_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10310_ _00054_ clknet_leaf_272_clk rf_ram.memory\[515\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_132_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_130_2809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11290_ _00005_ clknet_leaf_242_clk cpu.ctrl.pc_plus_4_cy_r vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10241_ _02819_ _05113_ _05114_ _01321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_120_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07747__A2 _03496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08944__A1 _03672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10172_ _02996_ _03134_ _05072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_121_1020 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_160_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_167_3488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06151__C net253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_167_3499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_1150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_1202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_5_9__f_clk_I clknet_3_2_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_1137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_182_clk_I clknet_5_29__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_309_clk clknet_5_5__leaf_clk clknet_leaf_309_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_85_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_62_clk_I clknet_5_8__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_1066 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09121__A1 _04367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_1099 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_197_clk_I clknet_5_28__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07683__A1 _02908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06486__A2 _01613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_1193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_72_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11626_ net76 net148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_13_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_181_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_77_clk_I clknet_5_8__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_182_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_154_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06238__A2 _01510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11557_ _01289_ clknet_leaf_129_clk rf_ram.memory\[44\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_120_clk_I clknet_5_13__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_94_2141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10508_ _00252_ clknet_leaf_219_clk rf_ram.memory\[255\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_94_2152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11488_ _01220_ clknet_leaf_181_clk rf_ram.memory\[274\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09188__A1 _04434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10439_ _00183_ clknet_leaf_222_clk rf_ram.memory\[498\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_55_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_1072 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_135_clk_I clknet_5_24__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06410__A2 _01856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05213__A3 _01385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05980_ rf_ram.memory\[8\]\[0\] _01643_ _01714_ rf_ram.memory\[9\]\[0\] _01653_ rf_ram.memory\[11\]\[0\]
+ _02176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XANTENNA_clkbuf_leaf_15_clk_I clknet_5_2__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_174_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07650_ _03458_ _03466_ _03468_ _00375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06568__I _02751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05472__I _01655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06601_ rf_ram.memory\[234\]\[1\] _02776_ _02778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_88_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07910__A2 _03547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07581_ rf_ram.memory\[356\]\[1\] _03423_ _03426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_149_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09320_ _04528_ _00985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09112__A1 _02959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06532_ _01497_ _01525_ _02718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_88_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_158_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08466__A3 _02709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09251_ _04476_ _04479_ _00965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_168_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07674__A1 _03455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06463_ _01599_ _02645_ _02657_ _01568_ _02658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_34_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_173_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08202_ rf_ram.memory\[537\]\[1\] _03811_ _03813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_28_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05685__B1 _01772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05414_ _01609_ _01610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_09182_ rf_ram.memory\[84\]\[1\] _04432_ _04435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_151_3201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06394_ _01972_ _02587_ _02588_ _02589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_28_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08133_ _03754_ _03769_ _03770_ _00556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_43_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06229__A2 _01801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07426__A1 _03323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05345_ rf_ram.memory\[516\]\[0\] _01538_ _01539_ rf_ram.memory\[517\]\[0\] _01540_
+ rf_ram.memory\[519\]\[0\] _01541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_16_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_114_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08064_ _03721_ _03726_ _03727_ _00530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05276_ _01383_ _01427_ _01449_ _01451_ _01474_ _01475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__05988__A1 _01349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11649__I net99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07015_ rf_ram.memory\[222\]\[1\] _03068_ _03070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_101_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08926__A1 _04266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_1183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_149_3163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05204__A3 _01341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08966_ rf_ram.memory\[118\]\[0\] _04299_ _04300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input31_I i_dbus_rdt[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07917_ _03619_ _03633_ _03634_ _00476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08897_ net243 _03547_ _04257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
Xclkbuf_leaf_95_clk clknet_5_14__leaf_clk clknet_leaf_95_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_127_2760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_162_3396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07848_ _02813_ _03559_ _03592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_162_Right_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_151_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output118_I net118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07779_ rf_ram.memory\[437\]\[0\] _03548_ _03549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_1217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_123_2679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09518_ cpu.immdec.imm19_12_20\[0\] _04646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_151_1057 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10790_ _00534_ clknet_leaf_332_clk rf_ram.memory\[561\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xserv_rf_top_255 o_dbus_adr[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_66_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_140_2993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07665__A1 _03458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06468__A2 _01514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09449_ _04600_ _01042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_13_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_136_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09406__A2 _03991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11411_ _01143_ clknet_leaf_18_clk rf_ram.memory\[187\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_50_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11342_ _01074_ clknet_leaf_216_clk cpu.immdec.imm19_12_20\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_34_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08090__A1 _03721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05979__A1 rf_ram.memory\[10\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_169_3528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_120_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_169_3539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_132_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11273_ _01008_ clknet_leaf_246_clk net208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_186_3842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_186_3853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09029__I _04037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10224_ _03892_ _03134_ _05104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_63_1272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_993 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10155_ rf_ram.memory\[450\]\[1\] _05060_ _05062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_33_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10086_ rf_ram.memory\[30\]\[0\] _05019_ _05020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_86_clk clknet_5_10__leaf_clk clknet_leaf_86_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09342__A1 net213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09342__B2 net224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06156__A1 _01675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_96_1092 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_18_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_18_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09645__A2 _01376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10988_ _00725_ clknet_leaf_27_clk rf_ram.memory\[129\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_128_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_155_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_48_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_169_1318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07656__A1 _03088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06459__A2 _01643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_182_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_170_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_155_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07408__A1 _03289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11609_ net87 net160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_26_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_108_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_10_clk clknet_5_2__leaf_clk clknet_leaf_10_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_05130_ cpu.decode.op21 _01333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_64_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06092__B1 _01721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_1313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06072__B _01615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_70_1708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09581__A1 _03992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08820_ net250 _04195_ _04210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07682__I _03355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08751_ _04129_ _04164_ _04166_ _00778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05963_ rf_ram.memory\[22\]\[0\] _01605_ _01624_ rf_ram.memory\[23\]\[0\] _01617_
+ rf_ram.memory\[21\]\[0\] _02159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_174_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_77_clk clknet_5_8__leaf_clk clknet_leaf_77_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_144_3071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08136__A2 _03009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09333__A1 net240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07702_ _03488_ _03500_ _03501_ _00394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08682_ _02821_ _04078_ _04123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05894_ rf_ram.memory\[94\]\[0\] _01770_ _02090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07633_ _03359_ _03458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_136_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_1127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_1176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_105_2343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_177_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_68_1659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_105_2354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07564_ rf_ram.memory\[318\]\[1\] _03413_ _03415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_85_1973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_85_1984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06515_ cpu.alu.i_rs1 _02699_ _02704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09303_ _03668_ _02909_ _04517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07495_ _03356_ _03371_ _03372_ _00316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_119_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09234_ rf_ram.memory\[329\]\[1\] _04464_ _04467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_29_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_3_Right_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06446_ _02638_ _02640_ _01493_ _02641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_111_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_91_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_160_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_1096 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09165_ rf_ram.memory\[87\]\[1\] _04422_ _04424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06377_ _02568_ _02569_ _02570_ _02571_ _01860_ _02572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_90_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_1250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_983 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_185_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08116_ rf_ram.memory\[553\]\[0\] _03759_ _03760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_146_1148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05328_ _01523_ _01524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_9_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08072__A1 _03724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09096_ _04367_ _04378_ _04380_ _00909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_86_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08047_ _03686_ _03715_ _03716_ _00524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05259_ _01380_ _01382_ _01456_ _01173_ _01458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_TAPCELL_ROW_129_2800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_164_3436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_164_3447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09998_ _04950_ _04964_ _04965_ _01227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_181_3750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_181_3761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08949_ _02983_ _04038_ _04289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_68_clk clknet_5_8__leaf_clk clknet_leaf_68_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_125_2719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06138__A1 _01675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_169_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_4_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_1216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10911_ _00655_ clknet_leaf_39_clk rf_ram.memory\[199\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_54_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10842_ _00586_ clknet_leaf_298_clk rf_ram.memory\[535\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_17_Left_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07638__A1 _03455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_149_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_1069 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10773_ _00517_ clknet_leaf_305_clk rf_ram.memory\[570\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_55_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06157__B _01684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_66_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06310__A1 _01552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_1313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05996__B _01528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_188_3904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06074__B1 _01688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07810__A1 _03557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11325_ _01058_ clknet_leaf_249_clk cpu.state.i_ctrl_misalign vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_26_Left_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_11256_ _00991_ clknet_leaf_77_clk rf_ram.memory\[99\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10207_ rf_ram.memory\[211\]\[1\] _05092_ _05094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_24_1075 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11187_ _00923_ clknet_leaf_57_clk rf_ram.memory\[91\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10138_ rf_ram.memory\[453\]\[0\] _05051_ _05052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_175_1322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_89_2051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_59_clk clknet_5_9__leaf_clk clknet_leaf_59_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10069_ rf_ram.memory\[508\]\[0\] _05008_ _05009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_82_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_187_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_159_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07877__A1 _03590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05337__C1 _01517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_35_Left_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_187_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05888__B1 _02019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09618__A2 _01460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05352__A2 _01532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_175_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06067__B _01599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06300_ rf_ram.memory\[160\]\[1\] _01846_ _01956_ _02495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_63_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_100_2251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_100_2262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_63_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07280_ _02836_ _02992_ _03238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_183_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_1881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06231_ rf_ram.memory\[406\]\[1\] _01623_ _01504_ _02426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_80_1892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_142_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_170_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08054__A1 _03690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06162_ rf_ram.memory\[481\]\[1\] _01697_ _02357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_124_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_44_Left_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06065__B1 _01519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06093_ _02284_ _02285_ _02286_ _02287_ _01658_ _02288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__07801__A1 _02866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05812__B1 _01848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09921_ _04887_ _04915_ _04917_ _01198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_0_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_146_3100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_146_3111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09852_ _01385_ _04487_ _04875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_08803_ net243 _03945_ _04199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09783_ rf_ram.memory\[187\]\[1\] _04831_ _04833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06995_ rf_ram.memory\[226\]\[1\] _03056_ _03058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_77_1238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08109__A2 _03729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08734_ _04129_ _04153_ _04155_ _00772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05946_ rf_ram.memory\[38\]\[0\] _01661_ _01607_ rf_ram.memory\[39\]\[0\] _01609_
+ rf_ram.memory\[37\]\[0\] _02142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_22_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_1_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_53_Left_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07868__A1 _02991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08665_ rf_ram.memory\[158\]\[1\] _04111_ _04113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05877_ _01768_ _02061_ _02072_ _01569_ _02073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_07616_ _03422_ _03446_ _03447_ _00362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_120_2627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_163_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06756__I _02893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08596_ rf_ram.memory\[166\]\[1\] _04068_ _04070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05660__I _01686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_1211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_166_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07547_ rf_ram.memory\[35\]\[0\] _03404_ _03405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_181_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07478_ _02728_ _02815_ _03362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08293__A1 _03230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08971__I _04037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_49_1307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09217_ rf_ram.memory\[67\]\[1\] _04454_ _04456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_162_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06429_ rf_ram.memory\[102\]\[1\] _01641_ _02004_ _02624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_134_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_118_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_62_Left_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08045__A1 _03008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09148_ _04397_ _04412_ _04413_ _00928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_118_2589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_20_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output185_I net185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09793__A1 _04837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09079_ _04364_ _04369_ _04370_ _00902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_47_1075 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11110_ _00846_ clknet_leaf_86_clk rf_ram.memory\[123\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_9_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_1242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11041_ _00778_ clknet_leaf_337_clk rf_ram.memory\[147\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08348__A2 _03903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_71_Left_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_157_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_1063 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09848__A2 _01413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_93_1040 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_1058 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_738 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_184_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10825_ _00569_ clknet_leaf_314_clk rf_ram.memory\[544\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_45_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_156_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_94_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07087__A2 _02911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10756_ _00500_ clknet_leaf_123_clk rf_ram.memory\[478\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_43_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06834__A2 _02941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10687_ _00431_ clknet_leaf_90_clk rf_ram.memory\[415\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_152_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_125_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_180_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_51_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_152_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08587__A2 _03949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09784__A1 _04637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_1115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_1321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06598__A1 _02766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11308_ _01041_ clknet_leaf_265_clk net73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_26_1159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09645__C _01385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11239_ _00975_ clknet_leaf_60_clk rf_ram.memory\[65\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05800_ rf_ram.memory\[168\]\[0\] _01510_ _01527_ _01996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06780_ _02909_ _02911_ _02912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09839__A2 _03984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05731_ rf_ram.memory\[442\]\[0\] _01719_ _01925_ rf_ram.memory\[443\]\[0\] _01926_
+ _01927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_188_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_171_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_65_1607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_102_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08450_ cpu.state.genblk1.misalign_trap_sync_r cpu.state.stage_two_req _03967_ _03968_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_05662_ rf_ram.memory\[473\]\[0\] _01787_ _01858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_72_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06522__B2 _01375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_82_1921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07401_ _03309_ _03083_ _03313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_82_1932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08381_ rf_ram.memory\[180\]\[0\] _03924_ _03925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05593_ rf_ram.memory\[290\]\[0\] _01785_ _01786_ rf_ram.memory\[291\]\[0\] _01788_
+ _01789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_110_1309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_129_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07332_ _03260_ _03268_ _03270_ _00255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_128_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08275__A1 _03852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07263_ _02738_ _02883_ _03227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_116_635 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06214_ rf_ram.memory\[393\]\[1\] _01697_ _02409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_09002_ _02953_ _04303_ _04322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_6_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08027__A1 _03686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07194_ _02813_ _02832_ _03184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_42_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_130_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_115_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06145_ rf_ram.memory\[318\]\[1\] _01804_ _01805_ _02340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__09775__A1 net243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06589__A1 _02748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06076_ rf_ram.memory\[336\]\[1\] _01692_ _01684_ _02271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_112_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11657__I net107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_113_2497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09904_ rf_ram.memory\[345\]\[1\] _04905_ _04907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_6_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_6_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06260__B _01756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10137__A2 _02836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09127__I _02747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07002__A2 _02904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09835_ rf_ram.memory\[61\]\[1\] _04863_ _04865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_77_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09766_ _04822_ _01137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06978_ _03018_ _03044_ _03046_ _00125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06761__A1 _02876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05564__A2 _01662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08717_ rf_ram.memory\[150\]\[1\] _04143_ _04145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_90_1202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05929_ rf_ram.memory\[96\]\[0\] _01922_ _01923_ _02125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09697_ _04740_ net33 _04775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_90_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05604__B _01602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08648_ rf_ram.memory\[161\]\[0\] _04102_ _04103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06513__A1 _01391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_159_3346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_178_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_166_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_176_3660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08579_ _04057_ _04058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_76_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_176_3671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_25_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10610_ _00354_ clknet_leaf_105_clk rf_ram.memory\[315\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_37_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11590_ _01322_ clknet_leaf_303_clk rf_ram.memory\[213\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10073__A1 _03445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_137_2932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_146_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06277__B1 _01953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10541_ _00285_ clknet_leaf_146_clk rf_ram.memory\[372\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_137_2943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_130_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_172_3579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_165_1310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06435__B net251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_40_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10472_ _00216_ clknet_leaf_104_clk rf_ram.memory\[424\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_162_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06029__B1 _01555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_115_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_1040 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07241__A2 _03040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05788__C1 _01702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11024_ _00761_ clknet_leaf_327_clk rf_ram.memory\[152\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08741__A2 _04158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_188_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06752__A1 _02873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_99_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_1000 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_68_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10808_ _00552_ clknet_leaf_321_clk rf_ram.memory\[552\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_60_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_16_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_6_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_103_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_184_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_82_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_1185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10739_ _00483_ clknet_leaf_55_clk rf_ram.memory\[440\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_103_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06345__B _01860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_1248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_97_2194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput105 net105 o_dbus_dat[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_140_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput116 net116 o_dbus_dat[26] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput127 net127 o_dbus_dat[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput138 net138 o_ext_rs1[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_23_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_58_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput149 net149 o_ext_rs1[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_58_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05243__A1 cpu.alu.i_rs1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09509__A1 _04634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_290_clk clknet_5_24__leaf_clk clknet_leaf_290_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_75_1791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07950_ rf_ram.memory\[456\]\[1\] _03652_ _03655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05794__A2 _01989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06901_ _02975_ _02993_ _02995_ _00099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07881_ rf_ram.memory\[446\]\[1\] _03610_ _03612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_128_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09620_ _04643_ _01393_ _04651_ _01094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06832_ rf_ram.memory\[304\]\[1\] _02947_ _02949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09551_ _01391_ cpu.immdec.imm24_20\[0\] _04670_ _04671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06763_ _02898_ _02899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_08502_ _03953_ _04006_ _04007_ _00688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05714_ rf_ram.memory\[436\]\[0\] _01510_ _01910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_37_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09482_ _04619_ _01056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06694_ _02820_ _02850_ _02851_ _00036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_188_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_53_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_148_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08433_ _03956_ _03954_ _03957_ _00669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05645_ rf_ram.memory\[496\]\[0\] _01644_ _01526_ _01841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_188_1310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05703__C1 _01721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_93_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_176_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08248__A1 _03820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_22_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05576_ _01617_ _01772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_135_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_22_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08364_ rf_ram.memory\[184\]\[0\] _03913_ _03914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_163_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06259__B1 _01810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10055__A1 _04982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_154_3254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07315_ _03017_ _03260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_61_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08295_ _03852_ _03869_ _03870_ _00618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_128_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06255__B _01650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07246_ _02882_ _03040_ _03216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07471__A2 _03101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_115_2526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_131_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_115_2537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_132_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07177_ rf_ram.memory\[482\]\[1\] _03172_ _03174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_132_2840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_132_2851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input61_I i_ibus_rdt[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06128_ rf_ram.memory\[296\]\[1\] _01692_ _01693_ _02323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08420__A1 _03922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_281_clk clknet_5_19__leaf_clk clknet_leaf_281_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_06059_ rf_ram.memory\[376\]\[1\] _01649_ _01650_ _02254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_111_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05785__A2 _01799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_888 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09818_ rf_ram.memory\[259\]\[0\] _04854_ _04855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06734__A1 _02795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05537__A2 _01367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09749_ _04804_ net19 _04811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_97_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_178_3700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08487__A1 _03956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06149__C _01658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_166_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_1016 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_174_3619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_1196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_1169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11642_ net123 net195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_65_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05170__B1 _01367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05988__C net254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_181_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11573_ _01305_ clknet_leaf_27_clk rf_ram.memory\[191\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput18 i_dbus_rdt[24] net18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput29 i_dbus_rdt[5] net29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10524_ _00268_ clknet_leaf_215_clk rf_ram.memory\[251\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_91_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_126_1124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10455_ _00199_ clknet_leaf_39_clk rf_ram.memory\[1\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_32_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10386_ _00130_ clknet_leaf_277_clk rf_ram.memory\[226\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_62_1167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_272_clk clknet_5_16__leaf_clk clknet_leaf_272_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_102_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_176_Right_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06973__A1 _03018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08714__A2 _04078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11007_ _00744_ clknet_leaf_295_clk rf_ram.memory\[15\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_176_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_133_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_176_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_90_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_157_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07150__A1 _03126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_185_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05430_ _01514_ _01626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_185_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_145_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05700__A2 _01634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_16_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_99_2234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_157_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10037__A1 _04985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_99_2245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05361_ _01548_ _01549_ _01553_ _01556_ _01494_ _01557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_55_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_5_26__f_clk_I clknet_3_6_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06075__B _01629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07100_ _03123_ _03124_ _03125_ _00168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_114_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08080_ _03721_ _03736_ _03737_ _00536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05292_ cpu.alu.i_rs1 cpu.alu.add_cy_r _01489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07031_ _03050_ _03079_ _03080_ _00144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_114_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_144_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_77_1831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_140_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_23_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08402__A1 _03919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07205__A2 _02941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09450__I0 net75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05216__A1 _01413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_263_clk clknet_5_17__leaf_clk clknet_leaf_263_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_41_1218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_110_2434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_1229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_110_2445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08982_ net242 _04303_ _04310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_11_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_303_clk_I clknet_5_6__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05767__A2 _01846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06964__A1 _03014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_143_Right_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07933_ rf_ram.memory\[440\]\[1\] _03642_ _03644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_177_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07864_ rf_ram.memory\[42\]\[0\] _03601_ _03602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06716__A1 _02826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09603_ _04643_ _04709_ _04710_ _04711_ _01085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_78_1174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06815_ rf_ram.memory\[288\]\[0\] _02936_ _02937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_318_clk_I clknet_5_5__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07795_ _03088_ _03559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_97_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_27_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09534_ _04526_ net38 _04660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_108_2396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08469__A1 _02714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06746_ _02876_ _02884_ _02886_ _00053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_148_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09465_ net82 net83 _04604_ _04609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_38_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06677_ _02838_ _02839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__07141__A1 _02795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08416_ _02959_ _03945_ _03946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_171_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_164_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_149_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05628_ _01821_ _01823_ _01746_ _01824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_09396_ net220 _04561_ _04564_ net221 _04571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_148_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_149_1102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09969__A1 _03672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08347_ _03902_ _03903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_11_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05559_ _01613_ _01755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_117_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07444__A2 _02815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08641__A1 _04097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08278_ _03230_ _02894_ _03860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_15_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_1107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_1313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_144_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07229_ rf_ram.memory\[424\]\[1\] _03204_ _03206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_15_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_104_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10240_ rf_ram.memory\[213\]\[0\] _05113_ _05114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_254_clk clknet_5_20__leaf_clk clknet_leaf_254_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08944__A2 _02899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10171_ _05049_ _05069_ _05071_ _01294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05758__A2 _01614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06955__A1 _03018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_167_3489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_110_Right_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_35_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06707__A1 _02752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_187_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07380__A1 _02775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06183__A2 _01785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11135__CLK clknet_5_10__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05930__A2 _01785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05999__B _01506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_182_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07683__A2 _03390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_154_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11625_ net75 net147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_13_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11556_ _01288_ clknet_leaf_112_clk rf_ram.memory\[450\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08632__A1 _04058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_94_2142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10507_ _00251_ clknet_leaf_190_clk rf_ram.memory\[272\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_94_2153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11487_ _01219_ clknet_leaf_183_clk rf_ram.memory\[274\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05997__A2 _01532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10438_ _00182_ clknet_leaf_222_clk rf_ram.memory\[498\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_110_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07199__A1 _02761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_55_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_245_clk clknet_5_21__leaf_clk clknet_leaf_245_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10369_ _00113_ clknet_leaf_38_clk rf_ram.memory\[206\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05749__A2 _01942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06946__A1 _02728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_100_1149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08699__A1 _02828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06600_ _02743_ _02776_ _02777_ _00016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_178_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07580_ _03359_ _03425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__10258__A1 _02825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09112__A2 _04005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06531_ _01498_ _01503_ _02717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__07123__A1 _03123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05702__B _01615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09250_ _04478_ cpu.bufreg.i_sh_signed _04479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_173_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06462_ _02648_ _02651_ _01599_ _02656_ _02657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__08871__A1 _04237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_185_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_875 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08201_ _03787_ _03811_ _03812_ _00582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_56_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05413_ _01513_ _01609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_06393_ rf_ram.memory\[70\]\[1\] _01719_ _01925_ rf_ram.memory\[71\]\[1\] _01912_
+ rf_ram.memory\[69\]\[1\] _02588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_09181_ _04400_ _04434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_151_3202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_141_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05344_ _01520_ _01540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_08132_ rf_ram.memory\[550\]\[0\] _03769_ _03770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_161_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_32_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08063_ rf_ram.memory\[563\]\[0\] _03726_ _03727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05275_ _01458_ _01468_ _01473_ _01474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_141_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_144_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07014_ _03050_ _03068_ _03069_ _00138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_144_1054 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_1174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_144_1076 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_242_clk_I clknet_5_21__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_236_clk clknet_5_22__leaf_clk clknet_leaf_236_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_149_3164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08965_ _03008_ _04038_ _04299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11665__I net116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07916_ rf_ram.memory\[45\]\[0\] _03633_ _03634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08896_ _04237_ _04254_ _04256_ _00833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_leaf_257_clk_I clknet_5_20__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input24_I i_dbus_rdt[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_127_2750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_127_2761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07847_ _03590_ _03588_ _03591_ _00449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_162_3397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06165__A2 _01735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07362__A1 _03260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_1101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07778_ _03547_ _03072_ _03548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05912__A2 _01856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10249__A1 _02838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09517_ _04643_ _04644_ _04645_ _01065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_94_701 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06729_ rf_ram.memory\[518\]\[0\] _02874_ _02875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07114__A1 _02716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xserv_rf_top_256 o_dbus_adr[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_151_1069 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_140_2994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09448_ net74 net75 _04593_ _04600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_82_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_109_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09379_ net211 _04561_ _04552_ net212 _04562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_46_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11410_ _01142_ clknet_leaf_20_clk rf_ram.memory\[77\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_124_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_164_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_152_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08614__A1 _04062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11341_ _01073_ clknet_leaf_216_clk cpu.immdec.imm19_12_20\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_62_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05979__A2 _01686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06443__B _01601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_169_3529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11272_ _01007_ clknet_leaf_246_clk net207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_186_3843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_227_clk clknet_5_23__leaf_clk clknet_leaf_227_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_123_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_186_3854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10223_ _05081_ _05101_ _05103_ _01314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_24_1235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_33_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10154_ _05046_ _05060_ _05061_ _01287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_33_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10085_ _02916_ _03035_ _05019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05573__I _01650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09342__A2 _03991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07353__A1 _03055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_1212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05903__A2 _01652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_173_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_1320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_18_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_187_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10987_ _00724_ clknet_leaf_330_clk rf_ram.memory\[164\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_85_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07656__A2 _03135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06313__C1 _01679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_139_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_154_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11608_ cpu.state.i_ctrl_misalign net149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_170_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08605__A1 _04058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_984 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11539_ _01271_ clknet_leaf_117_clk rf_ram.memory\[392\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_13_528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_180_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_218_clk clknet_5_22__leaf_clk clknet_leaf_218_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_0_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09030__A1 net247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_70_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07592__A1 _03425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08750_ rf_ram.memory\[147\]\[1\] _04164_ _04166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06579__I _02760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05962_ rf_ram.memory\[20\]\[0\] _01536_ _02158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_40_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05483__I _01624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07701_ rf_ram.memory\[400\]\[0\] _03500_ _03501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_144_3061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_144_3072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09333__A2 _04037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_1167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08681_ _04097_ _04120_ _04122_ _00752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_79_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06147__A2 _01808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05893_ _02077_ _02081_ _02085_ _02088_ _02089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_178_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07632_ _03455_ _03456_ _03457_ _00368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_105_2344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_178_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_75_1188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_105_2355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07563_ _03389_ _03413_ _03414_ _00342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_88_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09097__A1 net237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_948 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_85_1974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_85_1985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09302_ _04466_ _04514_ _04516_ _00979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06514_ _01388_ _02702_ _01399_ _01421_ _02703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_07494_ rf_ram.memory\[364\]\[0\] _03371_ _03372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_36_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_1240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08844__A1 _04205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_146_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_1104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09233_ _04400_ _04466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_06445_ rf_ram.memory\[34\]\[1\] _01605_ _01607_ rf_ram.memory\[35\]\[1\] _02639_
+ _02640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_119_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09839__B _02709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_173_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_72_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09164_ _04397_ _04422_ _04423_ _00934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06376_ rf_ram.memory\[248\]\[1\] _01863_ _01793_ rf_ram.memory\[249\]\[1\] _01696_
+ rf_ram.memory\[251\]\[1\] _02571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_32_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08115_ _02751_ _03729_ _03759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05327_ _01509_ _01523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_71_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_995 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09095_ rf_ram.memory\[97\]\[1\] _04378_ _04380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_31_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_181_clk_I clknet_5_29__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08046_ rf_ram.memory\[566\]\[0\] _03715_ _03716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05258_ _01442_ _01457_ _01453_ _01455_ _01173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_3_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_209_clk clknet_5_25__leaf_clk clknet_leaf_209_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA_clkbuf_leaf_61_clk_I clknet_5_9__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05189_ cpu.ctrl.pc _01389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_101_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_129_2801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_164_3437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_164_3448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_196_clk_I clknet_5_25__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09997_ rf_ram.memory\[276\]\[0\] _04964_ _04965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07583__A1 _02935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06386__A2 _01808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_181_3751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08948_ _04269_ _04286_ _04288_ _00853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_181_3762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_76_clk_I clknet_5_10__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output130_I net130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_4_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08879_ _04234_ _04245_ _04246_ _00826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_4_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07335__A1 _03257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10910_ _00654_ clknet_leaf_39_clk rf_ram.memory\[199\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_98_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_1239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10841_ _00585_ clknet_leaf_311_clk rf_ram.memory\[536\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_67_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_184_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10772_ _00516_ clknet_leaf_305_clk rf_ram.memory\[570\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08835__A1 _03672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05649__A1 _01600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_134_clk_I clknet_5_24__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_14_clk_I clknet_5_2__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_1037 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_188_3905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_149_clk_I clknet_5_26__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11324_ _01057_ clknet_leaf_249_clk net138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_50_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_160_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_120_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_29_clk_I clknet_5_1__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05821__A1 net251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11255_ _00003_ clknet_leaf_218_clk cpu.alu.add_cy_r vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09012__A1 _02774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10206_ _05078_ _05092_ _05093_ _01307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_11186_ _00922_ clknet_leaf_57_clk rf_ram.memory\[91\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_98_1133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_101_1244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10137_ _02794_ _02836_ _05051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_89_2052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_13_Right_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10068_ _02838_ _03158_ _05008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06129__A2 _01697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05337__B1 _01521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09079__A1 _04364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06348__B _01650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_159_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_169_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_100_2252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_63_1568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_63_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_100_2263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06301__A2 _01664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06230_ _02423_ _02424_ _01629_ _02425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_72_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_1882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_170_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_1893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_171_945 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_22_Right_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_110_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06161_ rf_ram.memory\[480\]\[1\] _01692_ _01693_ _02356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05478__I _01349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06092_ rf_ram.memory\[328\]\[1\] _01724_ _01721_ rf_ram.memory\[329\]\[1\] _01713_
+ rf_ram.memory\[331\]\[1\] _02287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_111_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07801__A2 _03234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_1171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_123_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09920_ rf_ram.memory\[343\]\[1\] _04915_ _04917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_40_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_1121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_146_3101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_146_3112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09851_ _02713_ _04487_ _04874_ _01170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_0_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09554__A2 _01491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07565__A1 _03393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06368__A2 _01989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08802_ _04170_ _04196_ _04198_ _00797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09782_ _04634_ _04831_ _04832_ _01143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06994_ _03050_ _03056_ _03057_ _00130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_31_Right_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08733_ rf_ram.memory\[148\]\[1\] _04153_ _04155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05945_ rf_ram.memory\[36\]\[0\] _01536_ _02141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07317__A1 _03260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_0_Left_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_1_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08664_ _04094_ _04111_ _04112_ _00745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_96_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07868__A2 _03559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05876_ _01600_ _02066_ _02071_ _02072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_15_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_178_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07615_ rf_ram.memory\[313\]\[0\] _03446_ _03447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_178_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_120_2617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08595_ _04058_ _04068_ _04069_ _00719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_120_2628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06258__B _01805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07546_ _02921_ _02889_ _03404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08817__A1 _04202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_165_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07477_ _03360_ _03357_ _03361_ _00309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09569__B _04678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_1070 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08293__A2 _02781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_666 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_40_Right_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_118_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_134_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09216_ _04431_ _04454_ _04455_ _00954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_107_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06428_ _02619_ _02620_ _02621_ _02622_ _01860_ _02623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_173_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_161_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_162_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_995 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09147_ rf_ram.memory\[8\]\[0\] _04412_ _04413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08045__A2 _03693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06359_ _02551_ _02553_ _01564_ _02554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_20_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_86_1070 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09078_ rf_ram.memory\[57\]\[0\] _04369_ _04370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_output178_I net178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_188_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08029_ _03690_ _03703_ _03705_ _00517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_97_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11040_ _00777_ clknet_leaf_0_clk rf_ram.memory\[147\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07556__A1 _02806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_1318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_188_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07308__A1 _03222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_1167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06531__A2 _01503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10824_ _00568_ clknet_leaf_314_clk rf_ram.memory\[544\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_170_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_138_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_45_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_165_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10755_ _00499_ clknet_leaf_203_clk rf_ram.memory\[46\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_165_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05800__B _01527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_137_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10686_ _00430_ clknet_leaf_90_clk rf_ram.memory\[415\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_129_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05298__I _01493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_180_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06598__A2 _02775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_10_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11307_ _01040_ clknet_leaf_265_clk net72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_50_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_65_1198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11238_ _00974_ clknet_leaf_61_clk rf_ram.memory\[65\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06350__C _01717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_5_27__f_clk clknet_3_6_0_clk clknet_5_27__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_11169_ _00905_ clknet_leaf_62_clk rf_ram.memory\[98\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_101_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07018__I _03071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_141_3020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_1115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05730_ rf_ram.memory\[441\]\[0\] _01918_ _01926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_175_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_1261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_1148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_158_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_65_1608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05661_ _01695_ _01857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_187_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_188_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06522__A2 _01376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_82_1922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07400_ _03292_ _03310_ _03312_ _00281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_129_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08380_ _03134_ _03903_ _03924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05592_ rf_ram.memory\[289\]\[0\] _01787_ _01788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_07331_ rf_ram.memory\[271\]\[1\] _03268_ _03270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_1170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_171_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07262_ _03225_ _03223_ _03226_ _00229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_183_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09001_ _04301_ _04319_ _04321_ _00873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_26_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06213_ rf_ram.memory\[392\]\[1\] _01692_ _01693_ _02408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_170_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09224__A1 _03319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07193_ _03161_ _03181_ _03183_ _00203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_60_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_182_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06144_ _02335_ _02336_ _02337_ _02338_ _01717_ _02339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__09775__A2 _04507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_987 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_112_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06075_ _02267_ _02269_ _01629_ _02270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_111_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_113_2498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09903_ _04884_ _04905_ _04906_ _01191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_6_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07538__A1 _03389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09834_ _04837_ _04863_ _04864_ _01163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05549__B1 _01696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09765_ net121 _04766_ _04760_ net122 _04821_ _04822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_06977_ rf_ram.memory\[427\]\[1\] _03044_ _03046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_77_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08468__B _03984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08716_ _04126_ _04143_ _04144_ _00765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_69_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05928_ rf_ram.memory\[100\]\[0\] _01863_ _01848_ rf_ram.memory\[101\]\[0\] _01696_
+ rf_ram.memory\[103\]\[0\] _02124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_09696_ _04774_ _01115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_68_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08647_ net238 _04067_ _04102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05859_ rf_ram.memory\[225\]\[0\] _01664_ _02055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_95_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07710__A1 net240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_159_3347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_1070 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08578_ _02742_ _04057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_176_3661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_25_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07529_ rf_ram.memory\[361\]\[1\] _03391_ _03394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_147_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_187_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_147_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_135_923 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_1132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10540_ _00284_ clknet_leaf_147_clk rf_ram.memory\[372\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10073__A2 _03134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_137_2933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_137_2944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_1322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_40_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10471_ _00215_ clknet_leaf_100_clk rf_ram.memory\[425\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_40_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_157_Right_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_103_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05788__B1 _01608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11023_ _00760_ clknet_leaf_41_clk rf_ram.memory\[39\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_86_2000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06677__I _02838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05581__I _01686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_188_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_87_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_87_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_184_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_170_1072 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_135_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_68_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_670 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10807_ _00551_ clknet_leaf_322_clk rf_ram.memory\[553\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_27_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_60_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10738_ _00482_ clknet_leaf_55_clk rf_ram.memory\[440\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_137_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_55_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09206__A1 _04431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_989 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10669_ _00413_ clknet_leaf_108_clk rf_ram.memory\[377\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_124_Right_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_88_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_97_2195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput106 net106 o_dbus_dat[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_11_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput117 net117 o_dbus_dat[27] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_105_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput128 net128 o_dbus_dat[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput139 net139 o_ext_rs1[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_58_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_142_1174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_75_1792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06900_ rf_ram.memory\[280\]\[1\] _02993_ _02995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07880_ _03587_ _03610_ _03611_ _00462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08193__A1 _03790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09390__B1 _04564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06831_ _02927_ _02947_ _02948_ _00076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07940__A1 _02781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09550_ _01391_ _04644_ _04669_ _04670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__05705__B _01504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06762_ _02750_ _02887_ _02898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__05491__I _01686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08501_ rf_ram.memory\[79\]\[0\] _04006_ _04007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05713_ _01756_ _01909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_37_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09481_ net89 _04618_ _01411_ _04619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_76_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06693_ rf_ram.memory\[524\]\[0\] _02850_ _02851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_176_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08432_ rf_ram.memory\[59\]\[1\] _03954_ _03957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_90_Left_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05644_ rf_ram.memory\[500\]\[0\] _01509_ _01668_ rf_ram.memory\[501\]\[0\] _01519_
+ rf_ram.memory\[503\]\[0\] _01840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XANTENNA__05703__B1 _01726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_176_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_188_1322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08363_ _02991_ _03903_ _03913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_110_1107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05575_ rf_ram.memory\[302\]\[0\] _01770_ _01771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_129_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_22_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07314_ _03257_ _03258_ _03259_ _00248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_128_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_34_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_1237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_154_3255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08294_ rf_ram.memory\[203\]\[0\] _03869_ _03870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_117_945 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09996__A2 _03135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07245_ _03193_ _03213_ _03215_ _00223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09847__B _01391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_115_2527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_115_2538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_132_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07176_ _03157_ _03172_ _03173_ _00196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_41_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07759__A1 _03521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_132_2841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11668__I net119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_132_2852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06127_ _01769_ _02320_ _02321_ _02322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_169_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06271__B _01956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input54_I i_ibus_rdt[29] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05234__A2 _01418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06058_ _01527_ _02251_ _02252_ _02253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_10_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08184__A1 _02838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_5_10__f_clk clknet_3_2_0_clk clknet_5_10__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09817_ net240 _03253_ _04854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06734__A2 _02846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_1132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09748_ _04810_ _01131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_154_1034 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_178_3701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_946 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09679_ net1 net28 _04736_ net124 _04761_ _04762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__06498__A1 _02690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_1066 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_1028 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_1077 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_670 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_90_1099 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11641_ net120 net192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__05170__A1 _01353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06446__B _01493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11572_ _01304_ clknet_leaf_30_clk rf_ram.memory\[210\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_65_876 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_135_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07998__A1 _03654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput19 i_dbus_rdt[25] net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10523_ _00267_ clknet_leaf_194_clk rf_ram.memory\[268\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_108_989 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_load_slew244_I _02821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_740 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05473__A2 _01500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10454_ _00198_ clknet_leaf_41_clk rf_ram.memory\[1\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_161_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_946 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_131_970 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10385_ _00129_ clknet_leaf_277_clk rf_ram.memory\[227\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05576__I _01617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_1266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_62_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06422__A1 _01909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08175__A1 _03787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11006_ _00743_ clknet_leaf_295_clk rf_ram.memory\[15\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_53_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07922__A1 _03619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_158_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06489__A1 _01348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06356__B _01551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_99_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_16_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05360_ rf_ram.memory\[530\]\[0\] _01501_ _01554_ rf_ram.memory\[531\]\[0\] _01555_
+ rf_ram.memory\[529\]\[0\] _01556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XTAP_TAPCELL_ROW_99_2246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07989__A1 _03672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05291_ _01486_ _01434_ _01438_ _01488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_67_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_915 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_113_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07030_ rf_ram.memory\[216\]\[0\] _03079_ _03080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_125_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06870__I _02825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_77_1832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_140_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06091__B _01602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09450__I1 net76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05486__I _01508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_110_2435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08981_ _04301_ _04307_ _04309_ _00865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_11_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_110_2446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07932_ _03619_ _03642_ _03643_ _00482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08797__I _04077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_1131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07863_ _02774_ _02869_ _03601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_120_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_1310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06814_ _02935_ _02904_ _02936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_39_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09602_ cpu.immdec.imm24_20\[3\] _04703_ _04526_ _04711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07794_ _03557_ _03555_ _03558_ _00429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_97_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_119_Left_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_27_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09533_ _04478_ cpu.immdec.imm19_12_20\[3\] _04659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06745_ rf_ram.memory\[516\]\[1\] _02884_ _02886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_108_2397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09666__A1 net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09464_ _04608_ _01049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_38_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06676_ _02716_ _02837_ _02838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_94_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07141__A2 _02911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08415_ _02996_ _03945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_93_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05627_ rf_ram.memory\[490\]\[0\] _01687_ _01688_ rf_ram.memory\[491\]\[0\] _01822_
+ _01823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_09395_ _04570_ _01018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_11_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1050 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1061 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_1114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08346_ _02731_ _02797_ _03902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_15_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05558_ _01527_ _01752_ _01753_ _01754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__09969__A2 _02946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_1094 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_172_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09577__B cpu.decode.opcode\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08277_ _03855_ _03857_ _03859_ _00611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05489_ rf_ram.memory\[344\]\[0\] _01683_ _01684_ _01685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_104_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_1089 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_128_Left_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_144_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07228_ _03190_ _03204_ _03205_ _00216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05455__A2 _01649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06652__A1 _02748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07159_ _02915_ _02946_ _03163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05207__A2 _01382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10170_ rf_ram.memory\[447\]\[1\] _05069_ _05071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_output160_I net160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_35_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_35_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_137_Left_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06707__A2 _02846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07904__A1 _03622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07380__A2 _03253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_1139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09657__A1 net98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_85_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_97_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05679__C1 _01810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_69_Right_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09409__A1 _01436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_190_clk clknet_5_28__leaf_clk clknet_leaf_190_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_154_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_154_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11624_ net74 net146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_33_1281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_13_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_146_Left_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_108_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_170_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11555_ _01287_ clknet_leaf_113_clk rf_ram.memory\[450\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_52_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_108_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05446__A2 _01641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10506_ _00250_ clknet_leaf_189_clk rf_ram.memory\[272\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_94_2143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11486_ _01218_ clknet_leaf_134_clk rf_ram.memory\[464\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_94_2154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10437_ _00181_ clknet_leaf_223_clk rf_ram.memory\[486\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_122_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_150_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_55_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07199__A2 _02941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_55_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_78_Right_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_0_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10368_ _00112_ clknet_leaf_38_clk rf_ram.memory\[206\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06946__A2 _02766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_1740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_178_1321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10299_ _00043_ clknet_leaf_316_clk rf_ram.memory\[521\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_155_Left_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08148__A1 _03754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06159__B1 _01688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08699__A2 _02921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09896__A1 _02828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09442__S _04593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_1073 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09648__A1 net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_87_Right_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_137_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06530_ _01512_ _01497_ _02716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_158_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_146_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06461_ _02652_ _02653_ _02654_ _02655_ rf_ram.i_raddr\[3\] _02656_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_158_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06086__B _01602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_181_clk clknet_5_29__leaf_clk clknet_leaf_181_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_EDGE_ROW_164_Left_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_157_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08200_ rf_ram.memory\[537\]\[0\] _03811_ _03812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_173_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_56_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05412_ _01607_ _01608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__05685__A2 _01711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09180_ _04431_ _04432_ _04433_ _00940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06882__A1 _02975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06392_ rf_ram.memory\[68\]\[1\] _01510_ _02587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_111_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_151_3203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08131_ _02805_ _03765_ _03769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_28_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05343_ _01516_ _01539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_71_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_172_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_16_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06634__A1 _02748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08062_ net242 _03693_ _03726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_05274_ _01381_ _01469_ _01472_ _01473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_114_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07013_ rf_ram.memory\[222\]\[0\] _03068_ _03069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_96_Right_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_113_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_114_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05842__C1 _01645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08387__A1 _03919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_110_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10194__A1 _03892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_149_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_173_Left_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_149_3165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08964_ _04057_ _04298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_45_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07915_ _02844_ _02869_ _03633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08895_ rf_ram.memory\[127\]\[1\] _04254_ _04256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07846_ rf_ram.memory\[431\]\[1\] _03588_ _03591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09860__B _02714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_127_2751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_127_2762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_162_3398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_169_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input17_I i_dbus_rdt[23] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07777_ _03039_ _03547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__09639__A1 _02971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_1135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_149_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06728_ _02806_ _02846_ _02874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09516_ _04524_ net57 _04645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10249__A2 _03035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_1292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_1172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xserv_rf_top_257 o_mdu_valid vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XPHY_EDGE_ROW_182_Left_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_140_2995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09447_ _04599_ _01041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_66_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06659_ _02820_ _02823_ _02824_ _00028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_94_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_172_clk clknet_5_30__leaf_clk clknet_leaf_172_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_136_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05676__A2 _01804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06873__A1 _02813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09378_ _03990_ _04561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_164_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_152_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08329_ _03887_ _03889_ _03891_ _00631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09811__A1 _04840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11340_ _01072_ clknet_leaf_215_clk cpu.immdec.imm19_12_20\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_90_985 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_166_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_1253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11271_ _01006_ clknet_leaf_247_clk net206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_105_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_1230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_186_3844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10222_ rf_ram.memory\[23\]\[1\] _05101_ _05103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_186_3855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10185__A1 _05078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_5_8__f_clk clknet_3_2_0_clk clknet_5_8__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__07050__A1 _02806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10153_ rf_ram.memory\[450\]\[0\] _05060_ _05061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_33_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10084_ _05017_ _05015_ _05018_ _01260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_50_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09878__A1 _04884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1023 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07353__A2 _02839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08550__A1 _04023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_173_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_57_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_18_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05803__B _01564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_186_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10986_ _00723_ clknet_leaf_331_clk rf_ram.memory\[164\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_168_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08302__A1 _03855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_163_clk clknet_5_30__leaf_clk clknet_leaf_163_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__05522__C _01717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06313__B1 _01793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_48_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_302_clk_I clknet_5_6__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_155_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_65_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11607_ cpu.csr_d_sel net137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_65_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_154_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_142_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_25_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09802__A1 net246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11538_ _01270_ clknet_leaf_110_clk rf_ram.memory\[312\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_317_clk_I clknet_5_5__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05824__C1 _01968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06092__A2 _01724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11469_ _01201_ clknet_leaf_170_clk rf_ram.memory\[341\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_151_884 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_96_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_110_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_21_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10176__A1 _05049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09030__A2 _04339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_0_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_188_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_input9_I i_dbus_rdt[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05961_ _01599_ _02144_ _02156_ _01568_ _02157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_40_1071 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09869__A1 _04884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_1124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07700_ _02945_ _03481_ _03500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_139_1135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_144_3062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_1270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_144_3073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08680_ rf_ram.memory\[559\]\[1\] _04120_ _04122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_75_1112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05892_ _01972_ _02086_ _02087_ _02088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__08541__A1 net246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_178_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07631_ rf_ram.memory\[388\]\[0\] _03456_ _03457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_152_1313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_105_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_105_2356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07562_ rf_ram.memory\[318\]\[0\] _03413_ _03414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09097__A2 _04339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_85_1975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09301_ rf_ram.memory\[66\]\[1\] _04514_ _04516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_122_2670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06513_ _01391_ _02701_ _02702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_75_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_85_1986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_154_clk clknet_5_26__leaf_clk clknet_leaf_154_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07493_ _02788_ _03101_ _03371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10100__A1 _02800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_146_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09232_ _04463_ _04464_ _04465_ _00960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_150_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_1032 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06444_ rf_ram.memory\[33\]\[1\] _01513_ _02639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_57_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_91_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_185_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_90_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09163_ rf_ram.memory\[87\]\[0\] _04422_ _04423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_145_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06375_ rf_ram.memory\[250\]\[1\] _01989_ _01783_ _02570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_clkbuf_5_10__f_clk_I clknet_3_2_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08114_ _03757_ _03755_ _03758_ _00549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_12_1195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05326_ rf_ram.memory\[524\]\[0\] _01511_ _01517_ rf_ram.memory\[525\]\[0\] _01521_
+ rf_ram.memory\[527\]\[0\] _01522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_31_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09094_ _04364_ _04378_ _04379_ _00908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_126_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_86_1274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05815__C1 _01786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08045_ _03008_ _03693_ _03715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07280__A1 _02836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05257_ cpu.mem_if.signbit _01457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_102_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05830__A2 _01537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10167__A1 _02908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05188_ _01384_ _01387_ _01388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_177_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_164_3438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09996_ _02940_ _03135_ _04964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_164_3449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07583__A2 _02839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_181_3752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08947_ rf_ram.memory\[449\]\[1\] _04286_ _04288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05607__C _01717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_181_3763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08878_ rf_ram.memory\[128\]\[0\] _04245_ _04246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_4_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07829_ rf_ram.memory\[412\]\[1\] _03578_ _03580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_93_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10840_ _00584_ clknet_leaf_312_clk rf_ram.memory\[536\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_67_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05897__A2 _01683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_183_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10771_ _00515_ clknet_leaf_305_clk rf_ram.memory\[571\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_145_clk clknet_5_26__leaf_clk clknet_leaf_145_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_67_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08835__A2 _03072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_136_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06454__B _01601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_43_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_188_3906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_151_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11323_ _01056_ clknet_leaf_254_clk net89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__06074__A2 _01623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07271__A1 _03222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11254_ _00990_ clknet_leaf_150_clk rf_ram.memory\[309\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_31_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_127_1094 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09484__C _03989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09012__A2 _03945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_1191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10205_ rf_ram.memory\[211\]\[0\] _05092_ _05093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07023__A1 _03053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11185_ _00921_ clknet_leaf_56_clk rf_ram.memory\[92\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08771__A1 _04170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10136_ _05049_ _05047_ _05050_ _01280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_59_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_89_2053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_1278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10067_ _04985_ _05005_ _05007_ _01254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08523__A1 _03956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05888__A2 _01804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_67_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_241_clk_I clknet_5_21__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_136_clk clknet_5_26__leaf_clk clknet_leaf_136_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_35_1173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10969_ _00706_ clknet_leaf_188_clk rf_ram.memory\[489\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_35_1184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06298__C1 _01516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_100_2253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_63_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_100_2264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09659__C _04740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_1894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_256_clk_I clknet_5_20__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06160_ _02352_ _02354_ _01746_ _02355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_108_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07262__A1 _03225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06065__A2 _01500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06091_ rf_ram.memory\[330\]\[1\] _01706_ _01602_ _02286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05812__A2 _01711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10149__A1 _05046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_146_3102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07014__A1 _03050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05708__B _01903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_146_3113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09850_ cpu.state.cnt_r\[3\] cpu.state.o_cnt\[2\] _04874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08762__A1 _02760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06222__C1 _01793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08801_ rf_ram.memory\[140\]\[1\] _04196_ _04198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06993_ rf_ram.memory\[226\]\[0\] _03056_ _03057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09781_ rf_ram.memory\[187\]\[0\] _04831_ _04832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_77_1218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08732_ _04126_ _04153_ _04154_ _00771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05944_ _02137_ _02139_ _01493_ _02140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08514__A1 _02787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_1_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08663_ rf_ram.memory\[158\]\[0\] _04111_ _04112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05875_ _02067_ _02068_ _02069_ _02070_ _01860_ _02071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_96_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07614_ _03445_ _02984_ _03446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__05879__A2 _01531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08594_ rf_ram.memory\[166\]\[0\] _04068_ _04069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_120_2618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_209_clk_I clknet_5_25__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_120_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_166_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07545_ _03393_ _03401_ _03403_ _00335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_138_Right_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_53_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_127_clk clknet_5_13__leaf_clk clknet_leaf_127_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_49_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_158_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07476_ rf_ram.memory\[366\]\[1\] _03357_ _03361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_146_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09215_ rf_ram.memory\[67\]\[0\] _04454_ _04455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06427_ rf_ram.memory\[104\]\[1\] _01677_ _01793_ rf_ram.memory\[105\]\[1\] _01679_
+ rf_ram.memory\[107\]\[1\] _02622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_146_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06274__B _01564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09146_ net250 _03035_ _04412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_161_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06358_ rf_ram.memory\[234\]\[1\] _01940_ _01959_ rf_ram.memory\[235\]\[1\] _02552_
+ _02553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_60_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_20_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06056__A2 _01641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05309_ _01504_ _01505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__07253__A1 _03190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09077_ _03668_ _02984_ _04369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_06289_ rf_ram.memory\[142\]\[1\] _01770_ _02484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_114_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08028_ rf_ram.memory\[570\]\[1\] _03703_ _03705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_102_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_163_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_141_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_9_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07556__A2 _03390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08753__A1 net236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09979_ rf_ram.memory\[274\]\[1\] _04951_ _04954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_157_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08505__A1 _01369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_110_Left_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_170_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_1146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_1179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_1059 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10823_ _00567_ clknet_leaf_321_clk rf_ram.memory\[545\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_118_clk clknet_5_12__leaf_clk clknet_leaf_118_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_EDGE_ROW_105_Right_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_45_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10754_ _00498_ clknet_leaf_132_clk rf_ram.memory\[46\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_138_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_598 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_94_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_165_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07492__A1 _03360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_125_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10685_ _00429_ clknet_leaf_80_clk rf_ram.memory\[436\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_109_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_82_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_1111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_670 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08992__A1 net248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11306_ _01039_ clknet_leaf_265_clk net71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__06452__C1 _01635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_1188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11237_ _00973_ clknet_leaf_257_clk cpu.genblk3.csr.mcause3_0\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_121_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08744__A1 _04157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11168_ _00904_ clknet_leaf_77_clk rf_ram.memory\[98\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05558__A1 _01527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10119_ _05017_ _05037_ _05039_ _01274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_11099_ _00835_ clknet_leaf_99_clk rf_ram.memory\[429\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_141_3010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_141_3021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09514__I _03992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_171_1018 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_1104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06359__B _01564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_1235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_117_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_leaf_180_clk_I clknet_5_31__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_65_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05660_ _01686_ _01856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__09450__S _04593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_82_1923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_109_clk clknet_5_15__leaf_clk clknet_leaf_109_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_58_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05591_ _01514_ _01787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA_clkbuf_leaf_60_clk_I clknet_5_9__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07330_ _03257_ _03268_ _03269_ _00254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_175_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_45_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07483__A1 _02844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07261_ rf_ram.memory\[418\]\[1\] _03223_ _03226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06286__A2 _01915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_195_clk_I clknet_5_25__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05710__C _01670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09000_ rf_ram.memory\[112\]\[1\] _04319_ _04321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_115_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05494__B1 _01688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06212_ _01769_ _02405_ _02406_ _02407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
Xclkbuf_3_7_0_clk clknet_0_clk clknet_3_7_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA_clkbuf_leaf_75_clk_I clknet_5_10__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07192_ rf_ram.memory\[473\]\[1\] _03181_ _03183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09224__A2 _02866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07235__A1 _03193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06143_ rf_ram.memory\[306\]\[1\] _01652_ _01726_ rf_ram.memory\[307\]\[1\] _01721_
+ rf_ram.memory\[305\]\[1\] _02338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_143_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_1255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_1266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06074_ rf_ram.memory\[346\]\[1\] _01623_ _01688_ rf_ram.memory\[347\]\[1\] _02268_
+ _02269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_41_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09902_ rf_ram.memory\[345\]\[0\] _04905_ _04906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_113_2488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_113_2499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09833_ rf_ram.memory\[61\]\[0\] _04863_ _04864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_133_clk_I clknet_5_24__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06210__A2 _01770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09764_ _04804_ net25 _04821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA_clkbuf_leaf_13_clk_I clknet_5_2__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06976_ _03014_ _03044_ _03045_ _00124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08715_ rf_ram.memory\[150\]\[0\] _04143_ _04144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_154_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05927_ rf_ram.memory\[102\]\[0\] _01631_ _02004_ _02123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09695_ net128 _04767_ _04768_ net129 _04773_ _04774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA_clkbuf_leaf_148_clk_I clknet_5_26__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08646_ _04097_ _04099_ _04101_ _00738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05858_ rf_ram.memory\[224\]\[0\] _01846_ _01956_ _02054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_95_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_68_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07710__A2 _02997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_159_3348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_28_clk_I clknet_5_3__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05789_ _01983_ _01984_ _01928_ _01985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08577_ _04026_ _04054_ _04056_ _00714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_166_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_166_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_1190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_1070 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_176_3662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_1032 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07528_ _03359_ _03393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_25_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_147_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_91_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07459_ _02954_ _03101_ _03349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_14_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06277__A2 _01958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_137_2934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_137_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_1106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10470_ _00214_ clknet_leaf_100_clk rf_ram.memory\[425\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_output190_I net190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_40_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_135_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_40_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_1139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_162_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07226__A1 _02728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06029__A2 _01538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09129_ rf_ram.memory\[92\]\[1\] _04398_ _04402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_60_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08974__A1 _04298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_124_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08726__A1 _04126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11022_ _00759_ clknet_leaf_41_clk rf_ram.memory\[39\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_99_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_95_1115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_86_2001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_339_clk clknet_5_0__leaf_clk clknet_leaf_339_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09151__A1 _02908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05712__A1 _01768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_1121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10806_ _00550_ clknet_leaf_322_clk rf_ram.memory\[553\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05811__B _01916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_1143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_60_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06268__A2 _01501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10737_ _00481_ clknet_leaf_50_clk rf_ram.memory\[458\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_125_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_1198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10668_ _00412_ clknet_leaf_108_clk rf_ram.memory\[377\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_153_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_97_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10599_ _00343_ clknet_leaf_106_clk rf_ram.memory\[318\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_51_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08965__A1 _03008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput107 net107 o_dbus_dat[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput118 net118 o_dbus_dat[28] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__06425__C1 _01625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput129 net129 o_dbus_dat[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__05779__A1 _01972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_58_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06440__A2 _01513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_1250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_75_1793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06830_ rf_ram.memory\[304\]\[0\] _02947_ _02948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05772__I _01918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07940__A2 _02869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06761_ _02876_ _02895_ _02897_ _00057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05951__A1 _01526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06089__B _01707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05712_ _01768_ _01894_ _01907_ net254 _01908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_08500_ _02953_ _04005_ _04006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09480_ _04616_ _04617_ _04618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06692_ _02788_ _02846_ _02850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_77_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_176_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_1065 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08431_ _03689_ _03956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_05643_ rf_ram.memory\[502\]\[0\] _01662_ _01504_ _01839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_175_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05721__B _01916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08362_ _03887_ _03910_ _03912_ _00643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_86_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05574_ _01530_ _01770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_86_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_22_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_738 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_22_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07313_ rf_ram.memory\[256\]\[0\] _03258_ _03259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06259__A2 _01666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07456__A1 _03323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_1318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08293_ _03230_ _02781_ _03869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_154_3256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_1287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_1249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07244_ rf_ram.memory\[421\]\[1\] _03213_ _03215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_171_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_61_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_171_3570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_171_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_5_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_115_2528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07175_ rf_ram.memory\[482\]\[0\] _03172_ _03173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_115_2539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_132_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_1172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_83_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08956__A1 _04266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_132_2853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06126_ rf_ram.memory\[300\]\[1\] _01863_ _01848_ rf_ram.memory\[301\]\[1\] _01773_
+ rf_ram.memory\[303\]\[1\] _02321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_83_1063 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06057_ rf_ram.memory\[380\]\[1\] _01666_ _01645_ rf_ram.memory\[381\]\[1\] _01646_
+ rf_ram.memory\[383\]\[1\] _02252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_2_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06431__A2 _01915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08708__A1 _04129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input47_I i_ibus_rdt[22] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08184__A2 _02846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09816_ _04840_ _04851_ _04853_ _01156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_185_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06195__A1 _01769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09747_ net114 _04790_ _04791_ net115 _04809_ _04810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_0_119_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06959_ rf_ram.memory\[230\]\[1\] _03032_ _03034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_178_3702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09133__A1 _04397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09678_ _04737_ _04758_ _04759_ _04760_ _04761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_179_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07695__A1 _02917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08629_ _04062_ _04088_ _04090_ _00732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_55_1176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11640_ net109 net181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_64_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_147_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05350__C _01495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_175_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11571_ _01303_ clknet_leaf_30_clk rf_ram.memory\[210\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_52_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10522_ _00266_ clknet_leaf_194_clk rf_ram.memory\[268\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_80_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10453_ _00197_ clknet_leaf_187_clk rf_ram.memory\[482\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_123_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_1201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06462__B _01599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10384_ _00128_ clknet_leaf_277_clk rf_ram.memory\[227\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06181__C net253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_102_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11005_ _00742_ clknet_leaf_338_clk rf_ram.memory\[160\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_53_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_1181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05394__C1 _01539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05933__A1 _01569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09124__A1 _02838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_172_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_133_1108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_29_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_1232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_1243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07438__A1 _03326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_16_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_99_2236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_40_clk clknet_5_7__leaf_clk clknet_leaf_40_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_126_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07989__A2 _02960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06110__A1 _01603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05290_ _01434_ _01438_ _01486_ _01487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_130_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_141_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_181_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_1204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_2_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_77_1822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_77_1833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08938__A1 _04269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_1214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07610__A1 _03422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06413__A2 _01787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08980_ rf_ram.memory\[116\]\[1\] _04307_ _04309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_110_2436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_110_2447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07931_ rf_ram.memory\[440\]\[0\] _03642_ _03643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_139_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07862_ _03590_ _03598_ _03600_ _00455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09601_ cpu.immdec.imm24_20\[4\] _04700_ _04710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06813_ _02800_ _02935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_155_1322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07793_ rf_ram.memory\[436\]\[1\] _03555_ _03558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_39_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09532_ _04656_ _04657_ _04658_ _01067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_06744_ _02873_ _02884_ _02885_ _00052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_108_2398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09666__A2 net24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07677__A1 _02923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09463_ net81 net82 _04604_ _04608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06675_ _02785_ _02810_ _02837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_176_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_94_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08414_ _03922_ _03942_ _03944_ _00663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05626_ rf_ram.memory\[489\]\[0\] _01626_ _01822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_175_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_173_3610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09394_ net219 _04561_ _04564_ net220 _04570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_47_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07429__A1 _02923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08345_ _03887_ _03899_ _03901_ _00637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05557_ rf_ram.memory\[268\]\[0\] _01644_ _01645_ rf_ram.memory\[269\]\[0\] _01636_
+ rf_ram.memory\[271\]\[0\] _01753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_0_7_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_163_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_31_clk clknet_5_6__leaf_clk clknet_leaf_31_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_184_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_163_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08276_ rf_ram.memory\[195\]\[1\] _03857_ _03859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_149_1159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05488_ _01550_ _01684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_105_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07227_ rf_ram.memory\[424\]\[0\] _03204_ _03205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_131_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08929__A1 net244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05860__B1 _01953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07158_ _03161_ _03159_ _03162_ _00189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_113_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06109_ rf_ram.memory\[284\]\[1\] _01634_ _01678_ rf_ram.memory\[285\]\[1\] _01625_
+ rf_ram.memory\[287\]\[1\] _02304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__06404__A2 _01863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_993 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07089_ _03087_ _03117_ _03118_ _00164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_121_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_125_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_121_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_98_clk clknet_5_14__leaf_clk clknet_leaf_98_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_35_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_1142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_35_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09354__B2 net232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05376__C1 _01521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09106__A1 _04367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05391__A2 _01502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_1058 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07668__A1 _03455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_84_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06457__B _01503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05679__B1 _01646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09409__A2 _01437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11623_ net73 net145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_108_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_108_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_22_clk clknet_5_3__leaf_clk clknet_leaf_22_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08093__A1 _02843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11554_ _01286_ clknet_leaf_113_clk rf_ram.memory\[451\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_25_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10505_ _00249_ clknet_leaf_197_clk rf_ram.memory\[256\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07840__A1 _03557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06192__B _01860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11485_ _01217_ clknet_leaf_124_clk rf_ram.memory\[464\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_94_2144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05587__I _01550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_880 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10436_ _00180_ clknet_leaf_223_clk rf_ram.memory\[486\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_150_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_55_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_993 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_55_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10367_ _00111_ clknet_leaf_275_clk rf_ram.memory\[228\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_72_1730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_72_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10298_ _00042_ clknet_leaf_316_clk rf_ram.memory\[521\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_89_clk clknet_5_11__leaf_clk clknet_leaf_89_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09896__A2 _03253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05906__A1 _01768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_1063 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05382__A2 _01524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_1182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_1193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06460_ rf_ram.memory\[50\]\[1\] _01499_ _01518_ rf_ram.memory\[51\]\[1\] _01655_
+ rf_ram.memory\[49\]\[1\] _02655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_157_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_133_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05411_ _01518_ _01607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_185_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_172_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_157_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06391_ _02583_ _02585_ _01978_ _02586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_44_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_13_clk clknet_5_2__leaf_clk clknet_leaf_13_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_151_3204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08130_ _03757_ _03766_ _03768_ _00555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_141_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05342_ _01537_ _01538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_83_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_32_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08061_ _03724_ _03722_ _03725_ _00529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_113_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07831__A1 _02945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05273_ _01470_ _01471_ _01472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_113_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05497__I _01550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07012_ _02738_ _02917_ _03068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05842__B1 _01636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_1143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_84_1180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06398__A1 _01769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_149_3155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10194__A2 _02923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_149_3166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_1099 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08963_ _04269_ _04295_ _04297_ _00859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_166_3480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07914_ _03622_ _03630_ _03632_ _00475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08894_ _04234_ _04254_ _04255_ _00832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_75_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_75_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07845_ _03359_ _03590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_127_2752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_127_2763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_162_3399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07776_ _03524_ _03544_ _03546_ _00423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09639__A2 _04507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09515_ cpu.immdec.imm31 _04644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_6_1209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06727_ _02819_ _02873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_151_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_149_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_79_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_91_1184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_177_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09446_ net73 net74 _04593_ _04599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_52_1146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06658_ rf_ram.memory\[347\]\[0\] _02823_ _02824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_140_2996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06322__A1 _01600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_1179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_849 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05609_ _01503_ _01805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_176_495 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06873__A2 _02941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09377_ _04560_ _01010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_46_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06589_ _02748_ _02767_ _02769_ _00013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_81_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08075__A1 _03721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08328_ rf_ram.memory\[21\]\[1\] _03889_ _03891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_145_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08259_ rf_ram.memory\[526\]\[1\] _03846_ _03848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_22_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11270_ _01005_ clknet_leaf_247_clk net205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_104_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10221_ _05078_ _05101_ _05102_ _01313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_186_3845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_max_cap247_I _02774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_1298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_186_3856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output78_I net78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10152_ _02831_ _02894_ _05060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07050__A2 _03089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09327__A1 _04466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10083_ rf_ram.memory\[350\]\[1\] _05015_ _05018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_50_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05349__C1 _01539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05364__A2 _01511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06561__A1 _01353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_1202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10985_ _00722_ clknet_leaf_339_clk rf_ram.memory\[165\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_97_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_139_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_1235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_1246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_736 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_48_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_167_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_155_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_48_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_154_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_183_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08066__A1 _03724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11606_ cpu.decode.co_mem_word net136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_0_1320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09802__A2 _04004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_136_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11537_ _01269_ clknet_leaf_110_clk rf_ram.memory\[312\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__07813__A1 _03554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_1310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_1137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05824__B1 _02019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11468_ _01200_ clknet_leaf_174_clk rf_ram.memory\[342\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_123_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10419_ _00163_ clknet_leaf_183_clk rf_ram.memory\[491\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11399_ _01131_ clknet_leaf_227_clk net114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__08421__I _03902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05960_ _02147_ _02150_ _01599_ _02155_ _02156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
Xclkbuf_leaf_2_clk clknet_5_1__leaf_clk clknet_leaf_2_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_139_1114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_119_Right_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_144_3063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05891_ rf_ram.memory\[70\]\[0\] _01719_ _01925_ rf_ram.memory\[71\]\[0\] _01912_
+ rf_ram.memory\[69\]\[0\] _02087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XTAP_TAPCELL_ROW_144_3074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07630_ _02882_ _03089_ _03456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08541__A2 _03949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_105_2346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_105_2357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07561_ _02935_ _02917_ _03413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_159_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_75_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_85_1976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09300_ _04463_ _04514_ _04515_ _00978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_122_2660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06512_ _01469_ cpu.decode.opcode\[1\] _02701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_122_2671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_85_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07492_ _03360_ _03368_ _03370_ _00315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10100__A2 _03083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09231_ rf_ram.memory\[329\]\[0\] _04464_ _04465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_146_635 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06443_ rf_ram.memory\[32\]\[1\] _01682_ _01601_ _02638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_8_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_173_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06374_ rf_ram.memory\[252\]\[1\] _01677_ _01678_ rf_ram.memory\[253\]\[1\] _01625_
+ rf_ram.memory\[255\]\[1\] _02569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_09162_ net235 _04418_ _04422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_17_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_173_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05325_ _01520_ _01521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_08113_ rf_ram.memory\[554\]\[1\] _03755_ _03758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_72_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09093_ rf_ram.memory\[97\]\[0\] _04378_ _04379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05815__B1 _01772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08044_ _03690_ _03712_ _03714_ _00523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_47_1248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05256_ _01342_ _01455_ _01456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07280__A2 _02992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_168_3520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05187_ _01386_ _01387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XANTENNA__10167__A2 _03547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09995_ _04953_ _04961_ _04963_ _01226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_110_771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_164_3439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_980 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08946_ _04266_ _04286_ _04287_ _00852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_181_3753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08877_ net237 _04077_ _04245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_98_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_4_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07828_ _03554_ _03578_ _03579_ _00442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_4_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05346__A2 _01524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07759_ _03521_ _03535_ _03536_ _00416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_output116_I net116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_165_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10770_ _00514_ clknet_leaf_304_clk rf_ram.memory\[571\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09429_ net95 net96 _02707_ _04590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_48_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_1321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_151_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_180_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_43_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09796__A1 _04840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_188_3907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11322_ _01055_ clknet_leaf_253_clk net88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_22_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11253_ _00989_ clknet_leaf_150_clk rf_ram.memory\[309\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_120_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06470__B _01493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10204_ _03892_ _02866_ _05092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08220__A1 _03823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11184_ _00920_ clknet_leaf_56_clk rf_ram.memory\[92\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10135_ rf_ram.memory\[454\]\[1\] _05047_ _05050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_100_281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06782__A1 _02873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10066_ rf_ram.memory\[307\]\[1\] _05005_ _05007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_89_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09571__I1 net53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05814__B _01505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05337__A2 _01532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_1000 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_1022 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05742__C1 _01811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_67_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_187_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_67_1651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_1066 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_58_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08287__A1 _03855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10968_ _00705_ clknet_leaf_188_clk rf_ram.memory\[489\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_58_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10094__A1 _05017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06298__B1 _01520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_156_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_100_2254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10899_ _00643_ clknet_leaf_14_clk rf_ram.memory\[183\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_100_2265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08039__A1 _03690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_80_1884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_80_1895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09787__A1 _04634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_1150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_5_2__f_clk_I clknet_3_0_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09448__S _04593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06090_ rf_ram.memory\[332\]\[1\] _01709_ _01715_ rf_ram.memory\[333\]\[1\] _01713_
+ rf_ram.memory\[335\]\[1\] _02285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_40_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06380__B _01597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_146_3103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08211__A1 _03787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_1183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_146_3114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_13_Left_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06222__B1 _01778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_1167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08800_ _04167_ _04196_ _04197_ _00796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08762__A2 _04152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09780_ net244 _04067_ _04831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06992_ _03055_ _02894_ _03056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06773__A1 _02873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_7_Right_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_77_1208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08731_ rf_ram.memory\[148\]\[0\] _04153_ _04154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05943_ rf_ram.memory\[34\]\[0\] _01605_ _01624_ rf_ram.memory\[35\]\[0\] _02138_
+ _02139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XTAP_TAPCELL_ROW_124_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08514__A2 _03949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08662_ _02916_ _04078_ _04111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09711__B2 net103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_1_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05874_ rf_ram.memory\[248\]\[0\] _01863_ _01793_ rf_ram.memory\[249\]\[0\] _01696_
+ rf_ram.memory\[251\]\[0\] _02070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_178_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07613_ _02800_ _03445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_156_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08593_ _02805_ _04067_ _04068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_95_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_120_2619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07544_ rf_ram.memory\[320\]\[1\] _03401_ _03403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_147_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08278__A1 _03230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_1203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_22_Left_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10085__A1 _02916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07475_ _03359_ _03360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_158_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09214_ net240 _04418_ _04454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_118_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06426_ rf_ram.memory\[106\]\[1\] _01989_ _01783_ _02621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_174_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_106_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_162_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09145_ _04401_ _04409_ _04411_ _00927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06357_ rf_ram.memory\[233\]\[1\] _01515_ _02552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_72_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_20_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09242__A3 net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_20_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05308_ _01503_ _01504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__08450__A1 cpu.state.genblk1.misalign_trap_sync_r vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06288_ _02481_ _02482_ _01978_ _02483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_09076_ _04367_ _04365_ _04368_ _00901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_130_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_135_2895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_163_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_114_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08027_ _03686_ _03703_ _03704_ _00516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_102_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05239_ _01434_ _01438_ _01439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_25_1321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_31_Left_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_130_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08753__A2 _04152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_301_clk_I clknet_5_6__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09978_ _04400_ _04953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__06764__A1 _02881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08929_ net244 _04038_ _04277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_output233_I net233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08505__A2 _01491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_1032 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_316_clk_I clknet_5_5__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_1027 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_169_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10822_ _00566_ clknet_leaf_321_clk rf_ram.memory\[545\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_95_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08269__A1 _03852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_45_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10753_ _00497_ clknet_leaf_129_clk rf_ram.memory\[47\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_137_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10684_ _00428_ clknet_leaf_80_clk rf_ram.memory\[436\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_168_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_180_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_164_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_1093 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08441__A1 _03953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_1313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11305_ _01038_ clknet_leaf_252_clk net70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__06452__B1 _01609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08992__A2 _04303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_1129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_120_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05809__B _02004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11236_ _00972_ clknet_leaf_257_clk cpu.genblk3.csr.mcause3_0\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_120_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10000__A1 _04953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09941__A1 _04918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11167_ _00903_ clknet_leaf_296_clk rf_ram.memory\[57\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_140_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06755__A1 _02773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10118_ rf_ram.memory\[373\]\[1\] _05037_ _05039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_175_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11098_ _00834_ clknet_leaf_99_clk rf_ram.memory\[429\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05963__C1 _01617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_141_3011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_141_3022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10049_ rf_ram.memory\[306\]\[0\] _04996_ _04997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07315__I _03017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05590_ _01695_ _01786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_82_1924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05730__A2 _01918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10067__A1 _04985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06375__B _01783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07260_ _03017_ _03225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__07483__A2 _03101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_27_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06211_ rf_ram.memory\[396\]\[1\] _01711_ _01772_ rf_ram.memory\[397\]\[1\] _01773_
+ rf_ram.memory\[399\]\[1\] _02406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_143_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07191_ _03157_ _03181_ _03182_ _00202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_14_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_1212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06142_ rf_ram.memory\[304\]\[1\] _01799_ _01602_ _02337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_14_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_1208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_53_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_130_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_117_2570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_1207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_293_clk clknet_5_7__leaf_clk clknet_leaf_293_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_06073_ rf_ram.memory\[345\]\[1\] _01626_ _02268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_111_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06994__A1 _03050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05797__A2 _01664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09901_ _03319_ _02984_ _04905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_112_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_888 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_113_2489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_6_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09832_ _03668_ _02960_ _04863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_171_Right_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05549__A2 _01687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06746__A1 _02876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09763_ _04820_ _01136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06975_ rf_ram.memory\[427\]\[0\] _03044_ _03045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_20_1251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08714_ _03008_ _04078_ _04143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05926_ _02118_ _02119_ _02120_ _02121_ _01860_ _02122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_20_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09694_ _04740_ net32 _04773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_83_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08645_ rf_ram.memory\[519\]\[1\] _04099_ _04101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_179_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05706__C1 _01763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05857_ _02050_ _02052_ _01564_ _02053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_90_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07171__A1 _03157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_159_3349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_179_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08576_ rf_ram.memory\[16\]\[1\] _04054_ _04056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_77_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_178_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_166_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05721__A2 _01915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05788_ rf_ram.memory\[138\]\[0\] _01606_ _01608_ rf_ram.memory\[139\]\[0\] _01702_
+ rf_ram.memory\[137\]\[0\] _01984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_49_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10058__A1 _02821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07527_ _03389_ _03391_ _03392_ _00328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_176_3663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_181_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_1112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07458_ _03326_ _03346_ _03348_ _00303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08671__A1 _04097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_137_2935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_137_2946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_146_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05485__A1 _01675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_107_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06409_ rf_ram.memory\[116\]\[1\] _01510_ _02604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_1129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_40_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07389_ _03292_ _03303_ _03305_ _00277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_40_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09128_ _04400_ _04401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__07226__A2 _03040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output183_I net183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_284_clk clknet_5_18__leaf_clk clknet_leaf_284_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09059_ _04334_ _04355_ _04357_ _00895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_102_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05629__B _01693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_128_1190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06985__A1 _02766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05788__A2 _01606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_240_clk_I clknet_5_21__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09923__A1 _04911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11021_ _00758_ clknet_leaf_330_clk rf_ram.memory\[153\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_25_1173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_1015 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06198__C1 _01713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1037 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_86_2002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05364__B _01552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_255_clk_I clknet_5_20__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06179__C _01670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09151__A2 _04077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_639 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_1183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10805_ _00549_ clknet_leaf_321_clk rf_ram.memory\[554\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_67_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_60_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_60_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10736_ _00480_ clknet_leaf_50_clk rf_ram.memory\[458\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08662__A1 _02916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_1207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_969 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10667_ _00411_ clknet_leaf_96_clk rf_ram.memory\[396\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08414__A1 _03922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_97_2197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10598_ _00342_ clknet_leaf_106_clk rf_ram.memory\[318\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05228__A1 _01375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_275_clk clknet_5_16__leaf_clk clknet_leaf_275_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__10221__A1 _05078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06425__B1 _01702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08965__A2 _04038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput108 net108 o_dbus_dat[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput119 net119 o_dbus_dat[29] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__06976__A1 _03014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_181_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_208_clk_I clknet_5_19__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_1165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_1127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09914__A1 _04884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_75_1794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11219_ _00955_ clknet_leaf_60_clk rf_ram.memory\[67\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_120_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06728__A1 _02806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput90 net90 o_dbus_adr[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_128_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06760_ rf_ram.memory\[514\]\[1\] _02895_ _02897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_163_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09461__S _04604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05711_ _01897_ _01900_ _01660_ _01906_ _01907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_06691_ _02826_ _02847_ _02849_ _00035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07153__A1 _02883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08430_ _03953_ _03954_ _03955_ _00668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_77_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06884__I _02983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05642_ _01836_ _01837_ _01629_ _01838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__05703__A2 _01801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_153_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08361_ rf_ram.memory\[183\]\[1\] _03910_ _03912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05573_ _01650_ _01769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_46_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_175_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_22_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07312_ _02904_ _03253_ _03258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_08292_ _03855_ _03866_ _03868_ _00617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_119_2610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06113__C1 _01646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_154_3246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_154_3257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07243_ _03190_ _03213_ _03214_ _00222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_15_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_143_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_186_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_171_3571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08405__A1 net236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_115_2529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_144_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07174_ _02894_ _03158_ _03172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_171_596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_131_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_266_clk clknet_5_17__leaf_clk clknet_leaf_266_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_42_775 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06125_ rf_ram.memory\[302\]\[1\] _01770_ _02320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_132_2843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_132_2854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_1184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_160_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06967__A1 _02797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_1037 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06056_ rf_ram.memory\[382\]\[1\] _01641_ _02251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09905__A1 _04887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09435__I _01411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09815_ rf_ram.memory\[7\]\[1\] _04851_ _04853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07392__A1 _03289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_1150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09746_ _04804_ net18 _04809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_06958_ _03014_ _03032_ _03033_ _00118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05942__A2 _01513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_178_3703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05909_ _01909_ _02103_ _02104_ _02105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_55_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09677_ _04739_ _04734_ _04760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_06889_ _02975_ _02985_ _02987_ _00095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08628_ rf_ram.memory\[539\]\[1\] _04088_ _04090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_51_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07695__A2 _03496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08892__A1 _02908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_6_Left_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_55_1188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_1079 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08559_ rf_ram.memory\[499\]\[0\] _04045_ _04046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_64_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08644__A1 _04094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11570_ _01302_ clknet_leaf_285_clk rf_ram.memory\[238\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_64_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10521_ _00265_ clknet_leaf_219_clk rf_ram.memory\[252\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_18_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10452_ _00196_ clknet_leaf_187_clk rf_ram.memory\[482\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09444__I0 net72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10203__A1 _05081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_257_clk clknet_5_20__leaf_clk clknet_leaf_257_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_60_561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_161_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_21_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10383_ _00127_ clknet_leaf_101_clk rf_ram.memory\[426\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_131_950 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_21_948 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06958__A1 _03014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11004_ _00741_ clknet_leaf_338_clk rf_ram.memory\[160\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_53_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_194_clk_I clknet_5_28__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06186__A2 _01697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05394__B1 _01540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_3_6_0_clk clknet_0_clk clknet_3_6_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA_clkbuf_leaf_74_clk_I clknet_5_10__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05933__A2 _02117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09124__A2 _04005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_29_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07135__A1 _03126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05697__A1 _01675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_158_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_89_clk_I clknet_5_11__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_185_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_99_2237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_132_clk_I clknet_5_24__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10719_ _00463_ clknet_leaf_78_clk rf_ram.memory\[446\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_67_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_12_clk_I clknet_5_2__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_181_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_77_1823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_130_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06372__C _01620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_141_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_248_clk clknet_5_21__leaf_clk clknet_leaf_248_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_77_1834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_147_clk_I clknet_5_26__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09060__A1 net241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_27_clk_I clknet_5_3__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_110_2437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05621__A1 _01597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_110_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07930_ _02991_ _03547_ _03642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_139_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_177_1036 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07861_ rf_ram.memory\[40\]\[1\] _03598_ _03600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07374__A1 _03292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06177__A2 _01644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09600_ net48 _04709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06812_ _02930_ _02932_ _02934_ _00071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_78_1166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07792_ _03359_ _03557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__05924__A2 _01989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09531_ _04526_ net37 _04658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06743_ rf_ram.memory\[516\]\[0\] _02884_ _02885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07126__A1 _02883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_108_2399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09462_ _04607_ _01048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_78_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_148_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06674_ _02831_ _02836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__08874__A1 _04234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08413_ rf_ram.memory\[177\]\[1\] _03942_ _03944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_114_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_176_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05625_ rf_ram.memory\[488\]\[0\] _01683_ _01684_ _01821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_173_3600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09393_ _04569_ _01017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_173_3611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_164_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05152__A3 _01344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08344_ rf_ram.memory\[214\]\[1\] _03899_ _03901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07429__A2 _03101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_1172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05556_ rf_ram.memory\[270\]\[0\] _01631_ _01752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_129_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_1240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_1194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_1036 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_149_1149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08275_ _03852_ _03857_ _03858_ _00610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05487_ _01682_ _01683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__06101__A2 _01626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_172_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07226_ _02728_ _03040_ _03204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_14_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_239_clk clknet_5_21__leaf_clk clknet_leaf_239_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08929__A2 _04038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07157_ rf_ram.memory\[484\]\[1\] _03159_ _03162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06108_ rf_ram.memory\[286\]\[1\] _01543_ _02303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07088_ rf_ram.memory\[490\]\[0\] _03117_ _03118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_30_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_121_1024 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06039_ _01351_ _02222_ _02233_ _01362_ _02234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_100_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_35_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09354__A2 _03991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05376__B1 _01517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05915__A2 _01918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09729_ _04797_ _01125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_69_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05642__B _01629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05361__C _01494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_139_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06340__A2 _01531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11622_ net72 net144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_167_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08617__A1 _04058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_13_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11553_ _01285_ clknet_leaf_113_clk rf_ram.memory\[451\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_52_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08093__A2 _03729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09290__A1 _04463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_163_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10504_ _00248_ clknet_leaf_196_clk rf_ram.memory\[256\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11484_ _01216_ clknet_leaf_139_clk rf_ram.memory\[295\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09417__I0 net87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_94_2145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10435_ _00179_ clknet_leaf_209_clk rf_ram.memory\[4\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09042__A1 _04331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_55_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10366_ _00110_ clknet_leaf_275_clk rf_ram.memory\[228\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_55_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_131_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_72_1731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_72_1742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10297_ _00041_ clknet_leaf_269_clk rf_ram.memory\[522\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_1243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06159__A2 _01687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_1318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_69_Left_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07108__A1 _03126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_185_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05410_ _01605_ _01606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_84_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08608__A1 _02731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06390_ rf_ram.memory\[66\]\[1\] _01808_ _02019_ rf_ram.memory\[67\]\[1\] _02584_
+ _02585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_150_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09678__C _04760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_151_3205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05341_ _01536_ _01537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_154_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06095__A1 _01350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_78_Left_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08060_ rf_ram.memory\[564\]\[1\] _03722_ _03725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_43_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05272_ cpu.ctrl.pc cpu.ctrl.pc_plus_4_cy_r _01471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_70_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07831__A2 _03234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07011_ _03053_ _03065_ _03067_ _00137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_148_1193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_70_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07595__A1 _03422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_149_3156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_149_3167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08962_ rf_ram.memory\[11\]\[1\] _04295_ _04297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_166_3470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07913_ rf_ram.memory\[443\]\[1\] _03630_ _03632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_166_3481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08893_ rf_ram.memory\[127\]\[0\] _04254_ _04255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07347__A1 _03260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_87_Left_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07844_ _03587_ _03588_ _03589_ _00448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_127_2753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_127_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07775_ rf_ram.memory\[374\]\[1\] _03544_ _03546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09514_ _03992_ _04643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_17_1212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06726_ _02826_ _02870_ _02872_ _00047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_78_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08847__A1 _04202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09445_ _04598_ _01040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06657_ _02815_ _02822_ _02823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_94_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_140_2997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_164_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_1169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_137_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05608_ _01640_ _01804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_75_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09376_ net210 _04549_ _04552_ net211 _04560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_164_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06588_ rf_ram.memory\[241\]\[1\] _02767_ _02769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_93_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08327_ _03884_ _03889_ _03890_ _00630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_96_Left_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05539_ _01536_ _01735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_34_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_172_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08258_ _03820_ _03846_ _03847_ _00604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_62_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07209_ rf_ram.memory\[262\]\[1\] _03191_ _03194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_105_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09024__A1 net246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08189_ _03668_ _03072_ _03805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_120_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_1232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_162_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_63_1243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10220_ rf_ram.memory\[23\]\[0\] _05101_ _05102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_104_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_186_3846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06389__A2 _01918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10151_ _05049_ _05057_ _05059_ _01286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_30_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10082_ _04400_ _05017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__07338__A1 _02958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_50_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05349__B1 _01540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10984_ _00721_ clknet_leaf_334_clk rf_ram.memory\[165\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_85_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_167_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07510__A1 _03356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_1258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06313__A2 _01677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_48_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_26_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11605_ cpu.bne_or_bge net135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09263__A1 _01484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11536_ _01268_ clknet_leaf_148_clk rf_ram.memory\[311\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_68_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_151_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_145_1322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11467_ _01199_ clknet_leaf_174_clk rf_ram.memory\[342\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_64_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09015__A1 rf_ram.memory\[10\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_1310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10418_ _00162_ clknet_leaf_183_clk rf_ram.memory\[491\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11398_ _01130_ clknet_leaf_228_clk net113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__07577__A1 _02882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05547__B _01684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10349_ _00093_ clknet_leaf_135_clk rf_ram.memory\[301\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_29_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_1051 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_144_3064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05890_ rf_ram.memory\[68\]\[0\] _01510_ _02086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_136_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_144_3075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_1136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_178_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07560_ _03393_ _03410_ _03412_ _00341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_105_2347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08829__A1 _04205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06511_ cpu.alu.i_rs1 cpu.bufreg.c_r _02699_ _02700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_122_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_159_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_85_1977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07491_ rf_ram.memory\[325\]\[1\] _03368_ _03370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_158_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_122_2672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_174_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06304__A2 _01510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_146_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09230_ net249 _02815_ _04464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_146_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06442_ _02634_ _02636_ _01563_ _02637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_115_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_185_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_173_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09161_ _04401_ _04419_ _04421_ _00933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09254__A1 _01356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06373_ rf_ram.memory\[254\]\[1\] _01641_ _02004_ _02568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_127_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_161_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06068__A1 _01600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08112_ _03689_ _03757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_05324_ _01519_ _01520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_09092_ net238 _04339_ _04378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_72_987 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08043_ rf_ram.memory\[567\]\[1\] _03712_ _03714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05255_ _01442_ _01453_ _01454_ _01455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09006__A1 _04301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_168_3510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_142_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_168_3521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_141_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05291__A2 _01434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05186_ cpu.mem_bytecnt\[1\] _01385_ cpu.state.o_cnt\[2\] _01386_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nor3_4
XANTENNA__07568__A1 _03389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09994_ rf_ram.memory\[296\]\[1\] _04961_ _04963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_50_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06240__A1 _01909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09309__A2 _01491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08945_ rf_ram.memory\[449\]\[0\] _04286_ _04287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_32_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_181_3754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08876_ _04237_ _04242_ _04244_ _00825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_99_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input22_I i_dbus_rdt[28] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07827_ rf_ram.memory\[412\]\[0\] _03578_ _03579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_4_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05904__C _01670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06288__B _01978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07758_ rf_ram.memory\[376\]\[0\] _03535_ _03536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06709_ _02820_ _02859_ _02860_ _00042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07689_ _02761_ _03481_ _03493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_177_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_137_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09428_ _04589_ _01032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05503__B1 _01696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09359_ net233 _04549_ _04540_ net203 _04551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_164_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09245__A1 cpu.genblk3.csr.o_new_irq vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_43_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_188_3908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_185_Right_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_5_16__f_clk clknet_3_4_0_clk clknet_5_16__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_22_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11321_ _01054_ clknet_leaf_253_clk net86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_50_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05806__A1 _01552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output90_I net90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05282__A2 cpu.alu.i_rs1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11252_ _00988_ clknet_leaf_77_clk rf_ram.memory\[109\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10203_ _05081_ _05089_ _05091_ _01306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_28_1193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11183_ _00919_ clknet_leaf_304_clk rf_ram.memory\[575\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_101_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10134_ _02747_ _05049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_24_1079 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_89_2044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10065_ _04982_ _05005_ _05006_ _01253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_89_2055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06534__A2 _01366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05742__B1 _01810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_134_1034 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_67_1641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_1652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_1131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10967_ _00704_ clknet_leaf_71_clk rf_ram.memory\[119\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05830__B _01551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_1077 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_167_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10898_ _00642_ clknet_leaf_13_clk rf_ram.memory\[183\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_100_2255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_183_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_182_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09236__A1 _03445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_1885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_26_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07798__A1 _03554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_152_Right_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_135_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11519_ _01251_ clknet_leaf_201_clk rf_ram.memory\[507\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_145_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_1184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_150_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_180_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_146_3104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_146_3115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06991_ _02765_ _03055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_08730_ _03134_ _04152_ _04153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_147_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05942_ rf_ram.memory\[33\]\[0\] _01513_ _02138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_124_2701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08661_ _04097_ _04108_ _04110_ _00744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_1_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05873_ rf_ram.memory\[250\]\[0\] _01989_ _01783_ _02069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_1_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07722__A1 _03488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07612_ _03425_ _03442_ _03444_ _00361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08592_ _03902_ _04067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_88_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07543_ _03389_ _03401_ _03402_ _00334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_89_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_1242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08278__A2 _02894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_158_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10085__A2 _03035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07474_ _02747_ _03359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_146_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09213_ _04434_ _04451_ _04453_ _00953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_147_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06425_ rf_ram.memory\[108\]\[1\] _01634_ _01702_ rf_ram.memory\[109\]\[1\] _01625_
+ rf_ram.memory\[111\]\[1\] _02620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_91_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09144_ rf_ram.memory\[90\]\[1\] _04409_ _04411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_44_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06356_ rf_ram.memory\[232\]\[1\] _01735_ _01551_ _02551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_71_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07789__A1 _03039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_1062 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05307_ rf_ram.i_raddr\[2\] _01503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_4
XTAP_TAPCELL_ROW_20_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09075_ rf_ram.memory\[81\]\[1\] _04365_ _04368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_60_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06287_ rf_ram.memory\[130\]\[1\] _01662_ _01636_ rf_ram.memory\[131\]\[1\] _01610_
+ rf_ram.memory\[129\]\[1\] _02482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XANTENNA__08450__A2 cpu.state.stage_two_req vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_135_2896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08026_ rf_ram.memory\[570\]\[0\] _03703_ _03704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05238_ net134 _01436_ _01437_ _01438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_47_1079 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08202__A2 _03811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05169_ _01353_ cpu.immdec.imm19_12_20\[7\] _01367_ cpu.immdec.imm24_20\[3\] _01372_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_60_1246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09977_ _04950_ _04951_ _04952_ _01219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06764__A2 _02899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07961__A1 _03654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08928_ _04269_ _04274_ _04276_ _00845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_98_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08859_ _04205_ _04231_ _04233_ _00819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_100_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_1164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05724__B1 _01911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10821_ _00565_ clknet_leaf_316_clk rf_ram.memory\[546\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_93_1099 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_149_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_45_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10752_ _00496_ clknet_leaf_128_clk rf_ram.memory\[47\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_137_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_45_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07421__I _03017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10683_ _00427_ clknet_leaf_98_clk rf_ram.memory\[416\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_62_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09218__A1 _04434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_1124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_180_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06481__B _01525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11304_ _01037_ clknet_leaf_252_clk net69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_120_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11235_ _00971_ clknet_leaf_255_clk cpu.genblk3.csr.mcause3_0\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_120_355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_8_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11166_ _00902_ clknet_leaf_296_clk rf_ram.memory\[57\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_105_1180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07952__A1 _02898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10117_ _05014_ _05037_ _05038_ _01273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_11097_ _00002_ clknet_leaf_280_clk cpu.alu.i_rs1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__05963__B1 _01624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_141_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10048_ _03445_ _02923_ _04996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_141_3023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_1107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07704__A1 _03491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_1253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_1264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_82_1914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_82_1925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_156_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09209__A1 net241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_1162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_156_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06210_ rf_ram.memory\[398\]\[1\] _01770_ _02405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_2_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05494__A2 _01687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09459__S _04604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06691__A1 _02826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07190_ rf_ram.memory\[473\]\[0\] _03181_ _03182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_143_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06141_ rf_ram.memory\[308\]\[1\] _01709_ _01715_ rf_ram.memory\[309\]\[1\] _01713_
+ rf_ram.memory\[311\]\[1\] _02336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XANTENNA_clkbuf_5_29__f_clk_I clknet_3_7_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_1258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06391__B _01978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_117_2571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06072_ rf_ram.memory\[344\]\[1\] _01683_ _01615_ _02267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_44_1219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09900_ _04887_ _04902_ _04904_ _01190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08196__A1 _03787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09831_ _04840_ _04860_ _04862_ _01162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_158_1321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06974_ _02781_ _03040_ _03044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09762_ net119 _04766_ _04760_ net121 _04819_ _04820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_0_77_1039 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08713_ _04129_ _04140_ _04142_ _00764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05925_ rf_ram.memory\[104\]\[0\] _01863_ _01793_ rf_ram.memory\[105\]\[0\] _01679_
+ rf_ram.memory\[107\]\[0\] _02121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_179_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09693_ _04772_ _01114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08644_ _04094_ _04099_ _04100_ _00737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_178_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05706__B1 _01656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05856_ rf_ram.memory\[234\]\[0\] _01940_ _01959_ rf_ram.memory\[235\]\[0\] _02051_
+ _02052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_83_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_159_3339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08575_ _04023_ _04054_ _04055_ _00713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05787_ rf_ram.memory\[136\]\[0\] _01922_ _01923_ _01983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_95_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_166_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07526_ rf_ram.memory\[361\]\[0\] _03391_ _03392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_178_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10058__A2 _03158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_176_3653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_176_3664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08120__A1 _02728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07457_ rf_ram.memory\[330\]\[1\] _03346_ _03348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_137_2936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_146_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_137_2947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06682__A1 _02826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06408_ _01768_ _02590_ _02602_ _01362_ _02603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_146_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07388_ rf_ram.memory\[24\]\[1\] _03303_ _03305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_40_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_40_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09127_ _02747_ _04400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_06339_ _02522_ _02526_ _02530_ _02533_ _02534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_162_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09620__A1 _04643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_161_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06434__A1 _01350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09058_ rf_ram.memory\[101\]\[1\] _04355_ _04357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_output176_I net176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06985__A2 _02889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08009_ _03692_ _03693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_41_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_1141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11020_ _00757_ clknet_leaf_330_clk rf_ram.memory\[153\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09384__B1 _04564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09923__A2 _03009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06198__B1 _01721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07934__A1 _03622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05645__B _01526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_86_2003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05380__B _01506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10804_ _00548_ clknet_leaf_321_clk rf_ram.memory\[554\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08111__A1 _03754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07151__I _03013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_60_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_60_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10735_ _00479_ clknet_leaf_77_clk rf_ram.memory\[441\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08662__A2 _04078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_137_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_180_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06673__A1 _02826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10666_ _00410_ clknet_leaf_94_clk rf_ram.memory\[396\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_82_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_458 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10597_ _00341_ clknet_leaf_155_clk rf_ram.memory\[358\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_2_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_97_2198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_180_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05228__A2 _01411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput109 net109 o_dbus_dat[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_146_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_1106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_1290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11218_ _00954_ clknet_leaf_58_clk rf_ram.memory\[67\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_75_1795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput80 net80 o_dbus_adr[23] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__06728__A2 _02846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput91 net91 o_dbus_adr[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_43_1296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07925__A1 _02774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11149_ _00885_ clknet_leaf_69_clk rf_ram.memory\[106\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_50_Left_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_37_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05400__A2 _01367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05710_ _01901_ _01902_ _01904_ _01905_ _01670_ _01906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_76_1050 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06690_ rf_ram.memory\[525\]\[1\] _02847_ _02849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_144_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08350__A1 _03884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07153__A2 _03158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_176_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05641_ rf_ram.memory\[506\]\[0\] _01652_ _01654_ rf_ram.memory\[507\]\[0\] _01715_
+ rf_ram.memory\[505\]\[0\] _01837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_153_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05164__A1 _01363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_175_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08360_ _03884_ _03910_ _03911_ _00642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_176_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05572_ _01660_ _01768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_175_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07061__I _03100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08102__A1 _03724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_22_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07311_ _03013_ _03257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_22_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_1207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08291_ rf_ram.memory\[192\]\[1\] _03866_ _03868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_119_2600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_119_2611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06113__B1 _01645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_154_3247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_300_clk_I clknet_5_7__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07242_ rf_ram.memory\[421\]\[0\] _03213_ _03214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05467__A2 _01662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_154_3258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06664__A1 _02779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_171_3561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_171_3572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05872__C1 _01625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07173_ _03161_ _03169_ _03171_ _00195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_42_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08405__A2 _03903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06124_ _01674_ _02306_ _02318_ _01361_ _02319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_83_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_132_2844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_631 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_132_2855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06967__A2 _02830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_315_clk_I clknet_5_5__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06055_ _02238_ _02242_ _02246_ _02249_ _02250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_140_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_995 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_78_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09814_ _04837_ _04851_ _04852_ _01155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09745_ _04808_ _01130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06957_ rf_ram.memory\[230\]\[0\] _03032_ _03033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_97_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_178_3704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05908_ rf_ram.memory\[118\]\[0\] _01706_ _01911_ rf_ram.memory\[119\]\[0\] _01931_
+ rf_ram.memory\[117\]\[0\] _02104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_06888_ rf_ram.memory\[281\]\[1\] _02985_ _02987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09676_ cpu.bufreg2.o_sh_done_r _04737_ _04759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_90_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08341__A1 _03892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08627_ _04058_ _04088_ _04089_ _00731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05839_ rf_ram.memory\[204\]\[0\] _01649_ _01912_ rf_ram.memory\[205\]\[0\] _01925_
+ rf_ram.memory\[207\]\[0\] _02035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_16_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08892__A2 _04038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_166_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08067__I _03692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08558_ _02865_ _03158_ _04045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_166_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07509_ rf_ram.memory\[323\]\[0\] _03380_ _03381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_147_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08489_ rf_ram.memory\[369\]\[0\] _03998_ _03999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_175_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09841__A1 _02714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06655__A1 _02779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10520_ _00264_ clknet_leaf_224_clk rf_ram.memory\[252\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_91_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_165_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05863__C1 _01968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10451_ _00195_ clknet_leaf_184_clk rf_ram.memory\[495\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09444__I1 net73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10382_ _00126_ clknet_leaf_100_clk rf_ram.memory\[426\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_32_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_33_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_107_Left_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_102_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05630__A2 _01697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07907__A1 _03619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11003_ _00740_ clknet_leaf_338_clk rf_ram.memory\[161\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05375__B _01506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_1072 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_53_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08580__A1 net250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_1183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_70_1692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09361__I _04539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_185_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08883__A2 _04248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06894__A1 _02975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_83_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_184_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_67_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09832__A1 _03668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_99_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_165_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06646__A1 _02736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10718_ _00462_ clknet_leaf_78_clk rf_ram.memory\[446\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09310__B _03967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10649_ _00393_ clknet_leaf_109_clk rf_ram.memory\[382\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_130_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08399__A1 _03922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_77_1824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_141_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_77_1835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_140_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_140_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09060__A2 _04339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05606__C1 _01721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07071__A1 _03092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_110_2438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_110_2449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07860_ _03587_ _03598_ _03599_ _00454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_78_1112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_177_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_1123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06031__C1 _01555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06811_ rf_ram.memory\[290\]\[1\] _02932_ _02934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07791_ _03554_ _03555_ _03556_ _00428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05385__A1 _01495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_1178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_155_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06742_ _02881_ _02883_ _02884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09530_ cpu.immdec.imm19_12_20\[1\] _04649_ _04657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07126__A2 _02997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09461_ net80 net81 _04604_ _04607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06673_ _02826_ _02833_ _02835_ _00031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06334__B1 _02019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_184_clk clknet_5_29__leaf_clk clknet_leaf_184_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_176_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05688__A2 _01697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06885__A1 _02958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08412_ _03919_ _03942_ _03943_ _00662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05624_ _01675_ _01818_ _01819_ _01820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_09392_ net218 _04561_ _04564_ net219 _04569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_173_3601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05304__I _01499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_173_3612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08343_ _03884_ _03899_ _03900_ _00636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05555_ _01738_ _01742_ _01747_ _01750_ _01751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_114_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_1106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06637__A1 _02801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06098__C1 _01678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_15_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08274_ rf_ram.memory\[195\]\[0\] _03857_ _03858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_144_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05486_ _01508_ _01682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_117_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07225_ _03193_ _03201_ _03203_ _00215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_89_1296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05845__C1 _01713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_144_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_254_clk_I clknet_5_20__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05860__A2 _01958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07156_ _03017_ _03161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_06107_ _02299_ _02301_ _01746_ _02302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07062__A1 _03082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07087_ _02775_ _02911_ _03117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA_input52_I i_ibus_rdt[27] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06038_ _02227_ _02232_ _01351_ _02233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_leaf_269_clk_I clknet_5_16__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_121_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_35_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08562__A1 _04026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_29_Right_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07989_ _03672_ _02960_ _03679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09728_ net107 _04790_ _04791_ net108 _04796_ _04797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_0_97_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_175_clk clknet_5_31__leaf_clk clknet_leaf_175_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09659_ net120 _04737_ _04744_ _04740_ _04745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_96_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05679__A2 _01801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_171_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_38_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_207_clk_I clknet_5_24__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11621_ net71 net143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_49_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_65_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_148_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_33_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09814__A1 _04837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_154_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06628__A1 _02797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_13_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_181_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11552_ _01284_ clknet_leaf_112_clk rf_ram.memory\[452\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_135_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_38_Right_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10503_ _00247_ clknet_leaf_202_clk rf_ram.memory\[257\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_162_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11483_ _01215_ clknet_leaf_139_clk rf_ram.memory\[295\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_135_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09417__I1 net90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09557__S _03967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10434_ _00178_ clknet_leaf_211_clk rf_ram.memory\[4\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_94_2146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05851__A2 _01501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10188__A1 _05081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_115_Left_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_122_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10365_ _00109_ clknet_leaf_138_clk rf_ram.memory\[297\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_55_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_1201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_55_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06261__C1 _01645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06800__A1 _02876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10296_ _00040_ clknet_leaf_269_clk rf_ram.memory\[522\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_72_1732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_178_1313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_72_1743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_47_Right_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08553__A1 net249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06013__C1 _01539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05833__B _01928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_124_Left_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_137_1054 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08305__A1 _03852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10112__A1 _05014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_1098 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06867__A1 _02935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_185_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_158_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_1059 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_1205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08608__A2 _02939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_173_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_157_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_56_Right_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_55_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06619__A1 _02748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05340_ _01508_ _01536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_151_3206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_1182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06095__A2 _02278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07292__A1 _03222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05271_ cpu.state.cnt_r\[2\] _01386_ _01470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_109_1101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_133_Left_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_183_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_181_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07010_ rf_ram.memory\[223\]\[1\] _03065_ _03067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_113_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09467__S _04604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_1100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05842__A2 _01662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10179__A1 _05046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_45_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07044__A1 _02829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_122_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08792__A1 net246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_149_3157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08961_ _04266_ _04295_ _04296_ _00858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_149_3168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_65_Right_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_166_3471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07912_ _03619_ _03630_ _03631_ _00474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_166_3482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08892_ _02908_ _04038_ _04254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07843_ rf_ram.memory\[431\]\[0\] _03588_ _03589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_142_Left_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_127_2754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07774_ _03521_ _03544_ _03545_ _00422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09513_ _04642_ _01064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06725_ rf_ram.memory\[51\]\[1\] _02870_ _02872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_157_clk clknet_5_26__leaf_clk clknet_leaf_157_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_67_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06858__A1 _02930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09444_ net72 net73 _04593_ _04598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06656_ _02821_ _02822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_140_2987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_1148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_166_Right_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_140_2998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_74_Right_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_93_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05607_ _01797_ _01798_ _01800_ _01802_ _01717_ _01803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_136_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09375_ _04559_ _01009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_46_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06587_ _02743_ _02767_ _02768_ _00012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_148_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05538_ _01347_ _01732_ _01733_ _01734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_74_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08326_ rf_ram.memory\[21\]\[0\] _03889_ _03890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_34_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_151_Left_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_61_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06086__A2 _01711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08257_ rf_ram.memory\[526\]\[0\] _03846_ _03847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_46_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05469_ rf_ram.memory\[372\]\[0\] _01509_ _01664_ rf_ram.memory\[373\]\[0\] _01519_
+ rf_ram.memory\[375\]\[0\] _01665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XTAP_TAPCELL_ROW_31_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_144_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_43_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_3_5_0_clk clknet_0_clk clknet_3_5_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_07208_ _03017_ _03193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA_clkbuf_leaf_73_clk_I clknet_5_10__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08188_ _03790_ _03802_ _03804_ _00577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_63_1211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09024__A2 _04303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_1245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07139_ rf_ram.memory\[498\]\[1\] _03148_ _03150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_63_1255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_186_3847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_83_Right_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10150_ rf_ram.memory\[451\]\[1\] _05057_ _05059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_88_clk_I clknet_5_11__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10081_ _05014_ _05015_ _05016_ _01259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_100_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_50_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08535__A1 _04026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07338__A2 _02972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_131_clk_I clknet_5_24__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_50_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06010__A2 _01532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_11_clk_I clknet_5_2__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05145__S _01347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_148_clk clknet_5_26__leaf_clk clknet_leaf_148_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_134_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10983_ _00720_ clknet_leaf_331_clk rf_ram.memory\[166\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_69_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_146_clk_I clknet_5_26__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_92_Right_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06849__A1 _02958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_48_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_133_Right_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_clkbuf_leaf_26_clk_I clknet_5_3__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_155_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06484__B _01503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_183_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_167_1003 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_139_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11604_ cpu.bufreg2.o_sh_done_r net125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_136_840 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_183_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_1322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06077__A2 _01697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_163_670 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11535_ _01267_ clknet_leaf_146_clk rf_ram.memory\[311\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_81_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_320_clk clknet_5_5__leaf_clk clknet_leaf_320_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_81_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06482__C1 _01653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05824__A2 _01940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11466_ _01198_ clknet_leaf_168_clk rf_ram.memory\[343\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_81_1322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07026__A1 _03050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10417_ _00161_ clknet_leaf_182_clk rf_ram.memory\[492\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11397_ _01129_ clknet_leaf_228_clk net112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__07577__A2 _03390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06234__C1 _01656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08774__A1 _04167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10348_ _00092_ clknet_leaf_134_clk rf_ram.memory\[301\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10279_ _00023_ clknet_leaf_137_clk rf_ram.memory\[293\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_144_3065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_144_3076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05563__B _01629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06001__A2 _01524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_161_3390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_177_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_105_2348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_139_clk clknet_5_27__leaf_clk clknet_leaf_139_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_06510_ _01382_ cpu.decode.opcode\[1\] _01381_ _02699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07490_ _03356_ _03368_ _03369_ _00314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_5_1200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_122_2662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_85_1978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_152_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_158_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_913 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06441_ rf_ram.memory\[42\]\[1\] _01605_ _01607_ rf_ram.memory\[43\]\[1\] _02635_
+ _02636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_5_1244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_100_Right_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_186_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_150_1073 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_146_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09160_ rf_ram.memory\[88\]\[1\] _04419_ _04421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_111_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06372_ _02563_ _02564_ _02565_ _02566_ _01620_ _02567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_174_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08111_ _03754_ _03755_ _03756_ _00548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05323_ _01518_ _01519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_12
XFILLER_0_173_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09091_ _04367_ _04375_ _04377_ _00907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07265__A1 _03222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_311_clk clknet_5_5__leaf_clk clknet_leaf_311_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_71_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08042_ _03686_ _03712_ _03713_ _00522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_9_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05254_ net98 net105 net128 net114 _01376_ _01375_ _01454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__05815__A2 _01799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07017__A1 _02750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_168_3511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_168_3522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05185_ cpu.mem_bytecnt\[0\] _01385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_101_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05579__A1 _01769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09993_ _04950_ _04961_ _04962_ _01225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08944_ _03672_ _02899_ _04286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09309__A3 _04013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_32_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_122_1197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_181_3755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08875_ rf_ram.memory\[12\]\[1\] _04242_ _04244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07826_ _02839_ _03559_ _03578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_98_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input15_I i_dbus_rdt[21] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07757_ _02991_ _03496_ _03535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05751__A1 _01674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06708_ rf_ram.memory\[521\]\[0\] _02859_ _02860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_17_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07688_ _03491_ _03489_ _03492_ _00389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_67_738 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09427_ net94 net95 _02707_ _04589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_48_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06639_ _02743_ _02807_ _02808_ _00024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_17_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_165_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09358_ _04550_ _01001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_35_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09245__A2 _01413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06059__A2 _01649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08309_ rf_ram.memory\[243\]\[0\] _03878_ _03879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_173_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_302_clk clknet_5_6__leaf_clk clknet_leaf_302_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09289_ rf_ram.memory\[65\]\[0\] _04508_ _04509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_151_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_188_3909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11320_ _01053_ clknet_leaf_264_clk net85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_16_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_166_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11251_ _00987_ clknet_leaf_70_clk rf_ram.memory\[109\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05648__B _01660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output83_I net83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10202_ rf_ram.memory\[191\]\[1\] _05089_ _05091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11182_ _00918_ clknet_leaf_303_clk rf_ram.memory\[575\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10133_ _05046_ _05047_ _05048_ _01279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06231__A2 _01623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10064_ rf_ram.memory\[307\]\[0\] _05005_ _05006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_89_2045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_89_2056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05990__A1 _02102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06479__B _01503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_526 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_159_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_67_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_187_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_67_1653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_1143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10966_ _00703_ clknet_leaf_71_clk rf_ram.memory\[119\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_39_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07495__A1 _03356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06298__A2 _01958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10897_ _00641_ clknet_leaf_13_clk rf_ram.memory\[182\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_100_2256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_156_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_911 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_109_851 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09236__A2 _02909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_1886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06455__C1 _01655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11518_ _01250_ clknet_leaf_200_clk rf_ram.memory\[34\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_180_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_1142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_111_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11449_ _01181_ clknet_leaf_276_clk rf_ram.memory\[239\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08747__A1 net242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_1148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_1125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_146_3105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_146_3116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06222__A2 _01777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06990_ _03053_ _03051_ _03054_ _00129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_163_3430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_186_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_input7_I i_dbus_rdt[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05941_ rf_ram.memory\[32\]\[0\] _01682_ _01550_ _02137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09172__A1 _03071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08660_ rf_ram.memory\[15\]\[1\] _04108_ _04110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05872_ rf_ram.memory\[252\]\[0\] _01677_ _01678_ rf_ram.memory\[253\]\[0\] _01625_
+ rf_ram.memory\[255\]\[0\] _02068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XTAP_TAPCELL_ROW_124_2702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07611_ rf_ram.memory\[353\]\[1\] _03442_ _03444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08591_ _04062_ _04064_ _04066_ _00718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_3_4_0_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07999__I _02742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_163_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07542_ rf_ram.memory\[320\]\[0\] _03401_ _03402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_152_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_5_22__f_clk clknet_3_5_0_clk clknet_5_22__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_76_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_1216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07473_ _03356_ _03357_ _03358_ _00308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_14_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06289__A2 _01770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_45_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09212_ rf_ram.memory\[68\]\[1\] _04451_ _04453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06424_ rf_ram.memory\[110\]\[1\] _01641_ _02004_ _02619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_16_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07238__A1 _03190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06355_ _01951_ _02548_ _02549_ _02550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09143_ _04397_ _04409_ _04410_ _00926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_161_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07789__A2 _03135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08986__A1 _04301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05306_ _01501_ _01502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_45_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09719__I _04766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09074_ _04061_ _04367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_20_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06286_ rf_ram.memory\[128\]\[1\] _01915_ _01923_ _02481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_71_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_135_2897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08025_ _02813_ _03693_ _03703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05237_ rf_ram.rdata\[0\] _01378_ rf_ram_if.rtrig1 _01437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_141_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08738__A1 _01369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05168_ _01369_ _01370_ _01371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__07410__A1 _03292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06213__A2 _01692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09976_ rf_ram.memory\[274\]\[0\] _04951_ _04952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08927_ rf_ram.memory\[124\]\[1\] _04274_ _04276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_99_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_157_1057 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08858_ rf_ram.memory\[131\]\[1\] _04231_ _04233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_93_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07809_ rf_ram.memory\[414\]\[1\] _03566_ _03568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_19_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08789_ _04167_ _04189_ _04190_ _00792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10820_ _00564_ clknet_leaf_316_clk rf_ram.memory\[546\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_79_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07477__A1 _03360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10751_ _00495_ clknet_leaf_51_clk rf_ram.memory\[470\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_45_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10682_ _00426_ clknet_leaf_97_clk rf_ram.memory\[416\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_36_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_62_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_137_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_180_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08977__A1 _03134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06437__C1 _01607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11303_ _01036_ clknet_leaf_252_clk net68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_65_1158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06452__A2 _01633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_1169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11234_ _00970_ clknet_leaf_256_clk cpu.genblk3.csr.mcause3_0\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06204__A2 _01649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07401__A1 _03309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06988__I _03017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11165_ _00901_ clknet_leaf_47_clk rf_ram.memory\[81\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07952__A2 _03158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10116_ rf_ram.memory\[373\]\[0\] _05037_ _05038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11096_ _00833_ clknet_leaf_84_clk rf_ram.memory\[127\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_141_3013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10047_ _04985_ _04993_ _04995_ _01246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_136_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08901__A1 _04237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05841__B _01916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_82_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_82_1926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07468__A1 _03326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10949_ _00687_ clknet_leaf_154_clk rf_ram.memory\[359\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_112_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_70_clk clknet_5_8__leaf_clk clknet_leaf_70_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_183_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09209__A2 _04418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_183_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_1174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_27_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06140_ rf_ram.memory\[310\]\[1\] _01719_ _01707_ _02335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_14_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_186_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_101_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_117_2572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07640__A1 _03458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06071_ _01675_ _02264_ _02265_ _02266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__06443__A2 _01682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_1269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09475__S _04604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_6_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09830_ rf_ram.memory\[62\]\[1\] _04860_ _04862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_10_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_120_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05254__I0 net98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09761_ _04804_ net23 _04819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_06973_ _03018_ _03041_ _03043_ _00123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_20_1231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_77_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09145__A1 _04401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_1253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08712_ rf_ram.memory\[151\]\[1\] _04140_ _04142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05924_ rf_ram.memory\[106\]\[0\] _01989_ _01783_ _02120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09692_ net127 _04767_ _04768_ net128 _04771_ _04772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__05307__I rf_ram.i_raddr\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08643_ rf_ram.memory\[519\]\[0\] _04099_ _04100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05855_ rf_ram.memory\[233\]\[0\] _01515_ _02051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_90_1218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_179_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05751__B _01946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08574_ rf_ram.memory\[16\]\[0\] _04054_ _04055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05786_ _01909_ _01980_ _01981_ _01982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_88_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_117_1074 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07525_ _02752_ _03390_ _03391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07459__A1 _02954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_176_3654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_176_3665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_61_clk clknet_5_9__leaf_clk clknet_leaf_61_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08120__A2 _03729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_91_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_174_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_64_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07456_ _03323_ _03346_ _03347_ _00302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_135_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_1136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_137_2937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06407_ _02593_ _02596_ _01660_ _02601_ _02602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_107_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_137_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07387_ _03289_ _03303_ _03304_ _00276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_106_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08959__A1 net246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_40_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09126_ _04397_ _04398_ _04399_ _00920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06338_ _01972_ _02531_ _02532_ _02533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_32_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06269_ rf_ram.memory\[156\]\[1\] _01614_ _01968_ rf_ram.memory\[157\]\[1\] _01953_
+ rf_ram.memory\[159\]\[1\] _02464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_09057_ _04331_ _04355_ _04356_ _00894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_103_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_130_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08008_ _02730_ _02732_ _02762_ _03692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_124_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_1175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09959_ _04911_ _02954_ _04941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09136__A1 net249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_86_2004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_170_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10803_ _00547_ clknet_leaf_322_clk rf_ram.memory\[555\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_170_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_68_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_138_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_1293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_52_clk clknet_5_9__leaf_clk clknet_leaf_52_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_138_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_60_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_24_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10734_ _00478_ clknet_leaf_77_clk rf_ram.memory\[441\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_137_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_153_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07870__A1 _03587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10665_ _00409_ clknet_leaf_109_clk rf_ram.memory\[378\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_36_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06492__B _01372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10596_ _00340_ clknet_leaf_155_clk rf_ram.memory\[358\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_35_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_97_2199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06425__A2 _01634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_121_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_1123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_142_1178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_75_1785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11217_ _00953_ clknet_leaf_64_clk rf_ram.memory\[68\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_75_1796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_112_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput70 net70 o_dbus_adr[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput81 net81 o_dbus_adr[24] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__07925__A2 _02832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput92 net92 o_dbus_adr[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_11148_ _00884_ clknet_leaf_67_clk rf_ram.memory\[106\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05936__A1 _01903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11079_ _00816_ clknet_leaf_14_clk rf_ram.memory\[132\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07689__A1 _02761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05640_ rf_ram.memory\[504\]\[0\] _01755_ _01756_ _01836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_187_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05164__A2 _01366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_149_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05571_ _01674_ _01751_ _01766_ _01361_ _01767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_86_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_43_clk clknet_5_13__leaf_clk clknet_leaf_43_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_50_1235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07310_ _03225_ _03254_ _03256_ _00247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_22_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_58_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_129_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08290_ _03852_ _03866_ _03867_ _00616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_128_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_119_2601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_119_2612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_154_3248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_1279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07241_ _02795_ _03040_ _03213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_154_3259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_171_3562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_171_3573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05872__B1 _01678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07172_ rf_ram.memory\[495\]\[1\] _03169_ _03171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_54_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06123_ _02309_ _02312_ _01349_ _02317_ _02318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_125_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06416__A2 _01915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_132_2845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_132_2856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06054_ _01527_ _02247_ _02248_ _02249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_41_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06719__A3 _02730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09813_ rf_ram.memory\[7\]\[0\] _04851_ _04852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09744_ net113 _04790_ _04791_ net114 _04807_ _04808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_06956_ _02766_ _02806_ _03032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_20_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05907_ rf_ram.memory\[116\]\[0\] _01510_ _02103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_118_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_1136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09675_ net124 _03976_ _04758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_179_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_178_3705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_154_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06887_ _02970_ _02985_ _02986_ _00094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_97_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_96_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_1135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08341__A2 _03009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08626_ rf_ram.memory\[539\]\[0\] _04088_ _04089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_55_1146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05838_ rf_ram.memory\[206\]\[0\] _01531_ _02034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05155__A2 cpu.decode.co_ebreak vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06352__A1 _01674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06296__C _01362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08557_ _04026_ _04042_ _04044_ _00706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05769_ rf_ram.memory\[146\]\[0\] _01958_ _01953_ rf_ram.memory\[147\]\[0\] _01964_
+ _01965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_49_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_34_clk clknet_5_6__leaf_clk clknet_leaf_34_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_92_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07508_ _03319_ _02889_ _03380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_64_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08488_ net248 _03496_ _03998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_135_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_147_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07852__A1 _03590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07439_ _02921_ _02883_ _03337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05863__B1 _01959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10450_ _00194_ clknet_leaf_184_clk rf_ram.memory\[495\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05500__I _01695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09109_ _04364_ _04387_ _04388_ _00914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10381_ _00125_ clknet_leaf_100_clk rf_ram.memory\[427\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_60_563 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_1128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_130_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_57_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09357__A1 net232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09357__B2 net233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11002_ _00739_ clknet_5_0__leaf_clk rf_ram.memory\[161\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_102_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_53_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09109__A1 _04364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_1173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08580__A2 _03949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05394__A2 _01544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_70_1693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05391__B _01506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_73_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_1219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_184_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_25_clk clknet_5_3__leaf_clk clknet_leaf_25_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_28_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_166_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09832__A2 _02960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_99_2239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06646__A2 _02799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10717_ _00461_ clknet_leaf_51_clk rf_ram.memory\[463\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_153_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_1321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_130_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10648_ _00392_ clknet_leaf_109_clk rf_ram.memory\[382\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_67_1039 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05410__I _01605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_183_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_530 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_738 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_77_1825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_114_2520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_77_1836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10579_ _00323_ clknet_leaf_159_clk rf_ram.memory\[323\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05606__B1 _01726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_121_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_110_2439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05566__B _01526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08020__A1 _02822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05909__A1 _01909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06031__B1 _01554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06810_ _02927_ _02932_ _02933_ _00070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07790_ rf_ram.memory\[436\]\[0\] _03555_ _03556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_78_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06582__A1 cpu.immdec.imm11_7\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_147_Right_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_39_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06741_ net241 _02883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_79_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09460_ _04606_ _01047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06672_ rf_ram.memory\[455\]\[1\] _02833_ _02835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_176_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08411_ rf_ram.memory\[177\]\[0\] _03942_ _03943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_114_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05623_ rf_ram.memory\[492\]\[0\] _01677_ _01793_ rf_ram.memory\[493\]\[0\] _01679_
+ rf_ram.memory\[495\]\[0\] _01819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_153_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06885__A2 _02984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09391_ _04568_ _01016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_59_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_173_3602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_16_clk clknet_5_2__leaf_clk clknet_leaf_16_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_173_3613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_171_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_1139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_47_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08087__A1 _03724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08342_ rf_ram.memory\[214\]\[0\] _03899_ _03900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_80_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05554_ _01603_ _01748_ _01749_ _01750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_129_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_1005 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_163_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1065 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06098__B1 _01679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_1129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05485_ _01675_ _01676_ _01680_ _01681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__06637__A2 _02806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_15_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08273_ _03230_ _02889_ _03857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_15_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05845__B1 _01721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07224_ rf_ram.memory\[425\]\[1\] _03201_ _03203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_27_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05320__I _01515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07155_ _03157_ _03159_ _03160_ _00188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_5_13__f_clk_I clknet_3_3_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_113_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06106_ rf_ram.memory\[282\]\[1\] _01687_ _01679_ rf_ram.memory\[283\]\[1\] _02300_
+ _02301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__07062__A2 _03101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07086_ _03092_ _03114_ _03116_ _00163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_112_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05476__B _01660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06037_ _02228_ _02229_ _02230_ _02231_ _01564_ _02232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_61_1150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_1026 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_1037 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_1292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input45_I i_ibus_rdt[20] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_100_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_35_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05376__A2 _01511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06573__A1 _02748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07988_ _03654_ _03676_ _03678_ _00503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_114_Right_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09727_ _04781_ net11 _04796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_06939_ rf_ram.memory\[228\]\[1\] _03020_ _03022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05781__C1 _01610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09511__A1 _04637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_179_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_1039 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09658_ _04737_ _03975_ _04743_ _04744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_85_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06100__B _01615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_166_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08609_ _04077_ _04078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_96_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_1133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09589_ _03967_ _04700_ _04701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_49_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_78_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11620_ net70 net142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_182_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_1252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08078__A1 _02945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07825__A1 _03557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11551_ _01283_ clknet_leaf_111_clk rf_ram.memory\[452\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06628__A2 _02799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_1296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_64_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10502_ _00246_ clknet_leaf_202_clk rf_ram.memory\[257\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11482_ _01214_ clknet_leaf_167_clk rf_ram.memory\[335\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_52_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_59_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_94_2136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_738 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10433_ _00177_ clknet_leaf_225_clk rf_ram.memory\[487\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_94_2147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_150_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08250__A1 _03823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10364_ _00108_ clknet_leaf_138_clk rf_ram.memory\[297\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_27_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_55_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06261__B1 _01646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05386__B _01505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10295_ _00039_ clknet_leaf_269_clk rf_ram.memory\[523\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_72_1733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_72_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06013__B1 _01540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09750__A1 net115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08553__A2 _03158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09750__B2 net116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_5_3__f_clk clknet_3_0_0_clk clknet_5_3__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_137_1077 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06010__B _01505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05405__I rf_ram.i_raddr\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_107_2390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_158_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_314_clk_I clknet_5_5__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06867__A2 _02972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_173_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_185_1318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07816__A1 _02959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_151_3207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_329_clk_I clknet_5_4__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05270_ cpu.decode.opcode\[0\] _01469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_71_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_154_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_1194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09569__A1 _04478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_1071 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_1135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_1172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07044__A2 _03089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_1134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08241__A1 _03668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08792__A2 _04152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08960_ rf_ram.memory\[11\]\[0\] _04295_ _04296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_149_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_5_clk clknet_5_1__leaf_clk clknet_leaf_5_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_149_3169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07911_ rf_ram.memory\[443\]\[0\] _03630_ _03631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_166_3472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08891_ _04237_ _04251_ _04253_ _00831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_166_3483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07842_ _02953_ _03234_ _03588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__06555__A1 _01353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_1111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_127_2755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05743__C _01658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07773_ rf_ram.memory\[374\]\[0\] _03544_ _03545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_155_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09512_ cpu.genblk3.csr.timer_irq_r _04471_ _04473_ _04642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06724_ _02820_ _02870_ _02871_ _00046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_78_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_177_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_1214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05315__I _01510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_149_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09443_ _04597_ _01039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_177_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06655_ _02779_ _02811_ _02821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_91_1176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_140_2988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_176_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05606_ rf_ram.memory\[306\]\[0\] _01801_ _01726_ rf_ram.memory\[307\]\[0\] _01721_
+ rf_ram.memory\[305\]\[0\] _01802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XTAP_TAPCELL_ROW_140_2999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09374_ net209 _04549_ _04552_ net210 _04559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_176_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06586_ rf_ram.memory\[241\]\[0\] _02767_ _02768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_19_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08325_ _03035_ _03072_ _03889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_19_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05537_ cpu.immdec.imm24_20\[2\] _01367_ _01733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_75_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_1072 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08256_ _02845_ _02972_ _03846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_144_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08480__A1 _02713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05468_ _01514_ _01664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_31_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_989 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07207_ _03190_ _03191_ _03192_ _00208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08187_ rf_ram.memory\[540\]\[1\] _03802_ _03804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_132_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05399_ cpu.immdec.imm19_12_20\[7\] _01595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_160_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07138_ _03123_ _03148_ _03149_ _00182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_186_3848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06243__B1 _01857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09980__A1 _04953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07069_ _03087_ _03105_ _03106_ _00156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06794__A1 _02773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output151_I net151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10080_ rf_ram.memory\[350\]\[0\] _05015_ _05016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_50_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05349__A2 _01544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06546__B2 _01347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10982_ _00719_ clknet_leaf_331_clk rf_ram.memory\[166\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06849__A2 _02960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_1238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_48_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_183_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_155_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09799__A1 _04837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11534_ _01266_ clknet_leaf_191_clk rf_ram.memory\[351\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08471__A1 _02714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_163_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_52_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06482__B1 _01714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11465_ _01197_ clknet_leaf_168_clk rf_ram.memory\[343\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_123_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_888 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08223__A1 _03820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10416_ _00160_ clknet_leaf_182_clk rf_ram.memory\[492\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_111_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11396_ _01128_ clknet_leaf_226_clk net111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_150_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_21_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06234__B1 _01763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09971__A1 _04918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10347_ _00091_ clknet_leaf_179_clk rf_ram.memory\[282\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_104_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05588__A2 _01782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06005__B _01505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10278_ _00022_ clknet_leaf_136_clk rf_ram.memory\[293\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_104_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09574__I1 net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05844__B _01805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_109_2430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_144_3066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_144_3077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_161_3380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_161_3391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_253_clk_I clknet_5_20__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_105_2349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10097__A1 _05014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_17_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_158_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_85_1979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_122_2663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06440_ rf_ram.memory\[41\]\[1\] _01513_ _02635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_173_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05512__A2 _01706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06170__C1 _01636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_5_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_174_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_111_1036 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_268_clk_I clknet_5_16__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_56_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06371_ rf_ram.memory\[242\]\[1\] _01606_ _01625_ rf_ram.memory\[243\]\[1\] _01702_
+ rf_ram.memory\[241\]\[1\] _02566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_17_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08110_ rf_ram.memory\[554\]\[0\] _03755_ _03756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_56_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05322_ _01512_ _01498_ _01518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_71_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_83_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_127_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_1177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09090_ rf_ram.memory\[569\]\[1\] _04375_ _04377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_160_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_16_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08041_ rf_ram.memory\[567\]\[0\] _03712_ _03713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06473__B1 _01624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05253_ _01385_ _01452_ cpu.mem_bytecnt\[1\] _01453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_86_1278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_3_0_0_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_168_3512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05184_ cpu.state.cnt_r\[0\] _01384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XTAP_TAPCELL_ROW_168_3523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10021__A1 _03309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09992_ rf_ram.memory\[296\]\[0\] _04961_ _04962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_12_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06776__A1 _02779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_110_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08943_ _04269_ _04283_ _04285_ _00851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_leaf_206_clk_I clknet_5_24__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_1165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_32_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09714__A1 net103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09714__B2 net104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_181_3756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08874_ _04234_ _04242_ _04243_ _00824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_36_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07825_ _03557_ _03575_ _03577_ _00441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05736__C1 _01857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07756_ _03524_ _03532_ _03534_ _00415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05751__A2 _01934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_1022 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06707_ _02752_ _02846_ _02859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_67_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_79_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07687_ rf_ram.memory\[383\]\[1\] _03489_ _03492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_39_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09426_ _04588_ _01031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_66_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_149_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06638_ rf_ram.memory\[294\]\[0\] _02807_ _02808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_94_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05503__A2 _01687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07260__I _03017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_1313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09357_ net232 _04549_ _04540_ net233 _04550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_63_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06569_ _02738_ _02752_ _02753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_180_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_945 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08308_ _03309_ _02866_ _03878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08453__A1 _01418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_180_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09288_ net238 _04507_ _04508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_117_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_1288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output199_I net199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_43_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_172_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08239_ rf_ram.memory\[530\]\[1\] _03834_ _03836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_50_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05929__B _01923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11250_ _00986_ clknet_leaf_279_clk cpu.immdec.imm11_7\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_4
XANTENNA__09402__B1 _04564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10201_ _05078_ _05089_ _05090_ _01305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09953__A1 _04921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_1098 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11181_ _00917_ clknet_leaf_62_clk rf_ram.memory\[93\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_140_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output76_I net76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10132_ rf_ram.memory\[454\]\[0\] _05047_ _05048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_100_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08508__A2 net134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_1149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10063_ _03445_ _02866_ _05005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_89_2046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_89_2057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05990__A2 _02129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_1150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_3_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_159_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05742__A2 _01666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10079__A1 _02814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_67_1643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_187_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10965_ _00702_ clknet_leaf_9_clk rf_ram.memory\[171\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_67_1654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_1177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_167_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_1188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10896_ _00640_ clknet_leaf_13_clk rf_ram.memory\[182\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_100_2257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_1120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_1887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08444__A1 _02945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_980 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10251__A1 _02819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06455__B1 _01653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11517_ _01249_ clknet_leaf_200_clk rf_ram.memory\[34\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_124_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_151_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11448_ _01180_ clknet_leaf_240_clk cpu.state.init_done vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_33_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_170_Left_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10003__A1 _04950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09944__A1 _04911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08747__A2 _04152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_1273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11379_ _01111_ clknet_leaf_232_clk net124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_146_3106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_163_3420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05940_ _02133_ _02135_ _01563_ _02136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_179_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09172__A2 _04418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05871_ rf_ram.memory\[254\]\[0\] _01641_ _02004_ _02067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_124_2703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_192_clk_I clknet_5_30__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07183__A1 _03161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_1_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07610_ _03422_ _03442_ _03443_ _00360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_1_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08590_ rf_ram.memory\[167\]\[1\] _04064_ _04066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_89_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_178_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_3_4_0_clk clknet_0_clk clknet_3_4_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_88_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_72_clk_I clknet_5_8__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_1200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07541_ _03319_ _02904_ _03401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_117_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_1244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_186_560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07472_ rf_ram.memory\[366\]\[0\] _03357_ _03358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_53_1266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06143__C1 _01721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09211_ _04431_ _04451_ _04452_ _00952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06423_ _02606_ _02610_ _02614_ _02617_ _01660_ _02618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_45_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_146_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_146_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09142_ rf_ram.memory\[90\]\[0\] _04409_ _04410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06354_ rf_ram.memory\[236\]\[1\] _01614_ _01968_ rf_ram.memory\[237\]\[1\] _01959_
+ rf_ram.memory\[239\]\[1\] _02549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_127_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_173_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_161_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_130_clk_I clknet_5_24__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_173_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_296_clk clknet_5_7__leaf_clk clknet_leaf_296_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_05305_ _01500_ _01501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_72_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09073_ _04364_ _04365_ _04366_ _00900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_126_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_1015 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06285_ _01972_ _02478_ _02479_ _02480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__06997__A1 _03055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_1026 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_10_clk_I clknet_5_2__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08024_ _03690_ _03700_ _03702_ _00515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_170_983 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_135_2898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05236_ rf_ram_if.rdata1 _01435_ _01436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_141_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_1205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_130_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_102_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_1302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_25_1313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08738__A2 _01496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_145_clk_I clknet_5_26__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05167_ _01338_ _01344_ _01370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09975_ _02922_ _03253_ _04951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA_clkbuf_leaf_25_clk_I clknet_5_3__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08926_ _04266_ _04274_ _04275_ _00844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_157_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_157_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08857_ _04202_ _04231_ _04232_ _00818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05709__C1 _01656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07174__A1 _02894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07808_ _03554_ _03566_ _03567_ _00434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_leaf_220_clk clknet_5_22__leaf_clk clknet_leaf_220_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08788_ rf_ram.memory\[149\]\[0\] _04189_ _04190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05724__A2 _01856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06382__C1 _01925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07739_ _03359_ _03524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA_output114_I net114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05931__C _01978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10750_ _00494_ clknet_leaf_51_clk rf_ram.memory\[470\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08674__A1 _04094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_45_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_177_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09409_ _01436_ _01437_ _01344_ _01388_ _04579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_10681_ _00425_ clknet_leaf_80_clk rf_ram.memory\[437\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_165_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_62_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_137_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08426__A1 _03922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_980 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_1105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10233__A1 _05081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_287_clk clknet_5_18__leaf_clk clknet_leaf_287_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__06437__B1 _01609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08977__A2 _04303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_1115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05659__B _01783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_181_1310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11302_ _01035_ clknet_leaf_252_clk net67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_133_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11233_ _00969_ clknet_leaf_256_clk cpu.genblk3.csr.mcause31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07401__A2 _03083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11164_ _00900_ clknet_leaf_48_clk rf_ram.memory\[81\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_8_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10115_ _03071_ _03100_ _05037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_101_1024 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11095_ _00832_ clknet_leaf_84_clk rf_ram.memory\[127\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_41_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05963__A2 _01605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10046_ rf_ram.memory\[506\]\[1\] _04993_ _04995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_141_3014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_211_clk clknet_5_28__leaf_clk clknet_leaf_211_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08901__A2 _04257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_1108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_187_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_82_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_82_1927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10948_ _00686_ clknet_leaf_155_clk rf_ram.memory\[359\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_39_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05413__I _01513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_744 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_2_1215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10879_ _00623_ clknet_leaf_32_clk rf_ram.memory\[221\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_186_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06140__A2 _01719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_156_3290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09465__I0 net82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10224__A1 _03892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_278_clk clknet_5_17__leaf_clk clknet_leaf_278_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_108_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06979__A1 _02775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_117_2562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_117_2573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06070_ rf_ram.memory\[348\]\[1\] _01677_ _01678_ rf_ram.memory\[349\]\[1\] _01688_
+ rf_ram.memory\[351\]\[1\] _02265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XANTENNA_1 _02839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09917__A1 _04911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05403__A1 _01347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05254__I1 net105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09760_ _04818_ _01135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06972_ rf_ram.memory\[428\]\[1\] _03041_ _03043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08711_ _04126_ _04140_ _04141_ _00763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05923_ rf_ram.memory\[108\]\[0\] _01677_ _01702_ rf_ram.memory\[109\]\[0\] _01625_
+ rf_ram.memory\[111\]\[0\] _02119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_09691_ _04740_ net31 _04771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
Xclkbuf_leaf_202_clk clknet_5_25__leaf_clk clknet_leaf_202_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08642_ _02828_ _02881_ _04099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05854_ rf_ram.memory\[232\]\[0\] _01735_ _01956_ _02050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05706__A2 _01509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_156_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05751__C _01569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08573_ _02945_ _03945_ _04054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05785_ rf_ram.memory\[140\]\[0\] _01799_ _01931_ rf_ram.memory\[141\]\[0\] _01857_
+ rf_ram.memory\[143\]\[0\] _01981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_49_525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_89_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07524_ _03100_ _03390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__07459__A2 _03101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08656__A1 _04097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_1159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06116__C1 _01715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_176_3655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05323__I _01518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_176_3666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_130_1220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07455_ rf_ram.memory\[330\]\[0\] _03346_ _03347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_76_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_563 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_57_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06406_ _02597_ _02598_ _02599_ _02600_ _01670_ _02601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XTAP_TAPCELL_ROW_137_2938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_137_2949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_130_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_9_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07386_ rf_ram.memory\[24\]\[0\] _03303_ _03304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_106_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_134_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_269_clk clknet_5_16__leaf_clk clknet_leaf_269_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09125_ rf_ram.memory\[92\]\[0\] _04398_ _04399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_40_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06337_ rf_ram.memory\[220\]\[1\] _01755_ _01912_ rf_ram.memory\[221\]\[1\] _02019_
+ rf_ram.memory\[223\]\[1\] _02532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__08959__A2 _03945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09081__A1 _04367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09056_ rf_ram.memory\[101\]\[0\] _04355_ _04356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_163_1040 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06268_ rf_ram.memory\[158\]\[1\] _01501_ _02463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_102_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09908__A1 _04884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08007_ _03690_ _03687_ _03691_ _00509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_130_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05219_ cpu.decode.opcode\[2\] cpu.branch_op cpu.csr_d_sel _01419_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_25_1110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06199_ rf_ram.memory\[458\]\[1\] _01706_ _01650_ _02394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_12_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05926__C _01860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06198__A2 _01709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09958_ _04921_ _04938_ _04940_ _01212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05945__A2 _01536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06103__B _01620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09136__A2 _04067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08909_ _04234_ _04263_ _04264_ _00838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_86_2005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09889_ rf_ram.memory\[219\]\[1\] _04896_ _04898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_170_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06370__A2 _01683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10802_ _00546_ clknet_leaf_322_clk rf_ram.memory\[555\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08647__A1 net238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05233__I net134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_1136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10733_ _00477_ clknet_leaf_127_clk rf_ram.memory\[45\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_32_1147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_24_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10664_ _00408_ clknet_leaf_108_clk rf_ram.memory\[378\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_138_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10206__A1 _05078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05881__A1 _01972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10595_ _00339_ clknet_leaf_204_clk rf_ram.memory\[31\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_69_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_133_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_1210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_1146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_128_Right_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_11216_ _00952_ clknet_leaf_61_clk rf_ram.memory\[68\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_112_2470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_75_1786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_112_2481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_75_1797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06189__A2 _01782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput71 net71 o_dbus_adr[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput82 net82 o_dbus_adr[25] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput93 net93 o_dbus_adr[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_11147_ _00883_ clknet_leaf_68_clk rf_ram.memory\[107\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_128_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11078_ _00815_ clknet_leaf_15_clk rf_ram.memory\[133\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07138__A1 _03123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10029_ _04982_ _04983_ _04984_ _01239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08886__A1 _04237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_1074 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05571__C _01361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_1069 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06361__A2 _01515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_148_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_158_3330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08638__A1 _04094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05570_ _01754_ _01759_ _01349_ _01765_ _01766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_74_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07310__A1 _03225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_119_2602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06113__A2 _01644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_73_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_119_2613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07240_ _03193_ _03210_ _03212_ _00221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_129_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_154_3249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09438__I0 net69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_171_3563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07171_ _03157_ _03169_ _03170_ _00194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_171_3574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_147_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06122_ _02313_ _02314_ _02315_ _02316_ _01670_ _02317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_108_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_132_2846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_132_2857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05624__A1 _01675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06053_ rf_ram.memory\[364\]\[1\] _01644_ _01610_ rf_ram.memory\[365\]\[1\] _01636_
+ rf_ram.memory\[367\]\[1\] _02248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_169_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_112_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07377__A1 _03289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09812_ _02828_ _03035_ _04851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05318__I _01513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05927__A2 _01631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06955_ _03018_ _03029_ _03031_ _00117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09743_ _04804_ net17 _04807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__07129__A1 rf_ram.memory\[4\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05906_ _01768_ _02089_ _02101_ _01362_ _02102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_154_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09674_ _04757_ _01110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06886_ rf_ram.memory\[281\]\[0\] _02985_ _02986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_20_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08877__A1 net237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06337__C1 _02019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_178_3706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_1005 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08625_ _02821_ _02881_ _04088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05837_ _02021_ _02025_ _02029_ _02032_ _02033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__08629__A1 _04062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08556_ rf_ram.memory\[489\]\[1\] _04042_ _04044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05768_ rf_ram.memory\[145\]\[0\] _01664_ _01964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_07507_ _03360_ _03377_ _03379_ _00321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_92_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08487_ _03956_ _03995_ _03997_ _00683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05699_ rf_ram.memory\[414\]\[0\] _01543_ _01895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06104__A2 _01692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07438_ _03326_ _03334_ _03336_ _00295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_175_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07369_ _03292_ _03290_ _03293_ _00269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09054__A1 _04334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_162_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09108_ rf_ram.memory\[94\]\[0\] _04387_ _04388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_66_1243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10380_ _00124_ clknet_leaf_100_clk rf_ram.memory\[427\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_116_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09039_ _04334_ _04343_ _04345_ _00887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_60_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05937__B _01601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09409__B _01344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_57_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11001_ _00738_ clknet_leaf_270_clk rf_ram.memory\[519\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10134__I _02747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05918__A2 _01770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_70_1694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_29_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_1236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07540__A1 _03393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06343__A2 _01915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09293__A1 net237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_99_2229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_166_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_138_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10716_ _00460_ clknet_leaf_51_clk rf_ram.memory\[463\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_55_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10647_ _00391_ clknet_leaf_95_clk rf_ram.memory\[401\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09045__A1 _02828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_181_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_77_1826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_114_2510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10578_ _00322_ clknet_leaf_164_clk rf_ram.memory\[323\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_114_2521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_77_1837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_1218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09348__A2 _03991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_2_Left_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08020__A2 _03693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_1147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06582__A2 _02730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06740_ _02716_ _02793_ _02882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__08449__I net34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08859__A1 _04205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_64_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06671_ _02820_ _02833_ _02834_ _00030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07531__A1 _03319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06334__A2 _01940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08410_ _02761_ _03903_ _03942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_114_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05622_ rf_ram.memory\[494\]\[0\] _01543_ _01818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_149_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09390_ net217 _04561_ _04564_ net218 _04568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_47_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_173_3603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_148_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08341_ _03892_ _03009_ _03899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_173_3614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_157_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05553_ rf_ram.memory\[284\]\[0\] _01634_ _01678_ rf_ram.memory\[285\]\[0\] _01625_
+ rf_ram.memory\[287\]\[0\] _01749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_188_1124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_74_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_144_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08272_ _03855_ _03853_ _03856_ _00609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05484_ rf_ram.memory\[348\]\[0\] _01677_ _01678_ rf_ram.memory\[349\]\[0\] _01679_
+ rf_ram.memory\[351\]\[0\] _01680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XTAP_TAPCELL_ROW_15_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_1077 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07223_ _03190_ _03201_ _03202_ _00214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_85_1107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_132_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07154_ rf_ram.memory\[484\]\[0\] _03159_ _03160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08912__I _04057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07598__A1 net239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06105_ rf_ram.memory\[281\]\[1\] _01626_ _02300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_30_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07085_ rf_ram.memory\[491\]\[1\] _03114_ _03116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_113_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07528__I _03359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06270__A1 _01951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06036_ rf_ram.memory\[570\]\[1\] _01544_ _01540_ rf_ram.memory\[571\]\[1\] _01539_
+ rf_ram.memory\[569\]\[1\] _02231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XTAP_TAPCELL_ROW_188_3890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_160_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_35_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input38_I i_ibus_rdt[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07987_ rf_ram.memory\[467\]\[1\] _03676_ _03678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06938_ _03014_ _03020_ _03021_ _00110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09726_ _04795_ _01124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__05781__B1 _01608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06869_ _02970_ _02973_ _02974_ _00088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09657_ net98 net109 _04743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_96_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07522__A1 _03360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06325__A2 _01510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08608_ _02731_ _02939_ _04077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_78_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09588_ _02709_ _04699_ _04700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_78_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_139_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_1145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08539_ rf_ram.memory\[19\]\[1\] _04031_ _04033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_38_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08078__A2 _03729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11550_ _01282_ clknet_leaf_122_clk rf_ram.memory\[453\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_65_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_9_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05511__I _01503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05836__A1 _01972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10501_ _00245_ clknet_leaf_196_clk rf_ram.memory\[258\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_52_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11481_ _01213_ clknet_leaf_168_clk rf_ram.memory\[335\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_18_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_123_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_107_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_59_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10432_ _00176_ clknet_leaf_225_clk rf_ram.memory\[487\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_33_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_94_2137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_94_2148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_1062 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10363_ _00107_ clknet_leaf_179_clk rf_ram.memory\[278\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_131_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10294_ _00038_ clknet_leaf_269_clk rf_ram.memory\[523\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_29_Left_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_72_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_1213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_72_1745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07761__A1 _03524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07513__A1 _02775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_107_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_107_2391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09602__B _04526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_185_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_75_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_38_Left_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_69_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_185_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07816__A2 _03559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_987 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05421__I _01513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_151_3208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_153_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09018__A1 _02787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_153_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_55_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_840 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09569__A2 net52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_180_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_180_Right_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_clkbuf_5_5__f_clk_I clknet_3_1_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08241__A2 _03135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_1184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_47_Left_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_59_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_149_3159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07910_ _02822_ _03547_ _03630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08890_ rf_ram.memory\[479\]\[1\] _04251_ _04253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_166_3473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_166_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_166_3484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06004__A1 _01495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07841_ _03355_ _03587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__07752__A1 _02781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07772_ _03008_ _03496_ _03544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_127_2756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06723_ rf_ram.memory\[51\]\[0\] _02870_ _02871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09511_ _04637_ _04639_ _04641_ _01063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_177_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_56_Left_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_79_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09442_ net71 net72 _04593_ _04597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06654_ _02819_ _02820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_91_1188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_140_2989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05605_ _01661_ _01801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_177_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09373_ _04558_ _01008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06585_ _02761_ _02766_ _02767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_8_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_164_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08324_ _03887_ _03885_ _03888_ _00629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05536_ cpu.immdec.imm19_12_20\[6\] _01732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_75_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05331__I _01526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08255_ _03823_ _03843_ _03845_ _00603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_61_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09009__A1 _04298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05467_ rf_ram.memory\[374\]\[0\] _01662_ _01504_ _01663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_6_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08480__A2 _03992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_31_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07206_ rf_ram.memory\[262\]\[0\] _03191_ _03192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06491__A1 net252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08186_ _03787_ _03802_ _03803_ _00576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05398_ _01570_ _01593_ _01594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_104_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_42_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_65_Left_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07137_ rf_ram.memory\[498\]\[0\] _03148_ _03149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_63_1235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_186_3838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_186_3849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07068_ rf_ram.memory\[494\]\[0\] _03105_ _03106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09980__A2 _04951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05451__C1 _01646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07991__A1 _03651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06019_ rf_ram.memory\[552\]\[1\] _01524_ _01528_ _02214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_101_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_989 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_50_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_1039 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05506__I _01609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_74_Left_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09709_ _04783_ _01119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_173_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10981_ _00718_ clknet_leaf_0_clk rf_ram.memory\[167\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_69_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_1206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_139_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_136_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_26_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_25_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_147_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11533_ _01265_ clknet_leaf_192_clk rf_ram.memory\[351\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_68_1146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_151_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_83_Left_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_68_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_81_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_162_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11464_ _01196_ clknet_leaf_141_clk rf_ram.memory\[344\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_29_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_1302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10415_ _00159_ clknet_leaf_182_clk rf_ram.memory\[493\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11395_ _01127_ clknet_leaf_226_clk net110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_33_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10346_ _00090_ clknet_leaf_179_clk rf_ram.memory\[282\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_104_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10277_ _00021_ clknet_leaf_281_clk rf_ram.memory\[236\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05993__B1 _01950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09383__I _04539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07734__A1 _03491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_109_2420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_92_Left_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_109_2431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_144_3067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_1106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_144_3078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_178_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_161_3381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_161_3392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09487__A1 _02690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_17_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_122_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06170__B1 _01645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_146_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_1184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06370_ rf_ram.memory\[240\]\[1\] _01683_ _01684_ _02565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_139_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_185_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_1194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05321_ _01516_ _01517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_16_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_71_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_154_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08040_ net235 _03693_ _03712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_05252_ cpu.bne_or_bge _01452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_142_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_153_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05183_ _01380_ _01381_ _01382_ _01383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XTAP_TAPCELL_ROW_168_3513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10021__A2 _03009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09991_ _02727_ _02801_ _04961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_126_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07973__A1 _03668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08942_ rf_ram.memory\[122\]\[1\] _04283_ _04285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_86_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_181_3746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08873_ rf_ram.memory\[12\]\[0\] _04242_ _04243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_181_3757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07725__A1 _02795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07824_ rf_ram.memory\[433\]\[1\] _03575_ _03577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05736__B1 _01931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07755_ rf_ram.memory\[395\]\[1\] _03532_ _03534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09478__A1 _02703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06706_ _02826_ _02856_ _02858_ _00041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05770__B _01494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07686_ _03359_ _03491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_56_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08150__A1 _03757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_165_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06637_ _02801_ _02806_ _02807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09425_ net93 net94 _02707_ _04588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_133_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_137_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06568_ _02751_ _02752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_09356_ _03990_ _04549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_75_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08307_ _03855_ _03875_ _03877_ _00623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05519_ _01714_ _01715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_62_423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09287_ _04004_ _04507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_117_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06499_ _01375_ _02690_ _01400_ net132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_117_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05267__A2 _01418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08238_ _03820_ _03834_ _03835_ _00596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_90_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_62_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_105_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05672__C1 _01713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08169_ rf_ram.memory\[543\]\[0\] _03792_ _03793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_43_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10200_ rf_ram.memory\[191\]\[0\] _05089_ _05090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_28_1163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11180_ _00916_ clknet_leaf_61_clk rf_ram.memory\[93\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_113_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_313_clk_I clknet_5_5__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07964__A1 _03651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10131_ _02805_ _02832_ _05047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_24_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_max_cap238_I _02898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output69_I net69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10062_ _04985_ _05002_ _05004_ _01252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_175_1318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_89_2047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_89_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_328_clk_I clknet_5_4__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_3_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_187_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_1101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10079__A2 _02917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_1026 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_67_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08547__I _04037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10964_ _00701_ clknet_leaf_9_clk rf_ram.memory\[171\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08141__A1 net241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_1313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10895_ _00639_ clknet_leaf_17_clk rf_ram.memory\[181\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_128_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_167_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_100_2247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_100_2258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_913 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_26_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_80_1877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_80_1888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08444__A2 _03949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09641__A1 _04634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11516_ _01248_ clknet_leaf_144_clk rf_ram.memory\[306\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11447_ _01179_ clknet_leaf_240_clk cpu.state.stage_two_req vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_150_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_111_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06207__A1 _01350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09944__A2 _02923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11378_ _01110_ clknet_leaf_231_clk net123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_104_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05415__C1 _01610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_146_3107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10329_ _00073_ clknet_leaf_147_clk rf_ram.memory\[288\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_81_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_163_3421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07707__A1 _03488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05870_ _02062_ _02063_ _02064_ _02065_ _01620_ _02066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__05146__I _01348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_124_2704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08380__A1 _03134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_1_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07540_ _03393_ _03398_ _03400_ _00333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07471_ _02972_ _03101_ _03357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_147_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06143__B1 _01726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_146_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09880__A1 _04887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06422_ _01909_ _02615_ _02616_ _02617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_57_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09210_ rf_ram.memory\[68\]\[0\] _04451_ _04452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06694__A1 _02820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09141_ net245 _04005_ _04409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06353_ rf_ram.memory\[238\]\[1\] _01501_ _02548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_44_423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_139_2980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05304_ _01499_ _01500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_12
XFILLER_0_142_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09072_ rf_ram.memory\[81\]\[0\] _04365_ _04366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_114_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06284_ rf_ram.memory\[132\]\[1\] _01799_ _01912_ rf_ram.memory\[133\]\[1\] _01911_
+ rf_ram.memory\[135\]\[1\] _02479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XANTENNA__05749__C _01717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_1076 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06997__A2 _02899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08023_ rf_ram.memory\[571\]\[1\] _03700_ _03702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_170_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_142_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05235_ rf_ram_if.rtrig1 _01435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_135_2899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08199__A1 _03798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09396__B1 _04564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05166_ _01347_ _01369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_60_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07946__A1 _02728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09974_ _04396_ _04950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_08925_ rf_ram.memory\[124\]\[0\] _04274_ _04275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05709__B1 _01763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08856_ rf_ram.memory\[131\]\[0\] _04231_ _04232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input20_I i_dbus_rdt[26] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07174__A2 _03158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_1145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07807_ rf_ram.memory\[414\]\[0\] _03566_ _03567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_98_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05999_ rf_ram.memory\[518\]\[1\] _01502_ _01506_ _02194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08787_ _03071_ _04152_ _04189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06382__B1 _01912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07738_ _03521_ _03522_ _03523_ _00408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_67_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output107_I net107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07669_ rf_ram.memory\[403\]\[1\] _03478_ _03480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06134__B1 _01786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06685__A1 _02730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09408_ cpu.ctrl.i_jump _01426_ _04577_ _04578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_10680_ _00424_ clknet_leaf_80_clk rf_ram.memory\[437\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_36_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_165_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09339_ _04539_ _04540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__09623__A1 _04634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_109_Right_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_30_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_180_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_152_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_69_1252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_161_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_1322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11301_ _01034_ clknet_leaf_251_clk net96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_16_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_252_clk_I clknet_5_20__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11232_ _00968_ clknet_leaf_238_clk cpu.genblk3.csr.mstatus_mpie vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_121_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_31_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07937__A1 _03619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11163_ _00899_ clknet_leaf_35_clk rf_ram.memory\[0\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_105_1150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_8_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10114_ _05017_ _05034_ _05036_ _01272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06070__C1 _01688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11094_ _00831_ clknet_leaf_121_clk rf_ram.memory\[479\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_179_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_leaf_267_clk_I clknet_5_17__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_1182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10045_ _04982_ _04993_ _04994_ _01245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_141_3015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08362__A1 _03887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05176__A1 _01353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08114__A1 _03757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_82_1917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_82_1928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10947_ _00685_ clknet_leaf_149_clk rf_ram.memory\[369\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06676__A1 _02716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_1121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_151_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_128_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10878_ _00622_ clknet_leaf_32_clk rf_ram.memory\[221\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_205_clk_I clknet_5_24__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_13_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_156_3291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09465__I1 net83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10224__A2 _03134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05569__C _01670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_1216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06979__A2 _03040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_117_2563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_117_2574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_2 _02839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05651__A2 _01846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09917__A2 _03083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_1071 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05585__B _01746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05939__B1 _01607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06600__A1 _02743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05403__A2 _01346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05254__I2 net128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06971_ _03014_ _03041_ _03042_ _00122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_20_1211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_158_1313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08710_ rf_ram.memory\[151\]\[0\] _04140_ _04141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05922_ rf_ram.memory\[110\]\[0\] _01641_ _02004_ _02118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09690_ _04770_ _01113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_174_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08353__A1 _03008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08641_ _04097_ _04095_ _04098_ _00736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05853_ _01951_ _02047_ _02048_ _02049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_83_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_117_1032 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08572_ _04026_ _04051_ _04053_ _00712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05784_ rf_ram.memory\[142\]\[0\] _01770_ _01980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_107_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08105__A1 _03721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07523_ _03355_ _03389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__06116__B1 _01654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09853__A1 _02713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_1098 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_176_3656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_176_3667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07454_ _02775_ _02815_ _03346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06667__A1 _02736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09520__B _02709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_1105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06405_ rf_ram.memory\[82\]\[1\] _01652_ _01654_ rf_ram.memory\[83\]\[1\] _01656_
+ rf_ram.memory\[81\]\[1\] _02600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_146_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07385_ _02992_ _02997_ _03303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_137_2939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09605__A1 _04524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_44_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06336_ rf_ram.memory\[222\]\[1\] _01531_ _02531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09124_ _02838_ _04005_ _04398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_40_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05890__A2 _01510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_161_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07092__A1 _02915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09055_ _02794_ _04339_ _04355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_103_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06267_ _01373_ _02348_ _02461_ _02462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_170_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_995 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_163_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05218_ _01417_ _01418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_08006_ rf_ram.memory\[465\]\[1\] _03687_ _03691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_41_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06198_ rf_ram.memory\[460\]\[1\] _01709_ _01721_ rf_ram.memory\[461\]\[1\] _01713_
+ rf_ram.memory\[463\]\[1\] _02393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_124_1036 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07919__A1 _03622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05495__B _01629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05149_ rf_ram_if.rtrig0 _01352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_TAPCELL_ROW_5_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09957_ rf_ram.memory\[336\]\[1\] _04938_ _04940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_99_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08908_ rf_ram.memory\[125\]\[0\] _04263_ _04264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_86_2006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09888_ _04884_ _04896_ _04897_ _01185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_output224_I net224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05158__A1 _01353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08839_ _04205_ _04219_ _04221_ _00811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10151__A1 _05049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_1132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_169_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_1143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_36_1251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10801_ _00545_ clknet_leaf_322_clk rf_ram.memory\[556\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_95_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_184_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_135_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08647__A2 _04067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09844__A1 _02714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_1115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10732_ _00476_ clknet_leaf_127_clk rf_ram.memory\[45\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_27_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_24_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_24_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10663_ _00407_ clknet_leaf_94_clk rf_ram.memory\[397\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_180_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_91_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10594_ _00338_ clknet_leaf_204_clk rf_ram.memory\[31\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_106_631 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_191_clk_I clknet_5_28__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_3_3_0_clk clknet_0_clk clknet_3_3_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__05633__A2 _01735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_71_clk_I clknet_5_8__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_107_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11215_ _00951_ clknet_leaf_40_clk rf_ram.memory\[6\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_75_1787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_112_2471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_112_2482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_75_1798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput72 net72 o_dbus_adr[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput83 net83 o_dbus_adr[26] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__05397__A1 _01351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11146_ _00882_ clknet_leaf_68_clk rf_ram.memory\[107\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xoutput94 net94 o_dbus_adr[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA_clkbuf_leaf_86_clk_I clknet_5_10__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11077_ _00814_ clknet_leaf_15_clk rf_ram.memory\[133\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08335__A1 _03887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10028_ rf_ram.memory\[327\]\[0\] _04983_ _04984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10142__A1 _03672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_196_clk clknet_5_25__leaf_clk clknet_leaf_196_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08886__A2 _04248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06897__A1 _02958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05424__I _01493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_158_3320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_59_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_158_3331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_144_clk_I clknet_5_27__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_46_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_119_2603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_24_clk_I clknet_5_3__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_119_2614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09438__I1 net70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07170_ rf_ram.memory\[495\]\[0\] _03169_ _03170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_171_3564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05872__A2 _01677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_171_3575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_171_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_159_clk_I clknet_5_27__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06121_ rf_ram.memory\[258\]\[1\] _01500_ _01519_ rf_ram.memory\[259\]\[1\] _01668_
+ rf_ram.memory\[257\]\[1\] _02316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_26_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07074__A1 _03087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_171_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_147_1069 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_120_clk clknet_5_13__leaf_clk clknet_leaf_120_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_112_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_132_2847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_39_clk_I clknet_5_7__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06052_ rf_ram.memory\[366\]\[1\] _01631_ _02247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_23_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_78_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06204__B _01756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06034__C1 _01554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09811_ _04840_ _04848_ _04850_ _01154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_10_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_185_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09742_ _04806_ _01129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_94_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06954_ rf_ram.memory\[231\]\[1\] _03029_ _03031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_158_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_1131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05905_ _02092_ _02095_ _01660_ _02100_ _02101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__10133__A1 _05046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09673_ net123 _04736_ _04756_ _04757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06337__B1 _01912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06885_ _02958_ _02984_ _02985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__08877__A2 _04077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_187_clk clknet_5_28__leaf_clk clknet_leaf_187_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_178_3707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_171_1310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08624_ _04062_ _04085_ _04087_ _00730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_55_1137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05836_ _01972_ _02030_ _02031_ _02032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_90_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05334__I _01499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_89_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_166_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05767_ rf_ram.memory\[144\]\[0\] _01846_ _01956_ _01963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08555_ _04023_ _04042_ _04043_ _00705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_178_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_166_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09826__A1 _04840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07506_ rf_ram.memory\[363\]\[1\] _03377_ _03379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08486_ rf_ram.memory\[379\]\[1\] _03995_ _03997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05698_ _01882_ _01886_ _01890_ _01893_ _01894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_64_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07437_ rf_ram.memory\[332\]\[1\] _03334_ _03336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_21_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05312__A1 _01496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_1073 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_9_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_174_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_31_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05863__A2 _01940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_169_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07368_ rf_ram.memory\[251\]\[1\] _03290_ _03293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_91_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09107_ _02916_ _04005_ _04387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_116_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06319_ rf_ram.memory\[176\]\[1\] _01922_ _01923_ _02514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xclkbuf_leaf_111_clk clknet_5_15__leaf_clk clknet_leaf_111_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_32_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07299_ _03225_ _03247_ _03249_ _00243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_131_921 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_1255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_1266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06812__A1 _02930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_96_2190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09038_ rf_ram.memory\[105\]\[1\] _04343_ _04345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09409__C _01388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_57_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08565__A1 _04023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11000_ _00737_ clknet_leaf_270_clk rf_ram.memory\[519\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06025__C1 _01517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_1020 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09762__B1 _04760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06040__A2 _02234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08317__A1 _03855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_70_1695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10124__A1 _05017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_178_clk clknet_5_31__leaf_clk clknet_leaf_178_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_38_1313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_29_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09817__A1 net240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_185_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_36_1070 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_157_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_83_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_161_Right_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09293__A2 _04507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05839__C1 _01925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10715_ _00459_ clknet_leaf_88_clk rf_ram.memory\[408\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05303__A1 _01496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_165_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_165_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05854__A2 _01735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10646_ _00390_ clknet_leaf_95_clk rf_ram.memory\[401\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_64_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09045__A2 _04339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_107_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_102_clk clknet_5_15__leaf_clk clknet_leaf_102_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_134_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_114_2511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10577_ _00321_ clknet_5_27__leaf_clk rf_ram.memory\[363\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_77_1827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_140_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_77_1838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_114_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05606__A2 _01801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_1020 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06024__B _01528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05419__I _01550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09753__B1 _04760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_1104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06031__A2 _01544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11129_ _00865_ clknet_leaf_76_clk rf_ram.memory\[116\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08308__A1 _03309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_169_clk clknet_5_30__leaf_clk clknet_leaf_169_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__10115__A1 _03071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06670_ rf_ram.memory\[455\]\[0\] _02833_ _02834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_153_1040 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07531__A2 _02899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05621_ _01597_ _01731_ _01816_ _01817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_59_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05542__A1 _01675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_153_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_176_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05552_ rf_ram.memory\[286\]\[0\] _01543_ _01748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_8_1288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08340_ _03887_ _03896_ _03898_ _00635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_86_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_173_3604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_173_3615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_103_Left_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_50_1034 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06098__A2 _01687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_1176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08271_ rf_ram.memory\[197\]\[1\] _03853_ _03856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07295__A1 _02984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_188_1158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_157_884 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05483_ _01624_ _01679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_129_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05145__I1 _01346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_15_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07222_ rf_ram.memory\[425\]\[0\] _03201_ _03202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_15_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05845__A2 _01724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_172_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07153_ _02883_ _03158_ _03159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07598__A2 _03390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06104_ rf_ram.memory\[280\]\[1\] _01692_ _01684_ _02299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07084_ _03087_ _03114_ _03115_ _00162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_160_1022 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06035_ rf_ram.memory\[568\]\[1\] _01524_ _01528_ _02230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_188_3880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_188_3891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05329__I rf_ram.i_raddr\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_5_28__f_clk clknet_3_7_0_clk clknet_5_28__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_61_1174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_35_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_1136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_35_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_1196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06022__A2 _01502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07986_ _03651_ _03676_ _03677_ _00502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_52_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09725_ net106 _04790_ _04791_ net107 _04794_ _04795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__10106__A1 rf_ram.memory\[312\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06937_ rf_ram.memory\[228\]\[0\] _03020_ _03021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_5_22__f_clk_I clknet_3_5_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09656_ _03973_ _04736_ _04741_ _04742_ _01107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06868_ rf_ram.memory\[302\]\[0\] _02973_ _02974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08607_ _04062_ _04074_ _04076_ _00724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_179_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05819_ _01600_ _02009_ _02014_ _02015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_167_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05533__A1 _01349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09587_ _01469_ _04698_ _04699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06799_ rf_ram.memory\[50\]\[1\] _02924_ _02926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08538_ _04023_ _04031_ _04032_ _00699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_65_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_77_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06089__A2 _01719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08469_ _02714_ _03985_ _00677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xclkbuf_leaf_332_clk clknet_5_4__leaf_clk clknet_leaf_332_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_92_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10500_ _00244_ clknet_leaf_196_clk rf_ram.memory\[258\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_162_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11480_ _01212_ clknet_leaf_177_clk rf_ram.memory\[336\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_33_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07038__A1 _03050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_59_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10431_ _00175_ clknet_leaf_224_clk rf_ram.memory\[500\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_94_2138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_94_2149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08786__A1 _04170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06623__I _02794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output99_I net99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10362_ _00106_ clknet_leaf_179_clk rf_ram.memory\[278\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_33_598 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_60_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06261__A2 _01801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10293_ _00037_ clknet_leaf_269_clk rf_ram.memory\[524\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_131_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_103_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08538__A1 _04023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_72_1735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_72_1746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_1247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06013__A2 _01544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07210__A1 _03193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_1132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_16_Right_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_77_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07513__A2 _03101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_107_2381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_150_1202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_69_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_107_2392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_150_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_157_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_173_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07277__A1 _03222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_323_clk clknet_5_4__leaf_clk clknet_leaf_323_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_83_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06019__B _01528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_12_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05827__A2 _01515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06485__C1 _01635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_181_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09018__A2 _04303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07029__A1 _02738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10629_ _00373_ clknet_leaf_92_clk rf_ram.memory\[387\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05858__B _01956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_25_Right_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_144_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07629__I _03355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08777__A1 _02971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_1114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_1163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_121_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_166_3474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_166_3485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07201__A1 _03157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07840_ _03557_ _03584_ _03586_ _00447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07771_ _03524_ _03541_ _03543_ _00421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_127_2757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_34_Right_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09510_ rf_ram.memory\[279\]\[1\] _04639_ _04641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06201__C _01658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06722_ _02866_ _02869_ _02870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_182_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08701__A1 _04126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09441_ _04596_ _01038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06653_ _02742_ _02819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XPHY_EDGE_ROW_111_Left_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__11614__I net94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05604_ rf_ram.memory\[304\]\[0\] _01799_ _01602_ _01800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09372_ net208 _04549_ _04552_ net209 _04558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09257__A2 _01484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06584_ _02765_ _02766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_46_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05612__I _01640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_176_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08323_ rf_ram.memory\[242\]\[1\] _03885_ _03888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_75_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05535_ _01368_ _01673_ _01730_ _01731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_117_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_314_clk clknet_5_5__leaf_clk clknet_leaf_314_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_74_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06476__C1 _01607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08254_ rf_ram.memory\[527\]\[1\] _03843_ _03845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05466_ _01661_ _01662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_90_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_43_Right_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08480__A3 _01418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_31_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_31_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07205_ _02806_ _02941_ _03191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_144_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08185_ rf_ram.memory\[540\]\[0\] _03802_ _03803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05397_ _01351_ _01581_ _01592_ _01362_ _01593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_166_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07136_ _02915_ _02923_ _03148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_127_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_186_3839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06243__A2 _01856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_1209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07067_ _02915_ _02972_ _03105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA_input50_I i_ibus_rdt[25] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_54_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05451__B1 _01645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06018_ rf_ram.memory\[556\]\[1\] _01511_ _01517_ rf_ram.memory\[557\]\[1\] _01521_
+ rf_ram.memory\[559\]\[1\] _02213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XANTENNA__09193__A1 _04434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_50_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07274__I _03039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_52_Right_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06400__C1 _01810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1018 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output137_I net137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07969_ _03651_ _03665_ _03666_ _00496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05754__A1 _01373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09708_ net101 _04767_ _04768_ net102 _04782_ _04783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_0_69_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10980_ _00717_ clknet_leaf_339_clk rf_ram.memory\[167\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09496__A2 _01388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09639_ _02971_ _04507_ _04728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_139_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_139_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07259__A1 _03222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_305_clk clknet_5_4__leaf_clk clknet_leaf_305_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_167_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_61_Right_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_154_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_843 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11532_ _01264_ clknet_leaf_144_clk rf_ram.memory\[310\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_53_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05809__A2 _01641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05678__B _01756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11463_ _01195_ clknet_leaf_192_clk rf_ram.memory\[344\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_80_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06482__A2 _01643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08759__A1 _01363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10414_ _00158_ clknet_leaf_183_clk rf_ram.memory\[493\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_123_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_1314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05397__C _01362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11394_ _01126_ clknet_leaf_226_clk net108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_60_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07431__A1 _03323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06234__A2 _01500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10345_ _00089_ clknet_leaf_136_clk rf_ram.memory\[302\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_104_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10276_ _00020_ clknet_leaf_281_clk rf_ram.memory\[236\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05993__A1 _01371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_70_Right_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09184__A1 net242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_5_11__f_clk clknet_3_2_0_clk clknet_5_11__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_40_1055 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_109_2421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08931__A1 _04266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1099 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_144_3068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_144_3079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_161_3382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_161_3393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07498__A1 _03319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_17_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_122_2654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_159_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_122_2665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_159_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_152_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_28_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_51_1162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_1293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_173_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05320_ _01515_ _01516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__06458__C1 _01518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_142_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05251_ _01381_ _01450_ _01451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07670__A1 _03458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05588__B _01783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06473__A2 _01686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_181_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05182_ cpu.decode.opcode\[0\] _01382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_0_141_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_168_3514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06225__A2 _01631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09990_ _04953_ _04958_ _04960_ _01224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_110_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07973__A2 _02972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08941_ _04266_ _04283_ _04284_ _00850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05984__A1 rf_ram.memory\[0\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11609__I net87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_1310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_32_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08872_ _02787_ _03945_ _04242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_181_3747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_1275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_181_3758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07725__A2 _02869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07823_ _03554_ _03575_ _03576_ _00440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07754_ _03521_ _03532_ _03533_ _00414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06705_ rf_ram.memory\[522\]\[1\] _02856_ _02858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07685_ _03488_ _03489_ _03490_ _00388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_leaf_91_clk clknet_5_11__leaf_clk clknet_leaf_91_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09424_ _04587_ _01030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_56_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06636_ _02805_ _02806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_94_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05342__I _01537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09355_ _04548_ _01000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_47_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_158_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06567_ _02750_ _02726_ _02751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__08989__A1 _04298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08306_ rf_ram.memory\[221\]\[1\] _03875_ _03877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11507__CLK clknet_5_30__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05518_ _01513_ _01714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_90_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09286_ _04506_ _00973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_35_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06498_ _02690_ _02691_ _01400_ net133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_7_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_173_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07661__A1 net238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05498__B _01693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08237_ rf_ram.memory\[530\]\[0\] _03834_ _03835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_43_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06464__A2 _01536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05449_ _01609_ _01645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_12
XFILLER_0_172_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05672__B1 _01721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08168_ _02881_ _02909_ _03792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_31_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07119_ rf_ram.memory\[500\]\[1\] _03136_ _03138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_105_1310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08099_ rf_ram.memory\[556\]\[0\] _03748_ _03749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_24_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10130_ _02742_ _05046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_30_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05975__A1 _01903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_1129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09166__A1 _04401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10061_ rf_ram.memory\[507\]\[1\] _05002_ _05004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08913__A1 _03039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05517__I _01653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_89_2048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_89_2059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_159_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05680__C _01717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10963_ _00700_ clknet_leaf_288_clk rf_ram.memory\[19\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_98_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_67_1645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_1173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_82_clk clknet_5_11__leaf_clk clknet_leaf_82_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08141__A2 _03765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06152__A1 net252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_183_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10894_ _00638_ clknet_leaf_15_clk rf_ram.memory\[181\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_85_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_100_2248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_167_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05360__C1 _01555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_100_2259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_183_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_26_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_1878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_170_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_80_1889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_164_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11515_ _01247_ clknet_leaf_165_clk rf_ram.memory\[306\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_108_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06455__A2 _01661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_135_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05663__B1 _01857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11446_ _01178_ clknet_leaf_289_clk rf_ram.memory\[60\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_46_1231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06016__C _01569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_145_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11377_ _01109_ clknet_leaf_231_clk net120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_150_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05415__B1 _01608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_146_3108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10328_ _00072_ clknet_leaf_136_clk rf_ram.memory\[288\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09157__A1 _02991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_163_3422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10259_ _02916_ _03692_ _05125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05427__I _01605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08904__A1 _04234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05718__A1 _01909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_124_2705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08380__A2 _03903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05871__B _02004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_73_clk clknet_5_10__leaf_clk clknet_leaf_73_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_88_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07470_ _03355_ _03356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_159_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06421_ rf_ram.memory\[124\]\[1\] _01799_ _01772_ rf_ram.memory\[125\]\[1\] _01786_
+ rf_ram.memory\[127\]\[1\] _02616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_146_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_173_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_56_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_118_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09140_ _04401_ _04406_ _04408_ _00925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_57_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06352_ _01674_ _02534_ _02546_ _01362_ _02547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XTAP_TAPCELL_ROW_139_2970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_139_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05303_ _01496_ _01498_ _01499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_72_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07643__A1 _03455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06283_ rf_ram.memory\[134\]\[1\] _01531_ _02478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09071_ net248 _04005_ _04365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_170_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_4_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_1066 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08022_ _03686_ _03700_ _03701_ _00514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05234_ _01432_ _01418_ _01420_ _01433_ _01434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_71_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_1099 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08199__A2 _02984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05165_ _01353_ cpu.immdec.imm19_12_20\[6\] _01367_ cpu.immdec.imm24_20\[2\] _01368_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_123_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07946__A2 _02832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09973_ _04921_ _04947_ _04949_ _01218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09148__A1 _04397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08924_ _02838_ _04038_ _04274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_41_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08855_ net240 _04195_ _04231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_157_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07806_ _02916_ _03559_ _03566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_2_Right_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08786_ _04170_ _04186_ _04188_ _00791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_58_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05998_ _02189_ _02190_ _02191_ _02192_ _02193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_93_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input13_I i_dbus_rdt[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07737_ rf_ram.memory\[378\]\[0\] _03522_ _03523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_49_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_170_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_79_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_64_clk clknet_5_8__leaf_clk clknet_leaf_64_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07668_ _03455_ _03478_ _03479_ _00382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_177_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_45_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09407_ cpu.ctrl.i_jump _01472_ _01344_ _04577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06619_ _02748_ _02789_ _02791_ _00021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07882__A1 _03590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07599_ rf_ram.memory\[354\]\[0\] _03436_ _03437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_153_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09338_ net65 _02696_ _04539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_36_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06437__A2 _01633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09269_ cpu.genblk3.csr.o_new_irq _04493_ _04494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_133_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_23_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_563 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06117__B _01629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11300_ _01033_ clknet_leaf_251_clk net95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_65_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_max_cap250_I _02727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11231_ _00967_ clknet_leaf_239_clk cpu.genblk3.csr.mie_mtie vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_output81_I net81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11162_ _00898_ clknet_leaf_35_clk rf_ram.memory\[0\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_101_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05675__C _01658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10113_ rf_ram.memory\[392\]\[1\] _05034_ _05036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06070__B1 _01678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_1184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11093_ _00830_ clknet_leaf_121_clk rf_ram.memory\[479\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_175_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10044_ rf_ram.memory\[506\]\[0\] _04993_ _04994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_141_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05691__B _01783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_1268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_55_clk clknet_5_9__leaf_clk clknet_leaf_55_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_39_1090 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_82_1918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10946_ _00684_ clknet_leaf_149_clk rf_ram.memory\[369\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_82_1929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10577__CLK clknet_5_27__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07873__A1 _02836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10877_ _00621_ clknet_leaf_214_clk rf_ram.memory\[244\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_128_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05884__B1 _01925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_183_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_156_3292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_738 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_164_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_1228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_117_2564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_117_2575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_3 _03009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11429_ _01161_ clknet_leaf_291_clk rf_ram.memory\[62\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05866__B _02004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_46_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_5_9__f_clk clknet_3_2_0_clk clknet_5_9__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08050__A1 _03071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06970_ rf_ram.memory\[428\]\[0\] _03041_ _03042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05254__I3 net114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_184_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_input5_I i_dbus_rdt[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_1223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05921_ _02105_ _02109_ _02113_ _02116_ _01660_ _02117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XANTENNA__09550__A1 _01391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08353__A2 _03903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08640_ rf_ram.memory\[162\]\[1\] _04095_ _04098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_179_805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_175_Right_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05852_ rf_ram.memory\[236\]\[0\] _01614_ _01968_ rf_ram.memory\[237\]\[0\] _01959_
+ rf_ram.memory\[239\]\[0\] _02048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XANTENNA__05167__A2 _01344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08571_ rf_ram.memory\[170\]\[1\] _04051_ _04053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05783_ _01976_ _01977_ _01978_ _01979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_53_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_46_clk clknet_5_12__leaf_clk clknet_leaf_46_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09302__A1 _04466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07522_ _03360_ _03386_ _03388_ _00327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_18_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_1005 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_1174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_176_3657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_312_clk_I clknet_5_5__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_176_3668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07453_ _03326_ _03343_ _03345_ _00301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06667__A2 _02830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_186_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11622__I net72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06404_ rf_ram.memory\[80\]\[1\] _01863_ _01602_ _02599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_29_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_174_565 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07384_ _03292_ _03300_ _03302_ _00275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_17_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09605__A2 net49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09123_ _04396_ _04397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_128_993 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07616__A1 _03422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_1318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06335_ _02527_ _02529_ _01928_ _02530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_72_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_327_clk_I clknet_5_4__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05627__B1 _01688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09054_ _04334_ _04352_ _04354_ _00893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07092__A2 _03009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06266_ _01372_ _02404_ _02460_ _02461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_115_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08005_ _03689_ _03690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_05217_ cpu.state.cnt_r\[3\] cpu.mem_bytecnt\[1\] _01385_ cpu.state.o_cnt\[2\] _01417_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_13_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_1173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06197_ rf_ram.memory\[462\]\[1\] _01719_ _01707_ _02392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xmax_cap250 _02727_ net250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_64_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05148_ _01350_ _01351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_09956_ _04918_ _04938_ _04939_ _01211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_5_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08907_ _02959_ _04038_ _04263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09887_ rf_ram.memory\[219\]\[0\] _04896_ _04897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_99_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08838_ rf_ram.memory\[469\]\[1\] _04219_ _04221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_142_Right_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06355__A1 _01951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_1100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_135_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08769_ _04167_ _04177_ _04178_ _00784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_170_1024 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_leaf_37_clk clknet_5_7__leaf_clk clknet_leaf_37_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10800_ _00544_ clknet_leaf_322_clk rf_ram.memory\[556\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_95_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_178_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_1285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10731_ _00475_ clknet_leaf_55_clk rf_ram.memory\[443\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07855__A1 _03587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_24_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10662_ _00406_ clknet_leaf_93_clk rf_ram.memory\[397\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06626__I cpu.immdec.imm11_7\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_180_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05530__I _01635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07607__A1 _03425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10593_ _00337_ clknet_leaf_203_clk rf_ram.memory\[35\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_149_Left_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08280__A1 _03852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_133_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11214_ _00950_ clknet_leaf_40_clk rf_ram.memory\[6\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08032__A1 _03686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_112_2472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_75_1788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_75_1799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09780__A1 net244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_112_2483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput73 net73 o_dbus_adr[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_11145_ _00881_ clknet_leaf_71_clk rf_ram.memory\[108\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xoutput84 net84 o_dbus_adr[27] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_101_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06594__A1 _02748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05397__A2 _01581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput95 net95 o_dbus_adr[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_11076_ _00813_ clknet_leaf_25_clk rf_ram.memory\[134\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_158_Left_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10027_ _04911_ _02829_ _04983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10142__A2 _02883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06897__A2 _02992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_28_clk clknet_5_3__leaf_clk clknet_leaf_28_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_58_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_158_3321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_158_3332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_188_1318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10929_ _00673_ clknet_leaf_7_clk rf_ram.memory\[175\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_129_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_184_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_119_2604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_160_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_67_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_119_2615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05440__I _01635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_167_Left_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_27_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_1069 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_171_3565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_171_3576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06120_ rf_ram.memory\[256\]\[1\] _01644_ _01526_ _02315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_81_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_152_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_950 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06051_ _02243_ _02245_ _01629_ _02246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_132_2848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07367__I _03017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_99_Right_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06034__B1 _01555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09810_ rf_ram.memory\[74\]\[1\] _04848_ _04850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_10_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05388__A2 _01511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06585__A1 _02761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_176_Left_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09741_ net112 _04790_ _04791_ net113 _04805_ _04806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_06953_ _03014_ _03029_ _03030_ _00116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11617__I net67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09523__A1 _03992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_1110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05904_ _02096_ _02097_ _02098_ _02099_ _01670_ _02100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_09672_ _04754_ _04755_ _04735_ _04756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_59_1241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06884_ _02983_ _02984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__06220__B _01790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05615__I _01635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_178_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08623_ rf_ram.memory\[529\]\[1\] _04085_ _04087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_178_3708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05835_ rf_ram.memory\[220\]\[0\] _01755_ _01968_ rf_ram.memory\[221\]\[0\] _02019_
+ rf_ram.memory\[223\]\[0\] _02031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_0_171_1322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_1296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_19_clk clknet_5_2__leaf_clk clknet_leaf_19_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA_clkbuf_leaf_251_clk_I clknet_5_20__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08554_ rf_ram.memory\[489\]\[0\] _04042_ _04043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05766_ _01957_ _01961_ _01564_ _01962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07505_ _03356_ _03377_ _03378_ _00320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_76_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08485_ _03953_ _03995_ _03996_ _00682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_147_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_37_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05697_ _01675_ _01891_ _01892_ _01893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_65_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_185_Left_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07436_ _03323_ _03334_ _03335_ _00294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_18_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_21_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_73_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_174_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_266_clk_I clknet_5_17__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07367_ _03017_ _03292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_134_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09106_ _04367_ _04384_ _04386_ _00913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_72_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06318_ rf_ram.memory\[180\]\[1\] _01711_ _01772_ rf_ram.memory\[181\]\[1\] _01773_
+ rf_ram.memory\[183\]\[1\] _02513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_131_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07298_ rf_ram.memory\[25\]\[1\] _03247_ _03249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_96_2180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06273__B1 _01959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_96_2191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09037_ _04331_ _04343_ _04344_ _00886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06249_ rf_ram.memory\[446\]\[1\] _01531_ _02444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_103_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08014__A1 _03690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_57_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_57_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_92_2099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06025__B1 _01521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09762__A1 net119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_1121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06576__A1 _02756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_102_1143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_204_clk_I clknet_5_24__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09939_ _02868_ _02899_ _04929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_70_1696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05525__I _01714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_219_clk_I clknet_5_22__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_185_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09817__A2 _03253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07828__A1 _03554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_95_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05839__B1 _01912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10714_ _00458_ clknet_leaf_89_clk rf_ram.memory\[408\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_166_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_181_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06500__A1 _01376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_1313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10645_ _00389_ clknet_leaf_107_clk rf_ram.memory\[383\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_153_3240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_563 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_181_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08253__A1 _03820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10576_ _00320_ clknet_leaf_159_clk rf_ram.memory\[363\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_180_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_2_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_12_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_114_2512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_77_1828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_114_2523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_77_1839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10060__A1 _04982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09753__A1 net116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_1075 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06567__A1 _02750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11128_ _00864_ clknet_leaf_76_clk rf_ram.memory\[116\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_78_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_1127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08308__A2 _02866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11059_ _00796_ clknet_leaf_12_clk rf_ram.memory\[140\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10115__A2 _03100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05435__I _01530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_188_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_87_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05620_ net252 _01767_ _01815_ _01816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_118_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_8_1245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_153_1074 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_147_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05551_ _01743_ _01745_ _01746_ _01747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_80_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_173_3605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08270_ _03689_ _03855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__08492__A1 _03956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05482_ _01617_ _01678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__07295__A2 _02997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_184_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07221_ _02752_ _03040_ _03201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_15_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_73_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_156_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_1109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_172_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07152_ _02910_ _03158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_15_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06103_ _02295_ _02297_ _01620_ _02298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_113_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07083_ rf_ram.memory\[491\]\[0\] _03114_ _03115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_8_clk clknet_5_0__leaf_clk clknet_leaf_8_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_42_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07097__I _03013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06034_ rf_ram.memory\[572\]\[1\] _01538_ _01555_ rf_ram.memory\[573\]\[1\] _01554_
+ rf_ram.memory\[575\]\[1\] _02229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_125_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_188_3881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_188_3892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_1142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_1284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09744__B2 net114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_35_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_35_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07985_ rf_ram.memory\[467\]\[0\] _03676_ _03677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_52_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09724_ _04781_ net10 _04794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_06936_ _02766_ _02883_ _03020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05781__A2 _01606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09655_ net1 net2 _04736_ _04742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06867_ _02935_ _02972_ _02973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_190_clk_I clknet_5_28__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08606_ rf_ram.memory\[164\]\[1\] _04074_ _04076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05818_ _02010_ _02011_ _02012_ _02013_ _01978_ _02014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
Xclkbuf_3_2_0_clk clknet_0_clk clknet_3_2_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_09586_ net134 _01339_ _04698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06730__A1 _02873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06798_ _02873_ _02924_ _02925_ _00066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_leaf_70_clk_I clknet_5_8__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08537_ rf_ram.memory\[19\]\[0\] _04031_ _04032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_77_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05749_ _01941_ _01942_ _01943_ _01944_ _01717_ _01945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_148_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_148_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08483__A1 net244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08468_ _03968_ _03969_ _03984_ _03985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_33_1277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_18_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_98_2220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07419_ rf_ram.memory\[371\]\[0\] _03324_ _03325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_46_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_85_clk_I clknet_5_10__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08399_ _03922_ _03933_ _03935_ _00657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_163_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10430_ _00174_ clknet_leaf_224_clk rf_ram.memory\[500\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08235__A1 _03823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_59_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_162_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_94_2139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10042__A1 _04985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09983__A1 _04950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10361_ _00105_ clknet_leaf_138_clk rf_ram.memory\[298\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_61_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_1075 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10292_ _00036_ clknet_leaf_269_clk rf_ram.memory\[524\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_104_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_72_1736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_143_clk_I clknet_5_27__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07735__I _03355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_23_clk_I clknet_5_3__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_158_clk_I clknet_5_27__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_107_2382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_38_clk_I clknet_5_7__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05524__A2 _01719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_107_2393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07470__I _03355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_186_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_111_1209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_83_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_95_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_28_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_138_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06485__B1 _01714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_12_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_187_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10628_ _00372_ clknet_leaf_92_clk rf_ram.memory\[387\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08226__A1 _03798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07029__A2 _02992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_1105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_181_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10033__A1 _02805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08777__A2 _04152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10559_ _00303_ clknet_leaf_158_clk rf_ram.memory\[330\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_161_1310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06788__A1 _02915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06035__B _01528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_110_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_121_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_166_3475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_166_3486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05748__C1 _01645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05212__A1 _01375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07770_ rf_ram.memory\[393\]\[1\] _03541_ _03543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_127_2747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06960__A1 _03018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_127_2758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_159_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06721_ _02868_ _02869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_91_1102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_78_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_188_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09440_ net70 net71 _04593_ _04596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06652_ _02748_ _02816_ _02818_ _00027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06173__C1 _01715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06712__A1 _02728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05603_ _01613_ _01799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_09371_ _04557_ _01007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_59_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06583_ _02731_ _02764_ _02765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_75_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_176_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_923 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08322_ _03689_ _03887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_86_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05534_ _01674_ _01705_ _01729_ _01361_ _01730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_46_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05279__A1 _01366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06476__B1 _01609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08253_ _03820_ _03843_ _03844_ _00602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_46_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05465_ _01499_ _01661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_62_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11630__I net80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07204_ _03013_ _03190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__08217__A1 _03820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_31_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08184_ _02838_ _02846_ _03802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_31_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_43_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05396_ _01586_ _01591_ _01351_ _01592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_132_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07135_ _03126_ _03145_ _03147_ _00181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_63_1215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_1226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_113_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07066_ _03092_ _03102_ _03104_ _00155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xoutput230 net230 o_ibus_adr[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_63_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_54_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06017_ rf_ram.memory\[558\]\[1\] _01502_ _01506_ _02212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09717__A1 net104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09717__B2 net105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_1070 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input43_I i_ibus_rdt[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_250_clk clknet_5_20__leaf_clk clknet_leaf_250_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__06400__B1 _01646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07968_ rf_ram.memory\[47\]\[0\] _03665_ _03666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06951__A1 _02766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05754__A2 _01817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06919_ _02785_ _02758_ _03007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_09707_ _04781_ net5 _04782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_07899_ _03622_ _03620_ _03623_ _00469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09638_ _04524_ _01391_ _04727_ _01104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_69_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_1208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_168_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09569_ _04478_ net52 _04678_ _04684_ _04685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_183_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11600_ _01330_ clknet_leaf_306_clk rf_ram.memory\[574\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_167_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_176_980 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_154_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_136_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_102_2290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_1220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11531_ _01263_ clknet_leaf_145_clk rf_ram.memory\[310\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10263__A1 _02825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_184_1321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_163_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11462_ _01194_ clknet_leaf_139_clk rf_ram.memory\[292\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08208__A1 _03790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06219__B1 _01786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10015__A1 _04953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09956__A1 _04918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08759__A2 _01366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10413_ _00157_ clknet_leaf_182_clk rf_ram.memory\[494\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_123_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_116_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11393_ _01125_ clknet_leaf_225_clk net107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_104_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10344_ _00088_ clknet_leaf_136_clk rf_ram.memory\[302\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_103_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05978__C1 _01653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05442__A1 _01527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09708__A1 net101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05694__B _01790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10275_ _00019_ clknet_leaf_278_clk rf_ram.memory\[235\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_148_3150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05993__A2 _01594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09184__A2 _04067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_241_clk clknet_5_21__leaf_clk clknet_leaf_241_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_109_2422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_144_3069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05745__A2 _01940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_161_3383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_159_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07498__A2 _02883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06155__C1 _01679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_17_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05713__I _01756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_186_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_122_2655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_1131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_122_2666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_1204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_158_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06170__A2 _01644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_1237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_1248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_185_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_173_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06458__B1 _01655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10254__A1 net249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_142_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05250_ _01399_ _01382_ _01450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_126_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05681__A1 _01350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05181_ cpu.branch_op _01381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_101_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_168_3515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08940_ rf_ram.memory\[122\]\[0\] _04283_ _04284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05984__A2 _01613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08871_ _04237_ _04239_ _04241_ _00823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_86_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_32_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07186__A1 _03157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_181_3748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_181_3759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07822_ rf_ram.memory\[433\]\[0\] _03575_ _03576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_232_clk clknet_5_23__leaf_clk clknet_leaf_232_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__05736__A2 _01799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07753_ rf_ram.memory\[395\]\[0\] _03532_ _03533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11625__I net75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06704_ _02820_ _02856_ _02857_ _00040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06146__C1 _01726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07684_ rf_ram.memory\[383\]\[0\] _03489_ _03490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08686__A1 _04097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09423_ net92 net93 _02707_ _04587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06635_ _02773_ _02793_ _02805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_177_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06161__A2 _01692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09354_ net231 _03991_ _04540_ net232 _04548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_59_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06566_ _01496_ _01497_ _02750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XTAP_TAPCELL_ROW_47_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08438__A1 _03956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_980 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08305_ _03852_ _03875_ _03876_ _00622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_164_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_299_clk clknet_5_7__leaf_clk clknet_leaf_299_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_05517_ _01653_ _01713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_09285_ cpu.genblk3.csr.mcause3_0\[3\] _04505_ _04497_ _04506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_7_530 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06497_ cpu.bne_or_bge _01375_ _02691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_173_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08236_ _03798_ _02923_ _03834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_173_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05448_ _01643_ _01644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_62_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07661__A2 _03089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09938__A1 _04921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08167_ _03790_ _03788_ _03791_ _00569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_166_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_160_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05379_ _01571_ _01572_ _01573_ _01574_ _01575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_67_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07118_ _03123_ _03136_ _03137_ _00174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08098_ _02787_ _03729_ _03748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08610__A1 net238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07049_ _03092_ _03090_ _03093_ _00149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_28_1198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_100_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10060_ _04982_ _05002_ _05003_ _01251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06122__C _01670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_223_clk clknet_5_29__leaf_clk clknet_leaf_223_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08913__A2 _03083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_89_2049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06924__A1 _02970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_173_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05961__C _01568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_3_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06629__I _02800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08677__A1 _02953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10962_ _00699_ clknet_leaf_283_clk rf_ram.memory\[19\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06137__C1 _01793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_67_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_104_2330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10893_ _00637_ clknet_leaf_30_clk rf_ram.memory\[214\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_84_1960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05360__B1 _01554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_100_2249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10236__A1 _02819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_80_1879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_130_Left_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_164_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11514_ _01246_ clknet_leaf_197_clk rf_ram.memory\[506\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_135_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_184_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_1102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09929__A1 _04911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11445_ _01177_ clknet_leaf_290_clk rf_ram.memory\[60\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_1270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11376_ _01108_ clknet_leaf_230_clk net109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_22_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_156_Right_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10327_ _00071_ clknet_leaf_122_clk rf_ram.memory\[290\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_146_3109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05966__A2 _01514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09157__A2 _04418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10258_ _02825_ _05122_ _05124_ _01328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_163_3423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07168__A1 _03161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06032__C _01494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_214_clk clknet_5_19__leaf_clk clknet_leaf_214_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_56_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10189_ _02765_ _02972_ _05083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06376__C1 _01696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_124_2706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_159_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06143__A2 _01652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07340__A1 _03257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06420_ rf_ram.memory\[126\]\[1\] _01770_ _02615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_53_1269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06351_ _02537_ _02540_ _01350_ _02545_ _02546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_127_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_139_2971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05302_ _01497_ _01498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_4
XTAP_TAPCELL_ROW_139_2982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09070_ _04057_ _04364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_06282_ _02465_ _02469_ _02473_ _02476_ _02477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_72_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08840__A1 _02805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08021_ rf_ram.memory\[571\]\[0\] _03700_ _03701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_60_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05654__A1 _01769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05233_ net134 _01433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_53_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_170_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05164_ _01363_ _01366_ _01357_ _01367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_141_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_1229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_123_Right_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09972_ rf_ram.memory\[464\]\[1\] _04947_ _04949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05957__A2 _01633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08923_ _04269_ _04271_ _04273_ _00843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07159__A1 _02915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_205_clk clknet_5_24__leaf_clk clknet_leaf_205_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08854_ _04205_ _04228_ _04230_ _00817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05709__A2 _01500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06906__A1 _02970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_97_1174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07805_ _03557_ _03563_ _03565_ _00433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_93_1016 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08785_ rf_ram.memory\[141\]\[1\] _04186_ _04188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05997_ rf_ram.memory\[522\]\[1\] _01532_ _01521_ rf_ram.memory\[523\]\[1\] _01517_
+ rf_ram.memory\[521\]\[1\] _02192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XANTENNA__06382__A2 _01649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07736_ _02813_ _03496_ _03522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_0_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_49_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_49_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08659__A1 _04094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06119__C1 _01519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07667_ rf_ram.memory\[403\]\[0\] _03478_ _03479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06134__A2 _01785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09406_ net226 _03991_ _04576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06618_ rf_ram.memory\[236\]\[1\] _02789_ _02791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_94_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09459__I0 net79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07598_ net239 _03390_ _03436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_36_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10218__A1 _05081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06549_ _02732_ _02734_ _02735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XTAP_TAPCELL_ROW_62_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09084__A1 _04364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09337_ _04466_ _04536_ _04538_ _00992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_180_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_164_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09268_ _01418_ _01464_ _01366_ _04493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_63_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08219_ rf_ram.memory\[534\]\[1\] _03821_ _03824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_106_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09199_ _02805_ _04418_ _04445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_160_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11230_ _00966_ clknet_leaf_238_clk cpu.genblk3.csr.mstatus_mie vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_31_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09631__I0 cpu.decode.opcode\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07398__A1 _03289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11161_ _00897_ clknet_leaf_67_clk rf_ram.memory\[100\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_output74_I net74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05528__I _01643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10112_ _05014_ _05034_ _05035_ _01271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_8_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11092_ _00829_ clknet_leaf_98_clk rf_ram.memory\[419\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_41_1173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05972__B _01563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10043_ _02812_ _03158_ _04993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_141_3006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_141_3017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07570__A1 _03393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06373__A2 _01641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09311__A2 net62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10945_ _00683_ clknet_leaf_108_clk rf_ram.memory\[379\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_82_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06125__A2 _01770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07322__A1 _03260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_1172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07873__A2 _02954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10876_ _00620_ clknet_leaf_283_clk rf_ram.memory\[244\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_156_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10209__A1 net245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_156_3293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07625__A2 _03452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08822__A1 _04202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_117_2565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_117_2576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_4 _01804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11428_ _01160_ clknet_leaf_212_clk rf_ram.memory\[249\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_134_2890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07389__A1 _03292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11359_ _01091_ clknet_leaf_22_clk rf_ram.memory\[72\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_158_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08050__A2 _03693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05438__I _01633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05939__A2 _01605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05920_ _01909_ _02114_ _02115_ _02116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__05882__B _01551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08889__A1 _04234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06349__C1 _01725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05851_ rf_ram.memory\[238\]\[0\] _01501_ _02047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_83_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07561__A1 _02935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06364__A2 _01523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08570_ _04023_ _04051_ _04052_ _00711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_89_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05782_ _01493_ _01978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_07521_ rf_ram.memory\[322\]\[1\] _03386_ _03388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_76_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06116__A2 _01652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07452_ rf_ram.memory\[368\]\[1\] _03343_ _03345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_176_3658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_176_3669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06403_ rf_ram.memory\[84\]\[1\] _01509_ _01656_ rf_ram.memory\[85\]\[1\] _01763_
+ rf_ram.memory\[87\]\[1\] _02598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_135_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07383_ rf_ram.memory\[266\]\[1\] _03300_ _03302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09066__A1 rf_ram.memory\[0\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09122_ _02742_ _04396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_06334_ rf_ram.memory\[218\]\[1\] _01940_ _02019_ rf_ram.memory\[219\]\[1\] _02528_
+ _02529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__07616__A2 _03446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_40_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_40_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_161_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09053_ rf_ram.memory\[102\]\[1\] _04352_ _04354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06265_ net252 _02432_ _02459_ _02460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_26_981 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08004_ _02747_ _03689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_128_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05216_ _01413_ _01415_ _01416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_124_1005 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06196_ _02379_ _02383_ _02387_ _02390_ _02391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_clkbuf_5_16__f_clk_I clknet_3_4_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_1102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xmax_cap240 _02888_ net240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_102_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xmax_cap251 net252 net251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_05147_ _01349_ _01350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_111_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05348__I _01543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09955_ rf_ram.memory\[336\]\[0\] _04938_ _04939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_5_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08906_ _04237_ _04260_ _04262_ _00837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09886_ _03892_ _02822_ _04896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08837_ _04202_ _04219_ _04220_ _00810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_99_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_170_1003 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08768_ rf_ram.memory\[144\]\[0\] _04177_ _04178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_169_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07719_ _03491_ _03509_ _03511_ _00401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_71_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_1167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07304__A1 _03225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08699_ _02828_ _02921_ _04134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_135_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10730_ _00474_ clknet_leaf_77_clk rf_ram.memory\[443\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_32_1128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_1188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_24_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09057__A1 _04331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10661_ _00405_ clknet_leaf_129_clk rf_ram.memory\[37\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_119_950 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06128__B _01693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08804__A1 rf_ram.memory\[13\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10592_ _00336_ clknet_leaf_204_clk rf_ram.memory\[35\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_152_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_1251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05618__A1 _01600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06291__A1 _01909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_160_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_79_1870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_142_1127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11213_ _00949_ clknet_leaf_65_clk rf_ram.memory\[70\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_142_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06043__A1 _01603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_112_2473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_75_1789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_112_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11144_ _00880_ clknet_leaf_71_clk rf_ram.memory\[108\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09780__A2 _04067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput74 net74 o_dbus_adr[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput85 net85 o_dbus_adr[28] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__07791__A1 _03554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput96 net96 o_dbus_adr[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_11075_ _00812_ clknet_leaf_25_clk rf_ram.memory\[134\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_76_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10026_ _04396_ _04982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__07543__A1 _03389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06346__A2 _01808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_188_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_76_1066 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_99_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_1099 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_158_3322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_158_3333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10928_ _00672_ clknet_leaf_7_clk rf_ram.memory\[175\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_86_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_129_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_119_2605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_183_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10859_ _00603_ clknet_leaf_314_clk rf_ram.memory\[527\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_119_2616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06038__B _01351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_171_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_136_2930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_171_3566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_171_3577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_147_1027 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_41_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05877__B _02072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_1173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_14_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06050_ rf_ram.memory\[362\]\[1\] _01606_ _01608_ rf_ram.memory\[363\]\[1\] _02244_
+ _02245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_48_1168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_132_2849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06552__I _02737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_1059 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_160_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_22_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07782__A1 _03524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06585__A2 _02766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06952_ rf_ram.memory\[231\]\[0\] _03029_ _03030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09740_ _04804_ net16 _04805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__08479__I _03967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
.ends

