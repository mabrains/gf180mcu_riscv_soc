magic
tech gf180mcuD
magscale 1 5
timestamp 1700747289
<< obsm1 >>
rect 672 1415 11392 8262
<< metal2 >>
rect 784 9600 840 10000
rect 2240 9600 2296 10000
rect 3696 9600 3752 10000
rect 5152 9600 5208 10000
rect 6608 9600 6664 10000
rect 8064 9600 8120 10000
rect 9520 9600 9576 10000
rect 10976 9600 11032 10000
rect 1568 0 1624 400
rect 1792 0 1848 400
rect 2016 0 2072 400
rect 2240 0 2296 400
rect 2464 0 2520 400
rect 2688 0 2744 400
rect 2912 0 2968 400
rect 3136 0 3192 400
rect 3360 0 3416 400
rect 3584 0 3640 400
rect 3808 0 3864 400
rect 4032 0 4088 400
rect 4256 0 4312 400
rect 4480 0 4536 400
rect 4704 0 4760 400
rect 4928 0 4984 400
rect 5152 0 5208 400
rect 5376 0 5432 400
rect 5600 0 5656 400
rect 5824 0 5880 400
rect 6048 0 6104 400
rect 6272 0 6328 400
rect 6496 0 6552 400
rect 6720 0 6776 400
rect 6944 0 7000 400
rect 7168 0 7224 400
rect 7392 0 7448 400
rect 7616 0 7672 400
rect 7840 0 7896 400
rect 8064 0 8120 400
rect 8288 0 8344 400
rect 8512 0 8568 400
rect 8736 0 8792 400
rect 8960 0 9016 400
rect 9184 0 9240 400
rect 9408 0 9464 400
rect 9632 0 9688 400
rect 9856 0 9912 400
rect 10080 0 10136 400
rect 10304 0 10360 400
<< obsm2 >>
rect 742 9570 754 9600
rect 870 9570 2210 9600
rect 2326 9570 3666 9600
rect 3782 9570 5122 9600
rect 5238 9570 6578 9600
rect 6694 9570 8034 9600
rect 8150 9570 9490 9600
rect 9606 9570 10946 9600
rect 11062 9570 11378 9600
rect 742 430 11378 9570
rect 742 400 1538 430
rect 1654 400 1762 430
rect 1878 400 1986 430
rect 2102 400 2210 430
rect 2326 400 2434 430
rect 2550 400 2658 430
rect 2774 400 2882 430
rect 2998 400 3106 430
rect 3222 400 3330 430
rect 3446 400 3554 430
rect 3670 400 3778 430
rect 3894 400 4002 430
rect 4118 400 4226 430
rect 4342 400 4450 430
rect 4566 400 4674 430
rect 4790 400 4898 430
rect 5014 400 5122 430
rect 5238 400 5346 430
rect 5462 400 5570 430
rect 5686 400 5794 430
rect 5910 400 6018 430
rect 6134 400 6242 430
rect 6358 400 6466 430
rect 6582 400 6690 430
rect 6806 400 6914 430
rect 7030 400 7138 430
rect 7254 400 7362 430
rect 7478 400 7586 430
rect 7702 400 7810 430
rect 7926 400 8034 430
rect 8150 400 8258 430
rect 8374 400 8482 430
rect 8598 400 8706 430
rect 8822 400 8930 430
rect 9046 400 9154 430
rect 9270 400 9378 430
rect 9494 400 9602 430
rect 9718 400 9826 430
rect 9942 400 10050 430
rect 10166 400 10274 430
rect 10390 400 11378 430
<< metal3 >>
rect 0 8624 400 8680
rect 11600 8624 12000 8680
rect 0 8400 400 8456
rect 0 8176 400 8232
rect 0 7952 400 8008
rect 0 7728 400 7784
rect 0 7504 400 7560
rect 0 7280 400 7336
rect 0 7056 400 7112
rect 0 6832 400 6888
rect 0 6608 400 6664
rect 0 6384 400 6440
rect 0 6160 400 6216
rect 11600 6160 12000 6216
rect 0 5936 400 5992
rect 0 5712 400 5768
rect 0 5488 400 5544
rect 0 5264 400 5320
rect 0 5040 400 5096
rect 0 4816 400 4872
rect 0 4592 400 4648
rect 0 4368 400 4424
rect 0 4144 400 4200
rect 0 3920 400 3976
rect 0 3696 400 3752
rect 11600 3696 12000 3752
rect 0 3472 400 3528
rect 0 3248 400 3304
rect 0 3024 400 3080
rect 0 2800 400 2856
rect 0 2576 400 2632
rect 0 2352 400 2408
rect 0 2128 400 2184
rect 0 1904 400 1960
rect 0 1680 400 1736
rect 0 1456 400 1512
rect 0 1232 400 1288
rect 11600 1232 12000 1288
<< obsm3 >>
rect 430 8594 11570 8666
rect 400 8486 11600 8594
rect 430 8370 11600 8486
rect 400 8262 11600 8370
rect 430 8146 11600 8262
rect 400 8038 11600 8146
rect 430 7922 11600 8038
rect 400 7814 11600 7922
rect 430 7698 11600 7814
rect 400 7590 11600 7698
rect 430 7474 11600 7590
rect 400 7366 11600 7474
rect 430 7250 11600 7366
rect 400 7142 11600 7250
rect 430 7026 11600 7142
rect 400 6918 11600 7026
rect 430 6802 11600 6918
rect 400 6694 11600 6802
rect 430 6578 11600 6694
rect 400 6470 11600 6578
rect 430 6354 11600 6470
rect 400 6246 11600 6354
rect 430 6130 11570 6246
rect 400 6022 11600 6130
rect 430 5906 11600 6022
rect 400 5798 11600 5906
rect 430 5682 11600 5798
rect 400 5574 11600 5682
rect 430 5458 11600 5574
rect 400 5350 11600 5458
rect 430 5234 11600 5350
rect 400 5126 11600 5234
rect 430 5010 11600 5126
rect 400 4902 11600 5010
rect 430 4786 11600 4902
rect 400 4678 11600 4786
rect 430 4562 11600 4678
rect 400 4454 11600 4562
rect 430 4338 11600 4454
rect 400 4230 11600 4338
rect 430 4114 11600 4230
rect 400 4006 11600 4114
rect 430 3890 11600 4006
rect 400 3782 11600 3890
rect 430 3666 11570 3782
rect 400 3558 11600 3666
rect 430 3442 11600 3558
rect 400 3334 11600 3442
rect 430 3218 11600 3334
rect 400 3110 11600 3218
rect 430 2994 11600 3110
rect 400 2886 11600 2994
rect 430 2770 11600 2886
rect 400 2662 11600 2770
rect 430 2546 11600 2662
rect 400 2438 11600 2546
rect 430 2322 11600 2438
rect 400 2214 11600 2322
rect 430 2098 11600 2214
rect 400 1990 11600 2098
rect 430 1874 11600 1990
rect 400 1766 11600 1874
rect 430 1650 11600 1766
rect 400 1542 11600 1650
rect 430 1426 11600 1542
rect 400 1318 11600 1426
rect 430 1246 11570 1318
<< metal4 >>
rect 1922 1538 2082 8262
rect 3252 1538 3412 8262
rect 4582 1538 4742 8262
rect 5912 1538 6072 8262
rect 7242 1538 7402 8262
rect 8572 1538 8732 8262
rect 9902 1538 10062 8262
rect 11232 1538 11392 8262
<< obsm4 >>
rect 910 1633 1892 6039
rect 2112 1633 3222 6039
rect 3442 1633 4552 6039
rect 4772 1633 5882 6039
rect 6102 1633 7212 6039
rect 7432 1633 8542 6039
rect 8762 1633 9842 6039
<< labels >>
rlabel metal3 s 11600 1232 12000 1288 6 buttons[0]
port 1 nsew signal input
rlabel metal3 s 11600 6160 12000 6216 6 buttons[1]
port 2 nsew signal input
rlabel metal3 s 11600 8624 12000 8680 6 buttons_enb[0]
port 3 nsew signal output
rlabel metal3 s 11600 3696 12000 3752 6 buttons_enb[1]
port 4 nsew signal output
rlabel metal2 s 9856 0 9912 400 6 clk
port 5 nsew signal input
rlabel metal2 s 10080 0 10136 400 6 clk2
port 6 nsew signal input
rlabel metal2 s 2240 0 2296 400 6 i_wb_addr[0]
port 7 nsew signal input
rlabel metal2 s 4928 0 4984 400 6 i_wb_addr[10]
port 8 nsew signal input
rlabel metal2 s 5152 0 5208 400 6 i_wb_addr[11]
port 9 nsew signal input
rlabel metal2 s 5376 0 5432 400 6 i_wb_addr[12]
port 10 nsew signal input
rlabel metal2 s 5600 0 5656 400 6 i_wb_addr[13]
port 11 nsew signal input
rlabel metal2 s 5824 0 5880 400 6 i_wb_addr[14]
port 12 nsew signal input
rlabel metal2 s 6048 0 6104 400 6 i_wb_addr[15]
port 13 nsew signal input
rlabel metal2 s 6272 0 6328 400 6 i_wb_addr[16]
port 14 nsew signal input
rlabel metal2 s 6496 0 6552 400 6 i_wb_addr[17]
port 15 nsew signal input
rlabel metal2 s 6720 0 6776 400 6 i_wb_addr[18]
port 16 nsew signal input
rlabel metal2 s 6944 0 7000 400 6 i_wb_addr[19]
port 17 nsew signal input
rlabel metal2 s 2688 0 2744 400 6 i_wb_addr[1]
port 18 nsew signal input
rlabel metal2 s 7168 0 7224 400 6 i_wb_addr[20]
port 19 nsew signal input
rlabel metal2 s 7392 0 7448 400 6 i_wb_addr[21]
port 20 nsew signal input
rlabel metal2 s 7616 0 7672 400 6 i_wb_addr[22]
port 21 nsew signal input
rlabel metal2 s 7840 0 7896 400 6 i_wb_addr[23]
port 22 nsew signal input
rlabel metal2 s 8064 0 8120 400 6 i_wb_addr[24]
port 23 nsew signal input
rlabel metal2 s 8288 0 8344 400 6 i_wb_addr[25]
port 24 nsew signal input
rlabel metal2 s 8512 0 8568 400 6 i_wb_addr[26]
port 25 nsew signal input
rlabel metal2 s 8736 0 8792 400 6 i_wb_addr[27]
port 26 nsew signal input
rlabel metal2 s 8960 0 9016 400 6 i_wb_addr[28]
port 27 nsew signal input
rlabel metal2 s 9184 0 9240 400 6 i_wb_addr[29]
port 28 nsew signal input
rlabel metal2 s 3136 0 3192 400 6 i_wb_addr[2]
port 29 nsew signal input
rlabel metal2 s 9408 0 9464 400 6 i_wb_addr[30]
port 30 nsew signal input
rlabel metal2 s 9632 0 9688 400 6 i_wb_addr[31]
port 31 nsew signal input
rlabel metal2 s 3360 0 3416 400 6 i_wb_addr[3]
port 32 nsew signal input
rlabel metal2 s 3584 0 3640 400 6 i_wb_addr[4]
port 33 nsew signal input
rlabel metal2 s 3808 0 3864 400 6 i_wb_addr[5]
port 34 nsew signal input
rlabel metal2 s 4032 0 4088 400 6 i_wb_addr[6]
port 35 nsew signal input
rlabel metal2 s 4256 0 4312 400 6 i_wb_addr[7]
port 36 nsew signal input
rlabel metal2 s 4480 0 4536 400 6 i_wb_addr[8]
port 37 nsew signal input
rlabel metal2 s 4704 0 4760 400 6 i_wb_addr[9]
port 38 nsew signal input
rlabel metal2 s 1568 0 1624 400 6 i_wb_cyc
port 39 nsew signal input
rlabel metal2 s 2464 0 2520 400 6 i_wb_data[0]
port 40 nsew signal input
rlabel metal2 s 2912 0 2968 400 6 i_wb_data[1]
port 41 nsew signal input
rlabel metal2 s 1792 0 1848 400 6 i_wb_stb
port 42 nsew signal input
rlabel metal2 s 2016 0 2072 400 6 i_wb_we
port 43 nsew signal input
rlabel metal2 s 6608 9600 6664 10000 6 led_enb[0]
port 44 nsew signal output
rlabel metal2 s 9520 9600 9576 10000 6 led_enb[1]
port 45 nsew signal output
rlabel metal2 s 8064 9600 8120 10000 6 leds[0]
port 46 nsew signal output
rlabel metal2 s 10976 9600 11032 10000 6 leds[1]
port 47 nsew signal output
rlabel metal3 s 0 1232 400 1288 6 o_wb_ack
port 48 nsew signal output
rlabel metal3 s 0 1680 400 1736 6 o_wb_data[0]
port 49 nsew signal output
rlabel metal3 s 0 3920 400 3976 6 o_wb_data[10]
port 50 nsew signal output
rlabel metal3 s 0 4144 400 4200 6 o_wb_data[11]
port 51 nsew signal output
rlabel metal3 s 0 4368 400 4424 6 o_wb_data[12]
port 52 nsew signal output
rlabel metal3 s 0 4592 400 4648 6 o_wb_data[13]
port 53 nsew signal output
rlabel metal3 s 0 4816 400 4872 6 o_wb_data[14]
port 54 nsew signal output
rlabel metal3 s 0 5040 400 5096 6 o_wb_data[15]
port 55 nsew signal output
rlabel metal3 s 0 5264 400 5320 6 o_wb_data[16]
port 56 nsew signal output
rlabel metal3 s 0 5488 400 5544 6 o_wb_data[17]
port 57 nsew signal output
rlabel metal3 s 0 5712 400 5768 6 o_wb_data[18]
port 58 nsew signal output
rlabel metal3 s 0 5936 400 5992 6 o_wb_data[19]
port 59 nsew signal output
rlabel metal3 s 0 1904 400 1960 6 o_wb_data[1]
port 60 nsew signal output
rlabel metal3 s 0 6160 400 6216 6 o_wb_data[20]
port 61 nsew signal output
rlabel metal3 s 0 6384 400 6440 6 o_wb_data[21]
port 62 nsew signal output
rlabel metal3 s 0 6608 400 6664 6 o_wb_data[22]
port 63 nsew signal output
rlabel metal3 s 0 6832 400 6888 6 o_wb_data[23]
port 64 nsew signal output
rlabel metal3 s 0 7056 400 7112 6 o_wb_data[24]
port 65 nsew signal output
rlabel metal3 s 0 7280 400 7336 6 o_wb_data[25]
port 66 nsew signal output
rlabel metal3 s 0 7504 400 7560 6 o_wb_data[26]
port 67 nsew signal output
rlabel metal3 s 0 7728 400 7784 6 o_wb_data[27]
port 68 nsew signal output
rlabel metal3 s 0 7952 400 8008 6 o_wb_data[28]
port 69 nsew signal output
rlabel metal3 s 0 8176 400 8232 6 o_wb_data[29]
port 70 nsew signal output
rlabel metal3 s 0 2128 400 2184 6 o_wb_data[2]
port 71 nsew signal output
rlabel metal3 s 0 8400 400 8456 6 o_wb_data[30]
port 72 nsew signal output
rlabel metal3 s 0 8624 400 8680 6 o_wb_data[31]
port 73 nsew signal output
rlabel metal3 s 0 2352 400 2408 6 o_wb_data[3]
port 74 nsew signal output
rlabel metal3 s 0 2576 400 2632 6 o_wb_data[4]
port 75 nsew signal output
rlabel metal3 s 0 2800 400 2856 6 o_wb_data[5]
port 76 nsew signal output
rlabel metal3 s 0 3024 400 3080 6 o_wb_data[6]
port 77 nsew signal output
rlabel metal3 s 0 3248 400 3304 6 o_wb_data[7]
port 78 nsew signal output
rlabel metal3 s 0 3472 400 3528 6 o_wb_data[8]
port 79 nsew signal output
rlabel metal3 s 0 3696 400 3752 6 o_wb_data[9]
port 80 nsew signal output
rlabel metal3 s 0 1456 400 1512 6 o_wb_stall
port 81 nsew signal output
rlabel metal2 s 10304 0 10360 400 6 reset
port 82 nsew signal input
rlabel metal4 s 1922 1538 2082 8262 6 vdd
port 83 nsew power bidirectional
rlabel metal4 s 4582 1538 4742 8262 6 vdd
port 83 nsew power bidirectional
rlabel metal4 s 7242 1538 7402 8262 6 vdd
port 83 nsew power bidirectional
rlabel metal4 s 9902 1538 10062 8262 6 vdd
port 83 nsew power bidirectional
rlabel metal4 s 3252 1538 3412 8262 6 vss
port 84 nsew ground bidirectional
rlabel metal4 s 5912 1538 6072 8262 6 vss
port 84 nsew ground bidirectional
rlabel metal4 s 8572 1538 8732 8262 6 vss
port 84 nsew ground bidirectional
rlabel metal4 s 11232 1538 11392 8262 6 vss
port 84 nsew ground bidirectional
rlabel metal2 s 2240 9600 2296 10000 6 xtal_clk[0]
port 85 nsew signal output
rlabel metal2 s 5152 9600 5208 10000 6 xtal_clk[1]
port 86 nsew signal output
rlabel metal2 s 784 9600 840 10000 6 xtal_clk_enb[0]
port 87 nsew signal output
rlabel metal2 s 3696 9600 3752 10000 6 xtal_clk_enb[1]
port 88 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 12000 10000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 420812
string GDS_FILE /home/farag/carvel_riscv_soc/gf180mcu_riscv_soc/openlane/wb_buttons_leds/runs/23_11_23_15_45/results/signoff/wb_buttons_leds.magic.gds
string GDS_START 138408
<< end >>

