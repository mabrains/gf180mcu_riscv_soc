magic
tech gf180mcuD
magscale 1 10
timestamp 1700928318
<< metal1 >>
rect 37202 46510 37214 46562
rect 37266 46559 37278 46562
rect 37874 46559 37886 46562
rect 37266 46513 37886 46559
rect 37266 46510 37278 46513
rect 37874 46510 37886 46513
rect 37938 46510 37950 46562
rect 1344 46282 38640 46316
rect 1344 46230 4024 46282
rect 4076 46230 4148 46282
rect 4200 46230 4272 46282
rect 4324 46230 4396 46282
rect 4448 46230 4520 46282
rect 4572 46230 4644 46282
rect 4696 46230 4768 46282
rect 4820 46230 4892 46282
rect 4944 46230 5016 46282
rect 5068 46230 5140 46282
rect 5192 46230 24024 46282
rect 24076 46230 24148 46282
rect 24200 46230 24272 46282
rect 24324 46230 24396 46282
rect 24448 46230 24520 46282
rect 24572 46230 24644 46282
rect 24696 46230 24768 46282
rect 24820 46230 24892 46282
rect 24944 46230 25016 46282
rect 25068 46230 25140 46282
rect 25192 46230 38640 46282
rect 1344 46196 38640 46230
rect 2706 45950 2718 46002
rect 2770 45950 2782 46002
rect 13570 45950 13582 46002
rect 13634 45950 13646 46002
rect 28802 45950 28814 46002
rect 28866 45950 28878 46002
rect 37874 45950 37886 46002
rect 37938 45950 37950 46002
rect 14814 45890 14866 45902
rect 3490 45838 3502 45890
rect 3554 45838 3566 45890
rect 14130 45838 14142 45890
rect 14194 45838 14206 45890
rect 14814 45826 14866 45838
rect 2046 45778 2098 45790
rect 2046 45714 2098 45726
rect 7870 45778 7922 45790
rect 7870 45714 7922 45726
rect 17726 45778 17778 45790
rect 17726 45714 17778 45726
rect 22654 45778 22706 45790
rect 22654 45714 22706 45726
rect 32510 45778 32562 45790
rect 32510 45714 32562 45726
rect 27918 45666 27970 45678
rect 27918 45602 27970 45614
rect 28366 45666 28418 45678
rect 28366 45602 28418 45614
rect 37214 45666 37266 45678
rect 37214 45602 37266 45614
rect 37438 45666 37490 45678
rect 37438 45602 37490 45614
rect 1344 45498 38640 45532
rect 1344 45446 14024 45498
rect 14076 45446 14148 45498
rect 14200 45446 14272 45498
rect 14324 45446 14396 45498
rect 14448 45446 14520 45498
rect 14572 45446 14644 45498
rect 14696 45446 14768 45498
rect 14820 45446 14892 45498
rect 14944 45446 15016 45498
rect 15068 45446 15140 45498
rect 15192 45446 34024 45498
rect 34076 45446 34148 45498
rect 34200 45446 34272 45498
rect 34324 45446 34396 45498
rect 34448 45446 34520 45498
rect 34572 45446 34644 45498
rect 34696 45446 34768 45498
rect 34820 45446 34892 45498
rect 34944 45446 35016 45498
rect 35068 45446 35140 45498
rect 35192 45446 38640 45498
rect 1344 45412 38640 45446
rect 2158 45330 2210 45342
rect 2158 45266 2210 45278
rect 1710 45218 1762 45230
rect 1710 45154 1762 45166
rect 2718 44994 2770 45006
rect 2718 44930 2770 44942
rect 1344 44714 38640 44748
rect 1344 44662 4024 44714
rect 4076 44662 4148 44714
rect 4200 44662 4272 44714
rect 4324 44662 4396 44714
rect 4448 44662 4520 44714
rect 4572 44662 4644 44714
rect 4696 44662 4768 44714
rect 4820 44662 4892 44714
rect 4944 44662 5016 44714
rect 5068 44662 5140 44714
rect 5192 44662 24024 44714
rect 24076 44662 24148 44714
rect 24200 44662 24272 44714
rect 24324 44662 24396 44714
rect 24448 44662 24520 44714
rect 24572 44662 24644 44714
rect 24696 44662 24768 44714
rect 24820 44662 24892 44714
rect 24944 44662 25016 44714
rect 25068 44662 25140 44714
rect 25192 44662 38640 44714
rect 1344 44628 38640 44662
rect 1344 43930 38640 43964
rect 1344 43878 14024 43930
rect 14076 43878 14148 43930
rect 14200 43878 14272 43930
rect 14324 43878 14396 43930
rect 14448 43878 14520 43930
rect 14572 43878 14644 43930
rect 14696 43878 14768 43930
rect 14820 43878 14892 43930
rect 14944 43878 15016 43930
rect 15068 43878 15140 43930
rect 15192 43878 34024 43930
rect 34076 43878 34148 43930
rect 34200 43878 34272 43930
rect 34324 43878 34396 43930
rect 34448 43878 34520 43930
rect 34572 43878 34644 43930
rect 34696 43878 34768 43930
rect 34820 43878 34892 43930
rect 34944 43878 35016 43930
rect 35068 43878 35140 43930
rect 35192 43878 38640 43930
rect 1344 43844 38640 43878
rect 1710 43650 1762 43662
rect 1710 43586 1762 43598
rect 38222 43314 38274 43326
rect 38222 43250 38274 43262
rect 1344 43146 38640 43180
rect 1344 43094 4024 43146
rect 4076 43094 4148 43146
rect 4200 43094 4272 43146
rect 4324 43094 4396 43146
rect 4448 43094 4520 43146
rect 4572 43094 4644 43146
rect 4696 43094 4768 43146
rect 4820 43094 4892 43146
rect 4944 43094 5016 43146
rect 5068 43094 5140 43146
rect 5192 43094 24024 43146
rect 24076 43094 24148 43146
rect 24200 43094 24272 43146
rect 24324 43094 24396 43146
rect 24448 43094 24520 43146
rect 24572 43094 24644 43146
rect 24696 43094 24768 43146
rect 24820 43094 24892 43146
rect 24944 43094 25016 43146
rect 25068 43094 25140 43146
rect 25192 43094 38640 43146
rect 1344 43060 38640 43094
rect 1344 42362 38640 42396
rect 1344 42310 14024 42362
rect 14076 42310 14148 42362
rect 14200 42310 14272 42362
rect 14324 42310 14396 42362
rect 14448 42310 14520 42362
rect 14572 42310 14644 42362
rect 14696 42310 14768 42362
rect 14820 42310 14892 42362
rect 14944 42310 15016 42362
rect 15068 42310 15140 42362
rect 15192 42310 34024 42362
rect 34076 42310 34148 42362
rect 34200 42310 34272 42362
rect 34324 42310 34396 42362
rect 34448 42310 34520 42362
rect 34572 42310 34644 42362
rect 34696 42310 34768 42362
rect 34820 42310 34892 42362
rect 34944 42310 35016 42362
rect 35068 42310 35140 42362
rect 35192 42310 38640 42362
rect 1344 42276 38640 42310
rect 1710 42082 1762 42094
rect 1710 42018 1762 42030
rect 1344 41578 38640 41612
rect 1344 41526 4024 41578
rect 4076 41526 4148 41578
rect 4200 41526 4272 41578
rect 4324 41526 4396 41578
rect 4448 41526 4520 41578
rect 4572 41526 4644 41578
rect 4696 41526 4768 41578
rect 4820 41526 4892 41578
rect 4944 41526 5016 41578
rect 5068 41526 5140 41578
rect 5192 41526 24024 41578
rect 24076 41526 24148 41578
rect 24200 41526 24272 41578
rect 24324 41526 24396 41578
rect 24448 41526 24520 41578
rect 24572 41526 24644 41578
rect 24696 41526 24768 41578
rect 24820 41526 24892 41578
rect 24944 41526 25016 41578
rect 25068 41526 25140 41578
rect 25192 41526 38640 41578
rect 1344 41492 38640 41526
rect 1710 40962 1762 40974
rect 1710 40898 1762 40910
rect 1344 40794 38640 40828
rect 1344 40742 14024 40794
rect 14076 40742 14148 40794
rect 14200 40742 14272 40794
rect 14324 40742 14396 40794
rect 14448 40742 14520 40794
rect 14572 40742 14644 40794
rect 14696 40742 14768 40794
rect 14820 40742 14892 40794
rect 14944 40742 15016 40794
rect 15068 40742 15140 40794
rect 15192 40742 34024 40794
rect 34076 40742 34148 40794
rect 34200 40742 34272 40794
rect 34324 40742 34396 40794
rect 34448 40742 34520 40794
rect 34572 40742 34644 40794
rect 34696 40742 34768 40794
rect 34820 40742 34892 40794
rect 34944 40742 35016 40794
rect 35068 40742 35140 40794
rect 35192 40742 38640 40794
rect 1344 40708 38640 40742
rect 1344 40010 38640 40044
rect 1344 39958 4024 40010
rect 4076 39958 4148 40010
rect 4200 39958 4272 40010
rect 4324 39958 4396 40010
rect 4448 39958 4520 40010
rect 4572 39958 4644 40010
rect 4696 39958 4768 40010
rect 4820 39958 4892 40010
rect 4944 39958 5016 40010
rect 5068 39958 5140 40010
rect 5192 39958 24024 40010
rect 24076 39958 24148 40010
rect 24200 39958 24272 40010
rect 24324 39958 24396 40010
rect 24448 39958 24520 40010
rect 24572 39958 24644 40010
rect 24696 39958 24768 40010
rect 24820 39958 24892 40010
rect 24944 39958 25016 40010
rect 25068 39958 25140 40010
rect 25192 39958 38640 40010
rect 1344 39924 38640 39958
rect 1710 39394 1762 39406
rect 1710 39330 1762 39342
rect 1344 39226 38640 39260
rect 1344 39174 14024 39226
rect 14076 39174 14148 39226
rect 14200 39174 14272 39226
rect 14324 39174 14396 39226
rect 14448 39174 14520 39226
rect 14572 39174 14644 39226
rect 14696 39174 14768 39226
rect 14820 39174 14892 39226
rect 14944 39174 15016 39226
rect 15068 39174 15140 39226
rect 15192 39174 34024 39226
rect 34076 39174 34148 39226
rect 34200 39174 34272 39226
rect 34324 39174 34396 39226
rect 34448 39174 34520 39226
rect 34572 39174 34644 39226
rect 34696 39174 34768 39226
rect 34820 39174 34892 39226
rect 34944 39174 35016 39226
rect 35068 39174 35140 39226
rect 35192 39174 38640 39226
rect 1344 39140 38640 39174
rect 1344 38442 38640 38476
rect 1344 38390 4024 38442
rect 4076 38390 4148 38442
rect 4200 38390 4272 38442
rect 4324 38390 4396 38442
rect 4448 38390 4520 38442
rect 4572 38390 4644 38442
rect 4696 38390 4768 38442
rect 4820 38390 4892 38442
rect 4944 38390 5016 38442
rect 5068 38390 5140 38442
rect 5192 38390 24024 38442
rect 24076 38390 24148 38442
rect 24200 38390 24272 38442
rect 24324 38390 24396 38442
rect 24448 38390 24520 38442
rect 24572 38390 24644 38442
rect 24696 38390 24768 38442
rect 24820 38390 24892 38442
rect 24944 38390 25016 38442
rect 25068 38390 25140 38442
rect 25192 38390 38640 38442
rect 1344 38356 38640 38390
rect 1710 37826 1762 37838
rect 1710 37762 1762 37774
rect 1344 37658 38640 37692
rect 1344 37606 14024 37658
rect 14076 37606 14148 37658
rect 14200 37606 14272 37658
rect 14324 37606 14396 37658
rect 14448 37606 14520 37658
rect 14572 37606 14644 37658
rect 14696 37606 14768 37658
rect 14820 37606 14892 37658
rect 14944 37606 15016 37658
rect 15068 37606 15140 37658
rect 15192 37606 34024 37658
rect 34076 37606 34148 37658
rect 34200 37606 34272 37658
rect 34324 37606 34396 37658
rect 34448 37606 34520 37658
rect 34572 37606 34644 37658
rect 34696 37606 34768 37658
rect 34820 37606 34892 37658
rect 34944 37606 35016 37658
rect 35068 37606 35140 37658
rect 35192 37606 38640 37658
rect 1344 37572 38640 37606
rect 1344 36874 38640 36908
rect 1344 36822 4024 36874
rect 4076 36822 4148 36874
rect 4200 36822 4272 36874
rect 4324 36822 4396 36874
rect 4448 36822 4520 36874
rect 4572 36822 4644 36874
rect 4696 36822 4768 36874
rect 4820 36822 4892 36874
rect 4944 36822 5016 36874
rect 5068 36822 5140 36874
rect 5192 36822 24024 36874
rect 24076 36822 24148 36874
rect 24200 36822 24272 36874
rect 24324 36822 24396 36874
rect 24448 36822 24520 36874
rect 24572 36822 24644 36874
rect 24696 36822 24768 36874
rect 24820 36822 24892 36874
rect 24944 36822 25016 36874
rect 25068 36822 25140 36874
rect 25192 36822 38640 36874
rect 1344 36788 38640 36822
rect 1710 36370 1762 36382
rect 1710 36306 1762 36318
rect 1344 36090 38640 36124
rect 1344 36038 14024 36090
rect 14076 36038 14148 36090
rect 14200 36038 14272 36090
rect 14324 36038 14396 36090
rect 14448 36038 14520 36090
rect 14572 36038 14644 36090
rect 14696 36038 14768 36090
rect 14820 36038 14892 36090
rect 14944 36038 15016 36090
rect 15068 36038 15140 36090
rect 15192 36038 34024 36090
rect 34076 36038 34148 36090
rect 34200 36038 34272 36090
rect 34324 36038 34396 36090
rect 34448 36038 34520 36090
rect 34572 36038 34644 36090
rect 34696 36038 34768 36090
rect 34820 36038 34892 36090
rect 34944 36038 35016 36090
rect 35068 36038 35140 36090
rect 35192 36038 38640 36090
rect 1344 36004 38640 36038
rect 1710 35810 1762 35822
rect 1710 35746 1762 35758
rect 1344 35306 38640 35340
rect 1344 35254 4024 35306
rect 4076 35254 4148 35306
rect 4200 35254 4272 35306
rect 4324 35254 4396 35306
rect 4448 35254 4520 35306
rect 4572 35254 4644 35306
rect 4696 35254 4768 35306
rect 4820 35254 4892 35306
rect 4944 35254 5016 35306
rect 5068 35254 5140 35306
rect 5192 35254 24024 35306
rect 24076 35254 24148 35306
rect 24200 35254 24272 35306
rect 24324 35254 24396 35306
rect 24448 35254 24520 35306
rect 24572 35254 24644 35306
rect 24696 35254 24768 35306
rect 24820 35254 24892 35306
rect 24944 35254 25016 35306
rect 25068 35254 25140 35306
rect 25192 35254 38640 35306
rect 1344 35220 38640 35254
rect 1344 34522 38640 34556
rect 1344 34470 14024 34522
rect 14076 34470 14148 34522
rect 14200 34470 14272 34522
rect 14324 34470 14396 34522
rect 14448 34470 14520 34522
rect 14572 34470 14644 34522
rect 14696 34470 14768 34522
rect 14820 34470 14892 34522
rect 14944 34470 15016 34522
rect 15068 34470 15140 34522
rect 15192 34470 34024 34522
rect 34076 34470 34148 34522
rect 34200 34470 34272 34522
rect 34324 34470 34396 34522
rect 34448 34470 34520 34522
rect 34572 34470 34644 34522
rect 34696 34470 34768 34522
rect 34820 34470 34892 34522
rect 34944 34470 35016 34522
rect 35068 34470 35140 34522
rect 35192 34470 38640 34522
rect 1344 34436 38640 34470
rect 1710 34242 1762 34254
rect 1710 34178 1762 34190
rect 1344 33738 38640 33772
rect 1344 33686 4024 33738
rect 4076 33686 4148 33738
rect 4200 33686 4272 33738
rect 4324 33686 4396 33738
rect 4448 33686 4520 33738
rect 4572 33686 4644 33738
rect 4696 33686 4768 33738
rect 4820 33686 4892 33738
rect 4944 33686 5016 33738
rect 5068 33686 5140 33738
rect 5192 33686 24024 33738
rect 24076 33686 24148 33738
rect 24200 33686 24272 33738
rect 24324 33686 24396 33738
rect 24448 33686 24520 33738
rect 24572 33686 24644 33738
rect 24696 33686 24768 33738
rect 24820 33686 24892 33738
rect 24944 33686 25016 33738
rect 25068 33686 25140 33738
rect 25192 33686 38640 33738
rect 1344 33652 38640 33686
rect 1344 32954 38640 32988
rect 1344 32902 14024 32954
rect 14076 32902 14148 32954
rect 14200 32902 14272 32954
rect 14324 32902 14396 32954
rect 14448 32902 14520 32954
rect 14572 32902 14644 32954
rect 14696 32902 14768 32954
rect 14820 32902 14892 32954
rect 14944 32902 15016 32954
rect 15068 32902 15140 32954
rect 15192 32902 34024 32954
rect 34076 32902 34148 32954
rect 34200 32902 34272 32954
rect 34324 32902 34396 32954
rect 34448 32902 34520 32954
rect 34572 32902 34644 32954
rect 34696 32902 34768 32954
rect 34820 32902 34892 32954
rect 34944 32902 35016 32954
rect 35068 32902 35140 32954
rect 35192 32902 38640 32954
rect 1344 32868 38640 32902
rect 1710 32674 1762 32686
rect 1710 32610 1762 32622
rect 1344 32170 38640 32204
rect 1344 32118 4024 32170
rect 4076 32118 4148 32170
rect 4200 32118 4272 32170
rect 4324 32118 4396 32170
rect 4448 32118 4520 32170
rect 4572 32118 4644 32170
rect 4696 32118 4768 32170
rect 4820 32118 4892 32170
rect 4944 32118 5016 32170
rect 5068 32118 5140 32170
rect 5192 32118 24024 32170
rect 24076 32118 24148 32170
rect 24200 32118 24272 32170
rect 24324 32118 24396 32170
rect 24448 32118 24520 32170
rect 24572 32118 24644 32170
rect 24696 32118 24768 32170
rect 24820 32118 24892 32170
rect 24944 32118 25016 32170
rect 25068 32118 25140 32170
rect 25192 32118 38640 32170
rect 1344 32084 38640 32118
rect 1710 31554 1762 31566
rect 1710 31490 1762 31502
rect 37662 31554 37714 31566
rect 38222 31554 38274 31566
rect 37874 31502 37886 31554
rect 37938 31502 37950 31554
rect 37662 31490 37714 31502
rect 38222 31490 38274 31502
rect 1344 31386 38640 31420
rect 1344 31334 14024 31386
rect 14076 31334 14148 31386
rect 14200 31334 14272 31386
rect 14324 31334 14396 31386
rect 14448 31334 14520 31386
rect 14572 31334 14644 31386
rect 14696 31334 14768 31386
rect 14820 31334 14892 31386
rect 14944 31334 15016 31386
rect 15068 31334 15140 31386
rect 15192 31334 34024 31386
rect 34076 31334 34148 31386
rect 34200 31334 34272 31386
rect 34324 31334 34396 31386
rect 34448 31334 34520 31386
rect 34572 31334 34644 31386
rect 34696 31334 34768 31386
rect 34820 31334 34892 31386
rect 34944 31334 35016 31386
rect 35068 31334 35140 31386
rect 35192 31334 38640 31386
rect 1344 31300 38640 31334
rect 1344 30602 38640 30636
rect 1344 30550 4024 30602
rect 4076 30550 4148 30602
rect 4200 30550 4272 30602
rect 4324 30550 4396 30602
rect 4448 30550 4520 30602
rect 4572 30550 4644 30602
rect 4696 30550 4768 30602
rect 4820 30550 4892 30602
rect 4944 30550 5016 30602
rect 5068 30550 5140 30602
rect 5192 30550 24024 30602
rect 24076 30550 24148 30602
rect 24200 30550 24272 30602
rect 24324 30550 24396 30602
rect 24448 30550 24520 30602
rect 24572 30550 24644 30602
rect 24696 30550 24768 30602
rect 24820 30550 24892 30602
rect 24944 30550 25016 30602
rect 25068 30550 25140 30602
rect 25192 30550 38640 30602
rect 1344 30516 38640 30550
rect 1710 29986 1762 29998
rect 1710 29922 1762 29934
rect 1344 29818 38640 29852
rect 1344 29766 14024 29818
rect 14076 29766 14148 29818
rect 14200 29766 14272 29818
rect 14324 29766 14396 29818
rect 14448 29766 14520 29818
rect 14572 29766 14644 29818
rect 14696 29766 14768 29818
rect 14820 29766 14892 29818
rect 14944 29766 15016 29818
rect 15068 29766 15140 29818
rect 15192 29766 34024 29818
rect 34076 29766 34148 29818
rect 34200 29766 34272 29818
rect 34324 29766 34396 29818
rect 34448 29766 34520 29818
rect 34572 29766 34644 29818
rect 34696 29766 34768 29818
rect 34820 29766 34892 29818
rect 34944 29766 35016 29818
rect 35068 29766 35140 29818
rect 35192 29766 38640 29818
rect 1344 29732 38640 29766
rect 1344 29034 38640 29068
rect 1344 28982 4024 29034
rect 4076 28982 4148 29034
rect 4200 28982 4272 29034
rect 4324 28982 4396 29034
rect 4448 28982 4520 29034
rect 4572 28982 4644 29034
rect 4696 28982 4768 29034
rect 4820 28982 4892 29034
rect 4944 28982 5016 29034
rect 5068 28982 5140 29034
rect 5192 28982 24024 29034
rect 24076 28982 24148 29034
rect 24200 28982 24272 29034
rect 24324 28982 24396 29034
rect 24448 28982 24520 29034
rect 24572 28982 24644 29034
rect 24696 28982 24768 29034
rect 24820 28982 24892 29034
rect 24944 28982 25016 29034
rect 25068 28982 25140 29034
rect 25192 28982 38640 29034
rect 1344 28948 38640 28982
rect 1710 28418 1762 28430
rect 1710 28354 1762 28366
rect 1344 28250 38640 28284
rect 1344 28198 14024 28250
rect 14076 28198 14148 28250
rect 14200 28198 14272 28250
rect 14324 28198 14396 28250
rect 14448 28198 14520 28250
rect 14572 28198 14644 28250
rect 14696 28198 14768 28250
rect 14820 28198 14892 28250
rect 14944 28198 15016 28250
rect 15068 28198 15140 28250
rect 15192 28198 34024 28250
rect 34076 28198 34148 28250
rect 34200 28198 34272 28250
rect 34324 28198 34396 28250
rect 34448 28198 34520 28250
rect 34572 28198 34644 28250
rect 34696 28198 34768 28250
rect 34820 28198 34892 28250
rect 34944 28198 35016 28250
rect 35068 28198 35140 28250
rect 35192 28198 38640 28250
rect 1344 28164 38640 28198
rect 1344 27466 38640 27500
rect 1344 27414 4024 27466
rect 4076 27414 4148 27466
rect 4200 27414 4272 27466
rect 4324 27414 4396 27466
rect 4448 27414 4520 27466
rect 4572 27414 4644 27466
rect 4696 27414 4768 27466
rect 4820 27414 4892 27466
rect 4944 27414 5016 27466
rect 5068 27414 5140 27466
rect 5192 27414 24024 27466
rect 24076 27414 24148 27466
rect 24200 27414 24272 27466
rect 24324 27414 24396 27466
rect 24448 27414 24520 27466
rect 24572 27414 24644 27466
rect 24696 27414 24768 27466
rect 24820 27414 24892 27466
rect 24944 27414 25016 27466
rect 25068 27414 25140 27466
rect 25192 27414 38640 27466
rect 1344 27380 38640 27414
rect 1710 26850 1762 26862
rect 1710 26786 1762 26798
rect 1344 26682 38640 26716
rect 1344 26630 14024 26682
rect 14076 26630 14148 26682
rect 14200 26630 14272 26682
rect 14324 26630 14396 26682
rect 14448 26630 14520 26682
rect 14572 26630 14644 26682
rect 14696 26630 14768 26682
rect 14820 26630 14892 26682
rect 14944 26630 15016 26682
rect 15068 26630 15140 26682
rect 15192 26630 34024 26682
rect 34076 26630 34148 26682
rect 34200 26630 34272 26682
rect 34324 26630 34396 26682
rect 34448 26630 34520 26682
rect 34572 26630 34644 26682
rect 34696 26630 34768 26682
rect 34820 26630 34892 26682
rect 34944 26630 35016 26682
rect 35068 26630 35140 26682
rect 35192 26630 38640 26682
rect 1344 26596 38640 26630
rect 1710 26402 1762 26414
rect 1710 26338 1762 26350
rect 1344 25898 38640 25932
rect 1344 25846 4024 25898
rect 4076 25846 4148 25898
rect 4200 25846 4272 25898
rect 4324 25846 4396 25898
rect 4448 25846 4520 25898
rect 4572 25846 4644 25898
rect 4696 25846 4768 25898
rect 4820 25846 4892 25898
rect 4944 25846 5016 25898
rect 5068 25846 5140 25898
rect 5192 25846 24024 25898
rect 24076 25846 24148 25898
rect 24200 25846 24272 25898
rect 24324 25846 24396 25898
rect 24448 25846 24520 25898
rect 24572 25846 24644 25898
rect 24696 25846 24768 25898
rect 24820 25846 24892 25898
rect 24944 25846 25016 25898
rect 25068 25846 25140 25898
rect 25192 25846 38640 25898
rect 1344 25812 38640 25846
rect 1344 25114 38640 25148
rect 1344 25062 14024 25114
rect 14076 25062 14148 25114
rect 14200 25062 14272 25114
rect 14324 25062 14396 25114
rect 14448 25062 14520 25114
rect 14572 25062 14644 25114
rect 14696 25062 14768 25114
rect 14820 25062 14892 25114
rect 14944 25062 15016 25114
rect 15068 25062 15140 25114
rect 15192 25062 34024 25114
rect 34076 25062 34148 25114
rect 34200 25062 34272 25114
rect 34324 25062 34396 25114
rect 34448 25062 34520 25114
rect 34572 25062 34644 25114
rect 34696 25062 34768 25114
rect 34820 25062 34892 25114
rect 34944 25062 35016 25114
rect 35068 25062 35140 25114
rect 35192 25062 38640 25114
rect 1344 25028 38640 25062
rect 1710 24834 1762 24846
rect 1710 24770 1762 24782
rect 1344 24330 38640 24364
rect 1344 24278 4024 24330
rect 4076 24278 4148 24330
rect 4200 24278 4272 24330
rect 4324 24278 4396 24330
rect 4448 24278 4520 24330
rect 4572 24278 4644 24330
rect 4696 24278 4768 24330
rect 4820 24278 4892 24330
rect 4944 24278 5016 24330
rect 5068 24278 5140 24330
rect 5192 24278 24024 24330
rect 24076 24278 24148 24330
rect 24200 24278 24272 24330
rect 24324 24278 24396 24330
rect 24448 24278 24520 24330
rect 24572 24278 24644 24330
rect 24696 24278 24768 24330
rect 24820 24278 24892 24330
rect 24944 24278 25016 24330
rect 25068 24278 25140 24330
rect 25192 24278 38640 24330
rect 1344 24244 38640 24278
rect 1344 23546 38640 23580
rect 1344 23494 14024 23546
rect 14076 23494 14148 23546
rect 14200 23494 14272 23546
rect 14324 23494 14396 23546
rect 14448 23494 14520 23546
rect 14572 23494 14644 23546
rect 14696 23494 14768 23546
rect 14820 23494 14892 23546
rect 14944 23494 15016 23546
rect 15068 23494 15140 23546
rect 15192 23494 34024 23546
rect 34076 23494 34148 23546
rect 34200 23494 34272 23546
rect 34324 23494 34396 23546
rect 34448 23494 34520 23546
rect 34572 23494 34644 23546
rect 34696 23494 34768 23546
rect 34820 23494 34892 23546
rect 34944 23494 35016 23546
rect 35068 23494 35140 23546
rect 35192 23494 38640 23546
rect 1344 23460 38640 23494
rect 1710 23266 1762 23278
rect 1710 23202 1762 23214
rect 1344 22762 38640 22796
rect 1344 22710 4024 22762
rect 4076 22710 4148 22762
rect 4200 22710 4272 22762
rect 4324 22710 4396 22762
rect 4448 22710 4520 22762
rect 4572 22710 4644 22762
rect 4696 22710 4768 22762
rect 4820 22710 4892 22762
rect 4944 22710 5016 22762
rect 5068 22710 5140 22762
rect 5192 22710 24024 22762
rect 24076 22710 24148 22762
rect 24200 22710 24272 22762
rect 24324 22710 24396 22762
rect 24448 22710 24520 22762
rect 24572 22710 24644 22762
rect 24696 22710 24768 22762
rect 24820 22710 24892 22762
rect 24944 22710 25016 22762
rect 25068 22710 25140 22762
rect 25192 22710 38640 22762
rect 1344 22676 38640 22710
rect 1710 22146 1762 22158
rect 1710 22082 1762 22094
rect 1344 21978 38640 22012
rect 1344 21926 14024 21978
rect 14076 21926 14148 21978
rect 14200 21926 14272 21978
rect 14324 21926 14396 21978
rect 14448 21926 14520 21978
rect 14572 21926 14644 21978
rect 14696 21926 14768 21978
rect 14820 21926 14892 21978
rect 14944 21926 15016 21978
rect 15068 21926 15140 21978
rect 15192 21926 34024 21978
rect 34076 21926 34148 21978
rect 34200 21926 34272 21978
rect 34324 21926 34396 21978
rect 34448 21926 34520 21978
rect 34572 21926 34644 21978
rect 34696 21926 34768 21978
rect 34820 21926 34892 21978
rect 34944 21926 35016 21978
rect 35068 21926 35140 21978
rect 35192 21926 38640 21978
rect 1344 21892 38640 21926
rect 1344 21194 38640 21228
rect 1344 21142 4024 21194
rect 4076 21142 4148 21194
rect 4200 21142 4272 21194
rect 4324 21142 4396 21194
rect 4448 21142 4520 21194
rect 4572 21142 4644 21194
rect 4696 21142 4768 21194
rect 4820 21142 4892 21194
rect 4944 21142 5016 21194
rect 5068 21142 5140 21194
rect 5192 21142 24024 21194
rect 24076 21142 24148 21194
rect 24200 21142 24272 21194
rect 24324 21142 24396 21194
rect 24448 21142 24520 21194
rect 24572 21142 24644 21194
rect 24696 21142 24768 21194
rect 24820 21142 24892 21194
rect 24944 21142 25016 21194
rect 25068 21142 25140 21194
rect 25192 21142 38640 21194
rect 1344 21108 38640 21142
rect 1710 20578 1762 20590
rect 1710 20514 1762 20526
rect 1344 20410 38640 20444
rect 1344 20358 14024 20410
rect 14076 20358 14148 20410
rect 14200 20358 14272 20410
rect 14324 20358 14396 20410
rect 14448 20358 14520 20410
rect 14572 20358 14644 20410
rect 14696 20358 14768 20410
rect 14820 20358 14892 20410
rect 14944 20358 15016 20410
rect 15068 20358 15140 20410
rect 15192 20358 34024 20410
rect 34076 20358 34148 20410
rect 34200 20358 34272 20410
rect 34324 20358 34396 20410
rect 34448 20358 34520 20410
rect 34572 20358 34644 20410
rect 34696 20358 34768 20410
rect 34820 20358 34892 20410
rect 34944 20358 35016 20410
rect 35068 20358 35140 20410
rect 35192 20358 38640 20410
rect 1344 20324 38640 20358
rect 1344 19626 38640 19660
rect 1344 19574 4024 19626
rect 4076 19574 4148 19626
rect 4200 19574 4272 19626
rect 4324 19574 4396 19626
rect 4448 19574 4520 19626
rect 4572 19574 4644 19626
rect 4696 19574 4768 19626
rect 4820 19574 4892 19626
rect 4944 19574 5016 19626
rect 5068 19574 5140 19626
rect 5192 19574 24024 19626
rect 24076 19574 24148 19626
rect 24200 19574 24272 19626
rect 24324 19574 24396 19626
rect 24448 19574 24520 19626
rect 24572 19574 24644 19626
rect 24696 19574 24768 19626
rect 24820 19574 24892 19626
rect 24944 19574 25016 19626
rect 25068 19574 25140 19626
rect 25192 19574 38640 19626
rect 1344 19540 38640 19574
rect 1710 19010 1762 19022
rect 1710 18946 1762 18958
rect 38222 19010 38274 19022
rect 38222 18946 38274 18958
rect 1344 18842 38640 18876
rect 1344 18790 14024 18842
rect 14076 18790 14148 18842
rect 14200 18790 14272 18842
rect 14324 18790 14396 18842
rect 14448 18790 14520 18842
rect 14572 18790 14644 18842
rect 14696 18790 14768 18842
rect 14820 18790 14892 18842
rect 14944 18790 15016 18842
rect 15068 18790 15140 18842
rect 15192 18790 34024 18842
rect 34076 18790 34148 18842
rect 34200 18790 34272 18842
rect 34324 18790 34396 18842
rect 34448 18790 34520 18842
rect 34572 18790 34644 18842
rect 34696 18790 34768 18842
rect 34820 18790 34892 18842
rect 34944 18790 35016 18842
rect 35068 18790 35140 18842
rect 35192 18790 38640 18842
rect 1344 18756 38640 18790
rect 1344 18058 38640 18092
rect 1344 18006 4024 18058
rect 4076 18006 4148 18058
rect 4200 18006 4272 18058
rect 4324 18006 4396 18058
rect 4448 18006 4520 18058
rect 4572 18006 4644 18058
rect 4696 18006 4768 18058
rect 4820 18006 4892 18058
rect 4944 18006 5016 18058
rect 5068 18006 5140 18058
rect 5192 18006 24024 18058
rect 24076 18006 24148 18058
rect 24200 18006 24272 18058
rect 24324 18006 24396 18058
rect 24448 18006 24520 18058
rect 24572 18006 24644 18058
rect 24696 18006 24768 18058
rect 24820 18006 24892 18058
rect 24944 18006 25016 18058
rect 25068 18006 25140 18058
rect 25192 18006 38640 18058
rect 1344 17972 38640 18006
rect 1710 17554 1762 17566
rect 1710 17490 1762 17502
rect 1344 17274 38640 17308
rect 1344 17222 14024 17274
rect 14076 17222 14148 17274
rect 14200 17222 14272 17274
rect 14324 17222 14396 17274
rect 14448 17222 14520 17274
rect 14572 17222 14644 17274
rect 14696 17222 14768 17274
rect 14820 17222 14892 17274
rect 14944 17222 15016 17274
rect 15068 17222 15140 17274
rect 15192 17222 34024 17274
rect 34076 17222 34148 17274
rect 34200 17222 34272 17274
rect 34324 17222 34396 17274
rect 34448 17222 34520 17274
rect 34572 17222 34644 17274
rect 34696 17222 34768 17274
rect 34820 17222 34892 17274
rect 34944 17222 35016 17274
rect 35068 17222 35140 17274
rect 35192 17222 38640 17274
rect 1344 17188 38640 17222
rect 1710 16994 1762 17006
rect 1710 16930 1762 16942
rect 1344 16490 38640 16524
rect 1344 16438 4024 16490
rect 4076 16438 4148 16490
rect 4200 16438 4272 16490
rect 4324 16438 4396 16490
rect 4448 16438 4520 16490
rect 4572 16438 4644 16490
rect 4696 16438 4768 16490
rect 4820 16438 4892 16490
rect 4944 16438 5016 16490
rect 5068 16438 5140 16490
rect 5192 16438 24024 16490
rect 24076 16438 24148 16490
rect 24200 16438 24272 16490
rect 24324 16438 24396 16490
rect 24448 16438 24520 16490
rect 24572 16438 24644 16490
rect 24696 16438 24768 16490
rect 24820 16438 24892 16490
rect 24944 16438 25016 16490
rect 25068 16438 25140 16490
rect 25192 16438 38640 16490
rect 1344 16404 38640 16438
rect 1344 15706 38640 15740
rect 1344 15654 14024 15706
rect 14076 15654 14148 15706
rect 14200 15654 14272 15706
rect 14324 15654 14396 15706
rect 14448 15654 14520 15706
rect 14572 15654 14644 15706
rect 14696 15654 14768 15706
rect 14820 15654 14892 15706
rect 14944 15654 15016 15706
rect 15068 15654 15140 15706
rect 15192 15654 34024 15706
rect 34076 15654 34148 15706
rect 34200 15654 34272 15706
rect 34324 15654 34396 15706
rect 34448 15654 34520 15706
rect 34572 15654 34644 15706
rect 34696 15654 34768 15706
rect 34820 15654 34892 15706
rect 34944 15654 35016 15706
rect 35068 15654 35140 15706
rect 35192 15654 38640 15706
rect 1344 15620 38640 15654
rect 1710 15426 1762 15438
rect 1710 15362 1762 15374
rect 1344 14922 38640 14956
rect 1344 14870 4024 14922
rect 4076 14870 4148 14922
rect 4200 14870 4272 14922
rect 4324 14870 4396 14922
rect 4448 14870 4520 14922
rect 4572 14870 4644 14922
rect 4696 14870 4768 14922
rect 4820 14870 4892 14922
rect 4944 14870 5016 14922
rect 5068 14870 5140 14922
rect 5192 14870 24024 14922
rect 24076 14870 24148 14922
rect 24200 14870 24272 14922
rect 24324 14870 24396 14922
rect 24448 14870 24520 14922
rect 24572 14870 24644 14922
rect 24696 14870 24768 14922
rect 24820 14870 24892 14922
rect 24944 14870 25016 14922
rect 25068 14870 25140 14922
rect 25192 14870 38640 14922
rect 1344 14836 38640 14870
rect 1344 14138 38640 14172
rect 1344 14086 14024 14138
rect 14076 14086 14148 14138
rect 14200 14086 14272 14138
rect 14324 14086 14396 14138
rect 14448 14086 14520 14138
rect 14572 14086 14644 14138
rect 14696 14086 14768 14138
rect 14820 14086 14892 14138
rect 14944 14086 15016 14138
rect 15068 14086 15140 14138
rect 15192 14086 34024 14138
rect 34076 14086 34148 14138
rect 34200 14086 34272 14138
rect 34324 14086 34396 14138
rect 34448 14086 34520 14138
rect 34572 14086 34644 14138
rect 34696 14086 34768 14138
rect 34820 14086 34892 14138
rect 34944 14086 35016 14138
rect 35068 14086 35140 14138
rect 35192 14086 38640 14138
rect 1344 14052 38640 14086
rect 1710 13858 1762 13870
rect 1710 13794 1762 13806
rect 1344 13354 38640 13388
rect 1344 13302 4024 13354
rect 4076 13302 4148 13354
rect 4200 13302 4272 13354
rect 4324 13302 4396 13354
rect 4448 13302 4520 13354
rect 4572 13302 4644 13354
rect 4696 13302 4768 13354
rect 4820 13302 4892 13354
rect 4944 13302 5016 13354
rect 5068 13302 5140 13354
rect 5192 13302 24024 13354
rect 24076 13302 24148 13354
rect 24200 13302 24272 13354
rect 24324 13302 24396 13354
rect 24448 13302 24520 13354
rect 24572 13302 24644 13354
rect 24696 13302 24768 13354
rect 24820 13302 24892 13354
rect 24944 13302 25016 13354
rect 25068 13302 25140 13354
rect 25192 13302 38640 13354
rect 1344 13268 38640 13302
rect 1710 12738 1762 12750
rect 1710 12674 1762 12686
rect 1344 12570 38640 12604
rect 1344 12518 14024 12570
rect 14076 12518 14148 12570
rect 14200 12518 14272 12570
rect 14324 12518 14396 12570
rect 14448 12518 14520 12570
rect 14572 12518 14644 12570
rect 14696 12518 14768 12570
rect 14820 12518 14892 12570
rect 14944 12518 15016 12570
rect 15068 12518 15140 12570
rect 15192 12518 34024 12570
rect 34076 12518 34148 12570
rect 34200 12518 34272 12570
rect 34324 12518 34396 12570
rect 34448 12518 34520 12570
rect 34572 12518 34644 12570
rect 34696 12518 34768 12570
rect 34820 12518 34892 12570
rect 34944 12518 35016 12570
rect 35068 12518 35140 12570
rect 35192 12518 38640 12570
rect 1344 12484 38640 12518
rect 1344 11786 38640 11820
rect 1344 11734 4024 11786
rect 4076 11734 4148 11786
rect 4200 11734 4272 11786
rect 4324 11734 4396 11786
rect 4448 11734 4520 11786
rect 4572 11734 4644 11786
rect 4696 11734 4768 11786
rect 4820 11734 4892 11786
rect 4944 11734 5016 11786
rect 5068 11734 5140 11786
rect 5192 11734 24024 11786
rect 24076 11734 24148 11786
rect 24200 11734 24272 11786
rect 24324 11734 24396 11786
rect 24448 11734 24520 11786
rect 24572 11734 24644 11786
rect 24696 11734 24768 11786
rect 24820 11734 24892 11786
rect 24944 11734 25016 11786
rect 25068 11734 25140 11786
rect 25192 11734 38640 11786
rect 1344 11700 38640 11734
rect 1710 11170 1762 11182
rect 1710 11106 1762 11118
rect 1344 11002 38640 11036
rect 1344 10950 14024 11002
rect 14076 10950 14148 11002
rect 14200 10950 14272 11002
rect 14324 10950 14396 11002
rect 14448 10950 14520 11002
rect 14572 10950 14644 11002
rect 14696 10950 14768 11002
rect 14820 10950 14892 11002
rect 14944 10950 15016 11002
rect 15068 10950 15140 11002
rect 15192 10950 34024 11002
rect 34076 10950 34148 11002
rect 34200 10950 34272 11002
rect 34324 10950 34396 11002
rect 34448 10950 34520 11002
rect 34572 10950 34644 11002
rect 34696 10950 34768 11002
rect 34820 10950 34892 11002
rect 34944 10950 35016 11002
rect 35068 10950 35140 11002
rect 35192 10950 38640 11002
rect 1344 10916 38640 10950
rect 11902 10610 11954 10622
rect 11902 10546 11954 10558
rect 12126 10610 12178 10622
rect 12126 10546 12178 10558
rect 12574 10610 12626 10622
rect 12574 10546 12626 10558
rect 12910 10610 12962 10622
rect 12910 10546 12962 10558
rect 12014 10498 12066 10510
rect 12014 10434 12066 10446
rect 13358 10498 13410 10510
rect 13358 10434 13410 10446
rect 12674 10334 12686 10386
rect 12738 10383 12750 10386
rect 13346 10383 13358 10386
rect 12738 10337 13358 10383
rect 12738 10334 12750 10337
rect 13346 10334 13358 10337
rect 13410 10334 13422 10386
rect 1344 10218 38640 10252
rect 1344 10166 4024 10218
rect 4076 10166 4148 10218
rect 4200 10166 4272 10218
rect 4324 10166 4396 10218
rect 4448 10166 4520 10218
rect 4572 10166 4644 10218
rect 4696 10166 4768 10218
rect 4820 10166 4892 10218
rect 4944 10166 5016 10218
rect 5068 10166 5140 10218
rect 5192 10166 24024 10218
rect 24076 10166 24148 10218
rect 24200 10166 24272 10218
rect 24324 10166 24396 10218
rect 24448 10166 24520 10218
rect 24572 10166 24644 10218
rect 24696 10166 24768 10218
rect 24820 10166 24892 10218
rect 24944 10166 25016 10218
rect 25068 10166 25140 10218
rect 25192 10166 38640 10218
rect 1344 10132 38640 10166
rect 12686 9938 12738 9950
rect 12686 9874 12738 9886
rect 9762 9774 9774 9826
rect 9826 9774 9838 9826
rect 7758 9714 7810 9726
rect 7758 9650 7810 9662
rect 8318 9714 8370 9726
rect 10546 9662 10558 9714
rect 10610 9662 10622 9714
rect 8318 9650 8370 9662
rect 1710 9602 1762 9614
rect 1710 9538 1762 9550
rect 7646 9602 7698 9614
rect 7646 9538 7698 9550
rect 13694 9602 13746 9614
rect 13694 9538 13746 9550
rect 1344 9434 38640 9468
rect 1344 9382 14024 9434
rect 14076 9382 14148 9434
rect 14200 9382 14272 9434
rect 14324 9382 14396 9434
rect 14448 9382 14520 9434
rect 14572 9382 14644 9434
rect 14696 9382 14768 9434
rect 14820 9382 14892 9434
rect 14944 9382 15016 9434
rect 15068 9382 15140 9434
rect 15192 9382 34024 9434
rect 34076 9382 34148 9434
rect 34200 9382 34272 9434
rect 34324 9382 34396 9434
rect 34448 9382 34520 9434
rect 34572 9382 34644 9434
rect 34696 9382 34768 9434
rect 34820 9382 34892 9434
rect 34944 9382 35016 9434
rect 35068 9382 35140 9434
rect 35192 9382 38640 9434
rect 1344 9348 38640 9382
rect 10446 9266 10498 9278
rect 10446 9202 10498 9214
rect 10782 9154 10834 9166
rect 10782 9090 10834 9102
rect 10222 9042 10274 9054
rect 10222 8978 10274 8990
rect 10446 9042 10498 9054
rect 11330 8990 11342 9042
rect 11394 8990 11406 9042
rect 10446 8978 10498 8990
rect 6414 8930 6466 8942
rect 6414 8866 6466 8878
rect 7422 8930 7474 8942
rect 7422 8866 7474 8878
rect 7870 8930 7922 8942
rect 7870 8866 7922 8878
rect 8430 8930 8482 8942
rect 8430 8866 8482 8878
rect 8766 8930 8818 8942
rect 8766 8866 8818 8878
rect 9662 8930 9714 8942
rect 13458 8878 13470 8930
rect 13522 8878 13534 8930
rect 9662 8866 9714 8878
rect 1344 8650 38640 8684
rect 1344 8598 4024 8650
rect 4076 8598 4148 8650
rect 4200 8598 4272 8650
rect 4324 8598 4396 8650
rect 4448 8598 4520 8650
rect 4572 8598 4644 8650
rect 4696 8598 4768 8650
rect 4820 8598 4892 8650
rect 4944 8598 5016 8650
rect 5068 8598 5140 8650
rect 5192 8598 24024 8650
rect 24076 8598 24148 8650
rect 24200 8598 24272 8650
rect 24324 8598 24396 8650
rect 24448 8598 24520 8650
rect 24572 8598 24644 8650
rect 24696 8598 24768 8650
rect 24820 8598 24892 8650
rect 24944 8598 25016 8650
rect 25068 8598 25140 8650
rect 25192 8598 38640 8650
rect 1344 8564 38640 8598
rect 7422 8370 7474 8382
rect 7422 8306 7474 8318
rect 7758 8370 7810 8382
rect 7758 8306 7810 8318
rect 5966 8258 6018 8270
rect 5966 8194 6018 8206
rect 10782 8258 10834 8270
rect 10782 8194 10834 8206
rect 12798 8258 12850 8270
rect 13458 8206 13470 8258
rect 13522 8206 13534 8258
rect 12798 8194 12850 8206
rect 1710 8146 1762 8158
rect 1710 8082 1762 8094
rect 5630 8146 5682 8158
rect 5630 8082 5682 8094
rect 8206 8146 8258 8158
rect 8206 8082 8258 8094
rect 8318 8146 8370 8158
rect 8318 8082 8370 8094
rect 9662 8146 9714 8158
rect 12898 8094 12910 8146
rect 12962 8094 12974 8146
rect 14242 8094 14254 8146
rect 14306 8094 14318 8146
rect 9662 8082 9714 8094
rect 3054 8034 3106 8046
rect 3054 7970 3106 7982
rect 3390 8034 3442 8046
rect 3390 7970 3442 7982
rect 3950 8034 4002 8046
rect 3950 7970 4002 7982
rect 4622 8034 4674 8046
rect 4622 7970 4674 7982
rect 5182 8034 5234 8046
rect 5182 7970 5234 7982
rect 5742 8034 5794 8046
rect 5742 7970 5794 7982
rect 6526 8034 6578 8046
rect 6526 7970 6578 7982
rect 6974 8034 7026 8046
rect 6974 7970 7026 7982
rect 7646 8034 7698 8046
rect 7646 7970 7698 7982
rect 7982 8034 8034 8046
rect 7982 7970 8034 7982
rect 8766 8034 8818 8046
rect 9202 7982 9214 8034
rect 9266 7982 9278 8034
rect 16482 7982 16494 8034
rect 16546 7982 16558 8034
rect 8766 7970 8818 7982
rect 1344 7866 38640 7900
rect 1344 7814 14024 7866
rect 14076 7814 14148 7866
rect 14200 7814 14272 7866
rect 14324 7814 14396 7866
rect 14448 7814 14520 7866
rect 14572 7814 14644 7866
rect 14696 7814 14768 7866
rect 14820 7814 14892 7866
rect 14944 7814 15016 7866
rect 15068 7814 15140 7866
rect 15192 7814 34024 7866
rect 34076 7814 34148 7866
rect 34200 7814 34272 7866
rect 34324 7814 34396 7866
rect 34448 7814 34520 7866
rect 34572 7814 34644 7866
rect 34696 7814 34768 7866
rect 34820 7814 34892 7866
rect 34944 7814 35016 7866
rect 35068 7814 35140 7866
rect 35192 7814 38640 7866
rect 1344 7780 38640 7814
rect 8878 7698 8930 7710
rect 8878 7634 8930 7646
rect 8990 7586 9042 7598
rect 13134 7586 13186 7598
rect 10098 7534 10110 7586
rect 10162 7534 10174 7586
rect 8990 7522 9042 7534
rect 13134 7522 13186 7534
rect 7534 7474 7586 7486
rect 2930 7422 2942 7474
rect 2994 7422 3006 7474
rect 7186 7422 7198 7474
rect 7250 7422 7262 7474
rect 7534 7410 7586 7422
rect 7758 7474 7810 7486
rect 7758 7410 7810 7422
rect 8206 7474 8258 7486
rect 8206 7410 8258 7422
rect 8654 7474 8706 7486
rect 8654 7410 8706 7422
rect 11678 7474 11730 7486
rect 11678 7410 11730 7422
rect 13694 7474 13746 7486
rect 13694 7410 13746 7422
rect 14702 7474 14754 7486
rect 14702 7410 14754 7422
rect 3502 7362 3554 7374
rect 1922 7310 1934 7362
rect 1986 7310 1998 7362
rect 3502 7298 3554 7310
rect 3950 7362 4002 7374
rect 7982 7362 8034 7374
rect 4274 7310 4286 7362
rect 4338 7310 4350 7362
rect 6402 7310 6414 7362
rect 6466 7310 6478 7362
rect 3950 7298 4002 7310
rect 7982 7298 8034 7310
rect 9774 7362 9826 7374
rect 9774 7298 9826 7310
rect 11790 7362 11842 7374
rect 11790 7298 11842 7310
rect 14254 7362 14306 7374
rect 14254 7298 14306 7310
rect 15150 7362 15202 7374
rect 15150 7298 15202 7310
rect 15598 7362 15650 7374
rect 15598 7298 15650 7310
rect 3490 7198 3502 7250
rect 3554 7247 3566 7250
rect 3938 7247 3950 7250
rect 3554 7201 3950 7247
rect 3554 7198 3566 7201
rect 3938 7198 3950 7201
rect 4002 7198 4014 7250
rect 14018 7198 14030 7250
rect 14082 7247 14094 7250
rect 14242 7247 14254 7250
rect 14082 7201 14254 7247
rect 14082 7198 14094 7201
rect 14242 7198 14254 7201
rect 14306 7247 14318 7250
rect 15586 7247 15598 7250
rect 14306 7201 15598 7247
rect 14306 7198 14318 7201
rect 15586 7198 15598 7201
rect 15650 7198 15662 7250
rect 1344 7082 38640 7116
rect 1344 7030 4024 7082
rect 4076 7030 4148 7082
rect 4200 7030 4272 7082
rect 4324 7030 4396 7082
rect 4448 7030 4520 7082
rect 4572 7030 4644 7082
rect 4696 7030 4768 7082
rect 4820 7030 4892 7082
rect 4944 7030 5016 7082
rect 5068 7030 5140 7082
rect 5192 7030 24024 7082
rect 24076 7030 24148 7082
rect 24200 7030 24272 7082
rect 24324 7030 24396 7082
rect 24448 7030 24520 7082
rect 24572 7030 24644 7082
rect 24696 7030 24768 7082
rect 24820 7030 24892 7082
rect 24944 7030 25016 7082
rect 25068 7030 25140 7082
rect 25192 7030 38640 7082
rect 1344 6996 38640 7030
rect 7198 6802 7250 6814
rect 1810 6750 1822 6802
rect 1874 6750 1886 6802
rect 17602 6750 17614 6802
rect 17666 6750 17678 6802
rect 7198 6738 7250 6750
rect 6526 6690 6578 6702
rect 21422 6690 21474 6702
rect 4722 6638 4734 6690
rect 4786 6638 4798 6690
rect 6738 6638 6750 6690
rect 6802 6638 6814 6690
rect 10210 6638 10222 6690
rect 10274 6638 10286 6690
rect 10658 6638 10670 6690
rect 10722 6638 10734 6690
rect 13458 6638 13470 6690
rect 13522 6638 13534 6690
rect 15474 6638 15486 6690
rect 15538 6638 15550 6690
rect 20514 6638 20526 6690
rect 20578 6638 20590 6690
rect 6526 6626 6578 6638
rect 21422 6626 21474 6638
rect 5742 6578 5794 6590
rect 3938 6526 3950 6578
rect 4002 6526 4014 6578
rect 5742 6514 5794 6526
rect 5854 6578 5906 6590
rect 7310 6578 7362 6590
rect 11230 6578 11282 6590
rect 16046 6578 16098 6590
rect 37886 6578 37938 6590
rect 5854 6514 5906 6526
rect 6190 6522 6242 6534
rect 5518 6466 5570 6478
rect 8642 6526 8654 6578
rect 8706 6526 8718 6578
rect 13570 6526 13582 6578
rect 13634 6526 13646 6578
rect 19730 6526 19742 6578
rect 19794 6526 19806 6578
rect 7310 6514 7362 6526
rect 11230 6514 11282 6526
rect 16046 6514 16098 6526
rect 37886 6514 37938 6526
rect 38222 6578 38274 6590
rect 38222 6514 38274 6526
rect 6190 6458 6242 6470
rect 6302 6466 6354 6478
rect 5518 6402 5570 6414
rect 6302 6402 6354 6414
rect 7086 6466 7138 6478
rect 7086 6402 7138 6414
rect 7758 6466 7810 6478
rect 7758 6402 7810 6414
rect 7870 6466 7922 6478
rect 7870 6402 7922 6414
rect 7982 6466 8034 6478
rect 7982 6402 8034 6414
rect 8206 6466 8258 6478
rect 8206 6402 8258 6414
rect 11118 6466 11170 6478
rect 11118 6402 11170 6414
rect 13022 6466 13074 6478
rect 37662 6466 37714 6478
rect 15474 6414 15486 6466
rect 15538 6414 15550 6466
rect 13022 6402 13074 6414
rect 37662 6402 37714 6414
rect 1344 6298 38640 6332
rect 1344 6246 14024 6298
rect 14076 6246 14148 6298
rect 14200 6246 14272 6298
rect 14324 6246 14396 6298
rect 14448 6246 14520 6298
rect 14572 6246 14644 6298
rect 14696 6246 14768 6298
rect 14820 6246 14892 6298
rect 14944 6246 15016 6298
rect 15068 6246 15140 6298
rect 15192 6246 34024 6298
rect 34076 6246 34148 6298
rect 34200 6246 34272 6298
rect 34324 6246 34396 6298
rect 34448 6246 34520 6298
rect 34572 6246 34644 6298
rect 34696 6246 34768 6298
rect 34820 6246 34892 6298
rect 34944 6246 35016 6298
rect 35068 6246 35140 6298
rect 35192 6246 38640 6298
rect 1344 6212 38640 6246
rect 6862 6130 6914 6142
rect 6862 6066 6914 6078
rect 20750 6130 20802 6142
rect 20750 6066 20802 6078
rect 2270 6018 2322 6030
rect 2270 5954 2322 5966
rect 5966 6018 6018 6030
rect 5966 5954 6018 5966
rect 6526 6018 6578 6030
rect 7646 6018 7698 6030
rect 7410 5966 7422 6018
rect 7474 5966 7486 6018
rect 6526 5954 6578 5966
rect 7646 5954 7698 5966
rect 8094 6018 8146 6030
rect 8094 5954 8146 5966
rect 8990 6018 9042 6030
rect 11330 5966 11342 6018
rect 11394 5966 11406 6018
rect 8990 5954 9042 5966
rect 6302 5906 6354 5918
rect 8542 5906 8594 5918
rect 1922 5854 1934 5906
rect 1986 5854 1998 5906
rect 5506 5854 5518 5906
rect 5570 5854 5582 5906
rect 6962 5854 6974 5906
rect 7026 5854 7038 5906
rect 6302 5842 6354 5854
rect 8542 5842 8594 5854
rect 8654 5906 8706 5918
rect 15374 5906 15426 5918
rect 14802 5854 14814 5906
rect 14866 5854 14878 5906
rect 8654 5842 8706 5854
rect 15374 5842 15426 5854
rect 6078 5794 6130 5806
rect 2034 5742 2046 5794
rect 2098 5742 2110 5794
rect 2594 5742 2606 5794
rect 2658 5742 2670 5794
rect 4722 5742 4734 5794
rect 4786 5742 4798 5794
rect 6078 5730 6130 5742
rect 7982 5794 8034 5806
rect 7982 5730 8034 5742
rect 8878 5794 8930 5806
rect 8878 5730 8930 5742
rect 15822 5794 15874 5806
rect 15822 5730 15874 5742
rect 16158 5794 16210 5806
rect 16158 5730 16210 5742
rect 16830 5794 16882 5806
rect 16830 5730 16882 5742
rect 17502 5794 17554 5806
rect 17502 5730 17554 5742
rect 17950 5794 18002 5806
rect 17950 5730 18002 5742
rect 24334 5794 24386 5806
rect 24334 5730 24386 5742
rect 7074 5630 7086 5682
rect 7138 5630 7150 5682
rect 1344 5514 38640 5548
rect 1344 5462 4024 5514
rect 4076 5462 4148 5514
rect 4200 5462 4272 5514
rect 4324 5462 4396 5514
rect 4448 5462 4520 5514
rect 4572 5462 4644 5514
rect 4696 5462 4768 5514
rect 4820 5462 4892 5514
rect 4944 5462 5016 5514
rect 5068 5462 5140 5514
rect 5192 5462 24024 5514
rect 24076 5462 24148 5514
rect 24200 5462 24272 5514
rect 24324 5462 24396 5514
rect 24448 5462 24520 5514
rect 24572 5462 24644 5514
rect 24696 5462 24768 5514
rect 24820 5462 24892 5514
rect 24944 5462 25016 5514
rect 25068 5462 25140 5514
rect 25192 5462 38640 5514
rect 1344 5428 38640 5462
rect 2158 5346 2210 5358
rect 2158 5282 2210 5294
rect 11566 5234 11618 5246
rect 6066 5182 6078 5234
rect 6130 5182 6142 5234
rect 11566 5170 11618 5182
rect 3390 5122 3442 5134
rect 2818 5070 2830 5122
rect 2882 5070 2894 5122
rect 3390 5058 3442 5070
rect 4062 5122 4114 5134
rect 12126 5122 12178 5134
rect 11106 5070 11118 5122
rect 11170 5070 11182 5122
rect 4062 5058 4114 5070
rect 12126 5058 12178 5070
rect 12238 5122 12290 5134
rect 28142 5122 28194 5134
rect 32286 5122 32338 5134
rect 13794 5070 13806 5122
rect 13858 5070 13870 5122
rect 14354 5070 14366 5122
rect 14418 5070 14430 5122
rect 16594 5070 16606 5122
rect 16658 5070 16670 5122
rect 22194 5070 22206 5122
rect 22258 5070 22270 5122
rect 26002 5070 26014 5122
rect 26066 5070 26078 5122
rect 30146 5070 30158 5122
rect 30210 5070 30222 5122
rect 12238 5058 12290 5070
rect 28142 5058 28194 5070
rect 32286 5058 32338 5070
rect 34974 5122 35026 5134
rect 34974 5058 35026 5070
rect 4398 5010 4450 5022
rect 3714 4958 3726 5010
rect 3778 4958 3790 5010
rect 4398 4946 4450 4958
rect 5070 5010 5122 5022
rect 5070 4946 5122 4958
rect 11678 5010 11730 5022
rect 11678 4946 11730 4958
rect 12574 5010 12626 5022
rect 12574 4946 12626 4958
rect 14030 5010 14082 5022
rect 14030 4946 14082 4958
rect 15598 5010 15650 5022
rect 15598 4946 15650 4958
rect 17054 5010 17106 5022
rect 17054 4946 17106 4958
rect 22878 5010 22930 5022
rect 22878 4946 22930 4958
rect 24894 5010 24946 5022
rect 32846 5010 32898 5022
rect 30258 4958 30270 5010
rect 30322 4958 30334 5010
rect 24894 4946 24946 4958
rect 32846 4946 32898 4958
rect 1710 4898 1762 4910
rect 1710 4834 1762 4846
rect 4846 4898 4898 4910
rect 4846 4834 4898 4846
rect 4958 4898 5010 4910
rect 4958 4834 5010 4846
rect 11454 4898 11506 4910
rect 11454 4834 11506 4846
rect 12462 4898 12514 4910
rect 12462 4834 12514 4846
rect 15150 4898 15202 4910
rect 15150 4834 15202 4846
rect 18734 4898 18786 4910
rect 18734 4834 18786 4846
rect 19518 4898 19570 4910
rect 19518 4834 19570 4846
rect 20526 4898 20578 4910
rect 20526 4834 20578 4846
rect 21534 4898 21586 4910
rect 21534 4834 21586 4846
rect 21982 4898 22034 4910
rect 21982 4834 22034 4846
rect 23774 4898 23826 4910
rect 23774 4834 23826 4846
rect 26462 4898 26514 4910
rect 26462 4834 26514 4846
rect 26910 4898 26962 4910
rect 34414 4898 34466 4910
rect 33842 4846 33854 4898
rect 33906 4846 33918 4898
rect 26910 4834 26962 4846
rect 34414 4834 34466 4846
rect 1344 4730 38640 4764
rect 1344 4678 14024 4730
rect 14076 4678 14148 4730
rect 14200 4678 14272 4730
rect 14324 4678 14396 4730
rect 14448 4678 14520 4730
rect 14572 4678 14644 4730
rect 14696 4678 14768 4730
rect 14820 4678 14892 4730
rect 14944 4678 15016 4730
rect 15068 4678 15140 4730
rect 15192 4678 34024 4730
rect 34076 4678 34148 4730
rect 34200 4678 34272 4730
rect 34324 4678 34396 4730
rect 34448 4678 34520 4730
rect 34572 4678 34644 4730
rect 34696 4678 34768 4730
rect 34820 4678 34892 4730
rect 34944 4678 35016 4730
rect 35068 4678 35140 4730
rect 35192 4678 38640 4730
rect 1344 4644 38640 4678
rect 6862 4562 6914 4574
rect 6862 4498 6914 4510
rect 8206 4562 8258 4574
rect 11118 4562 11170 4574
rect 16382 4562 16434 4574
rect 8978 4510 8990 4562
rect 9042 4510 9054 4562
rect 9874 4510 9886 4562
rect 9938 4510 9950 4562
rect 11666 4510 11678 4562
rect 11730 4510 11742 4562
rect 25330 4510 25342 4562
rect 25394 4510 25406 4562
rect 8206 4498 8258 4510
rect 11118 4498 11170 4510
rect 16382 4498 16434 4510
rect 7646 4450 7698 4462
rect 3826 4398 3838 4450
rect 3890 4398 3902 4450
rect 5394 4398 5406 4450
rect 5458 4398 5470 4450
rect 6066 4398 6078 4450
rect 6130 4398 6142 4450
rect 7410 4398 7422 4450
rect 7474 4398 7486 4450
rect 7646 4386 7698 4398
rect 8094 4450 8146 4462
rect 8094 4386 8146 4398
rect 12126 4450 12178 4462
rect 12126 4386 12178 4398
rect 14702 4450 14754 4462
rect 19406 4450 19458 4462
rect 17378 4398 17390 4450
rect 17442 4398 17454 4450
rect 14702 4386 14754 4398
rect 19406 4386 19458 4398
rect 20862 4450 20914 4462
rect 25902 4450 25954 4462
rect 23762 4398 23774 4450
rect 23826 4398 23838 4450
rect 20862 4386 20914 4398
rect 25902 4386 25954 4398
rect 27918 4450 27970 4462
rect 27918 4386 27970 4398
rect 33070 4450 33122 4462
rect 33070 4386 33122 4398
rect 33742 4450 33794 4462
rect 33742 4386 33794 4398
rect 34750 4450 34802 4462
rect 34750 4386 34802 4398
rect 35086 4450 35138 4462
rect 35086 4386 35138 4398
rect 6414 4338 6466 4350
rect 7982 4338 8034 4350
rect 16046 4338 16098 4350
rect 4610 4286 4622 4338
rect 4674 4286 4686 4338
rect 5282 4286 5294 4338
rect 5346 4286 5358 4338
rect 6850 4286 6862 4338
rect 6914 4286 6926 4338
rect 8754 4286 8766 4338
rect 8818 4286 8830 4338
rect 9874 4286 9886 4338
rect 9938 4286 9950 4338
rect 10098 4286 10110 4338
rect 10162 4286 10174 4338
rect 11554 4286 11566 4338
rect 11618 4286 11630 4338
rect 13570 4286 13582 4338
rect 13634 4286 13646 4338
rect 6414 4274 6466 4286
rect 7982 4274 8034 4286
rect 16046 4274 16098 4286
rect 18286 4338 18338 4350
rect 25342 4338 25394 4350
rect 20402 4286 20414 4338
rect 20466 4286 20478 4338
rect 24098 4286 24110 4338
rect 24162 4286 24174 4338
rect 27458 4286 27470 4338
rect 27522 4286 27534 4338
rect 33282 4286 33294 4338
rect 33346 4286 33358 4338
rect 33954 4286 33966 4338
rect 34018 4286 34030 4338
rect 34402 4286 34414 4338
rect 34466 4286 34478 4338
rect 35298 4286 35310 4338
rect 35362 4286 35374 4338
rect 18286 4274 18338 4286
rect 25342 4274 25394 4286
rect 11230 4226 11282 4238
rect 1698 4174 1710 4226
rect 1762 4174 1774 4226
rect 9986 4174 9998 4226
rect 10050 4174 10062 4226
rect 11230 4162 11282 4174
rect 16942 4226 16994 4238
rect 16942 4162 16994 4174
rect 17726 4226 17778 4238
rect 24558 4226 24610 4238
rect 18610 4174 18622 4226
rect 18674 4174 18686 4226
rect 17726 4162 17778 4174
rect 24558 4162 24610 4174
rect 29486 4226 29538 4238
rect 29486 4162 29538 4174
rect 29934 4226 29986 4238
rect 30494 4226 30546 4238
rect 30146 4174 30158 4226
rect 30210 4174 30222 4226
rect 29934 4162 29986 4174
rect 7074 4062 7086 4114
rect 7138 4062 7150 4114
rect 22754 4062 22766 4114
rect 22818 4062 22830 4114
rect 29362 4062 29374 4114
rect 29426 4111 29438 4114
rect 30161 4111 30207 4174
rect 30494 4162 30546 4174
rect 31838 4226 31890 4238
rect 31838 4162 31890 4174
rect 32510 4226 32562 4238
rect 32510 4162 32562 4174
rect 35982 4226 36034 4238
rect 35982 4162 36034 4174
rect 36542 4226 36594 4238
rect 36542 4162 36594 4174
rect 37438 4226 37490 4238
rect 37438 4162 37490 4174
rect 34414 4114 34466 4126
rect 29426 4065 30207 4111
rect 29426 4062 29438 4065
rect 31490 4062 31502 4114
rect 31554 4111 31566 4114
rect 31826 4111 31838 4114
rect 31554 4065 31838 4111
rect 31554 4062 31566 4065
rect 31826 4062 31838 4065
rect 31890 4062 31902 4114
rect 34414 4050 34466 4062
rect 1344 3946 38640 3980
rect 1344 3894 4024 3946
rect 4076 3894 4148 3946
rect 4200 3894 4272 3946
rect 4324 3894 4396 3946
rect 4448 3894 4520 3946
rect 4572 3894 4644 3946
rect 4696 3894 4768 3946
rect 4820 3894 4892 3946
rect 4944 3894 5016 3946
rect 5068 3894 5140 3946
rect 5192 3894 24024 3946
rect 24076 3894 24148 3946
rect 24200 3894 24272 3946
rect 24324 3894 24396 3946
rect 24448 3894 24520 3946
rect 24572 3894 24644 3946
rect 24696 3894 24768 3946
rect 24820 3894 24892 3946
rect 24944 3894 25016 3946
rect 25068 3894 25140 3946
rect 25192 3894 38640 3946
rect 1344 3860 38640 3894
rect 9438 3778 9490 3790
rect 11442 3726 11454 3778
rect 11506 3726 11518 3778
rect 9438 3714 9490 3726
rect 3054 3666 3106 3678
rect 2146 3614 2158 3666
rect 2210 3614 2222 3666
rect 3054 3602 3106 3614
rect 9326 3666 9378 3678
rect 27694 3666 27746 3678
rect 13458 3614 13470 3666
rect 13522 3614 13534 3666
rect 32050 3614 32062 3666
rect 32114 3614 32126 3666
rect 9326 3602 9378 3614
rect 27694 3602 27746 3614
rect 1710 3554 1762 3566
rect 1710 3490 1762 3502
rect 3278 3554 3330 3566
rect 3278 3490 3330 3502
rect 3950 3554 4002 3566
rect 5742 3554 5794 3566
rect 8430 3554 8482 3566
rect 4722 3502 4734 3554
rect 4786 3502 4798 3554
rect 6514 3502 6526 3554
rect 6578 3502 6590 3554
rect 7858 3502 7870 3554
rect 7922 3502 7934 3554
rect 3950 3490 4002 3502
rect 5742 3490 5794 3502
rect 8430 3490 8482 3502
rect 9774 3554 9826 3566
rect 11118 3554 11170 3566
rect 17950 3554 18002 3566
rect 10546 3502 10558 3554
rect 10610 3502 10622 3554
rect 11666 3502 11678 3554
rect 11730 3502 11742 3554
rect 12562 3502 12574 3554
rect 12626 3502 12638 3554
rect 14018 3502 14030 3554
rect 14082 3502 14094 3554
rect 15250 3502 15262 3554
rect 15314 3502 15326 3554
rect 16146 3502 16158 3554
rect 16210 3502 16222 3554
rect 17266 3502 17278 3554
rect 17330 3502 17342 3554
rect 9774 3490 9826 3502
rect 11118 3490 11170 3502
rect 17950 3490 18002 3502
rect 18846 3554 18898 3566
rect 18846 3490 18898 3502
rect 19742 3554 19794 3566
rect 19742 3490 19794 3502
rect 21534 3554 21586 3566
rect 21534 3490 21586 3502
rect 22430 3554 22482 3566
rect 26350 3554 26402 3566
rect 32286 3554 32338 3566
rect 23426 3502 23438 3554
rect 23490 3502 23502 3554
rect 27122 3502 27134 3554
rect 27186 3502 27198 3554
rect 28578 3502 28590 3554
rect 28642 3502 28654 3554
rect 34402 3502 34414 3554
rect 34466 3502 34478 3554
rect 36194 3502 36206 3554
rect 36258 3502 36270 3554
rect 36978 3502 36990 3554
rect 37042 3502 37054 3554
rect 37874 3502 37886 3554
rect 37938 3502 37950 3554
rect 22430 3490 22482 3502
rect 26350 3490 26402 3502
rect 32286 3490 32338 3502
rect 4958 3442 5010 3454
rect 6750 3442 6802 3454
rect 8094 3442 8146 3454
rect 3602 3390 3614 3442
rect 3666 3390 3678 3442
rect 4274 3390 4286 3442
rect 4338 3390 4350 3442
rect 6066 3390 6078 3442
rect 6130 3390 6142 3442
rect 7410 3390 7422 3442
rect 7474 3390 7486 3442
rect 4958 3378 5010 3390
rect 6750 3378 6802 3390
rect 8094 3378 8146 3390
rect 8766 3442 8818 3454
rect 8766 3378 8818 3390
rect 10110 3442 10162 3454
rect 10110 3378 10162 3390
rect 10782 3442 10834 3454
rect 16382 3442 16434 3454
rect 12450 3390 12462 3442
rect 12514 3390 12526 3442
rect 14802 3390 14814 3442
rect 14866 3390 14878 3442
rect 10782 3378 10834 3390
rect 16382 3378 16434 3390
rect 17054 3442 17106 3454
rect 17054 3378 17106 3390
rect 18286 3442 18338 3454
rect 18286 3378 18338 3390
rect 19182 3442 19234 3454
rect 19182 3378 19234 3390
rect 20078 3442 20130 3454
rect 20078 3378 20130 3390
rect 20750 3442 20802 3454
rect 20750 3378 20802 3390
rect 21086 3442 21138 3454
rect 21086 3378 21138 3390
rect 21870 3442 21922 3454
rect 21870 3378 21922 3390
rect 22766 3442 22818 3454
rect 22766 3378 22818 3390
rect 23662 3442 23714 3454
rect 23662 3378 23714 3390
rect 24558 3442 24610 3454
rect 24558 3378 24610 3390
rect 24894 3442 24946 3454
rect 24894 3378 24946 3390
rect 25230 3442 25282 3454
rect 25230 3378 25282 3390
rect 25566 3442 25618 3454
rect 25566 3378 25618 3390
rect 26014 3442 26066 3454
rect 26014 3378 26066 3390
rect 26910 3442 26962 3454
rect 26910 3378 26962 3390
rect 28366 3442 28418 3454
rect 28366 3378 28418 3390
rect 29038 3442 29090 3454
rect 29038 3378 29090 3390
rect 29374 3442 29426 3454
rect 29374 3378 29426 3390
rect 29710 3442 29762 3454
rect 29710 3378 29762 3390
rect 30046 3442 30098 3454
rect 30046 3378 30098 3390
rect 30494 3442 30546 3454
rect 30494 3378 30546 3390
rect 30830 3442 30882 3454
rect 30830 3378 30882 3390
rect 31278 3442 31330 3454
rect 33730 3390 33742 3442
rect 33794 3390 33806 3442
rect 34514 3390 34526 3442
rect 34578 3390 34590 3442
rect 31278 3378 31330 3390
rect 7086 3330 7138 3342
rect 7086 3266 7138 3278
rect 31614 3330 31666 3342
rect 31614 3266 31666 3278
rect 35982 3330 36034 3342
rect 35982 3266 36034 3278
rect 36766 3330 36818 3342
rect 36766 3266 36818 3278
rect 37662 3330 37714 3342
rect 37662 3266 37714 3278
rect 1344 3162 38640 3196
rect 1344 3110 14024 3162
rect 14076 3110 14148 3162
rect 14200 3110 14272 3162
rect 14324 3110 14396 3162
rect 14448 3110 14520 3162
rect 14572 3110 14644 3162
rect 14696 3110 14768 3162
rect 14820 3110 14892 3162
rect 14944 3110 15016 3162
rect 15068 3110 15140 3162
rect 15192 3110 34024 3162
rect 34076 3110 34148 3162
rect 34200 3110 34272 3162
rect 34324 3110 34396 3162
rect 34448 3110 34520 3162
rect 34572 3110 34644 3162
rect 34696 3110 34768 3162
rect 34820 3110 34892 3162
rect 34944 3110 35016 3162
rect 35068 3110 35140 3162
rect 35192 3110 38640 3162
rect 1344 3076 38640 3110
rect 7074 2942 7086 2994
rect 7138 2991 7150 2994
rect 9650 2991 9662 2994
rect 7138 2945 9662 2991
rect 7138 2942 7150 2945
rect 9650 2942 9662 2945
rect 9714 2942 9726 2994
<< via1 >>
rect 37214 46510 37266 46562
rect 37886 46510 37938 46562
rect 4024 46230 4076 46282
rect 4148 46230 4200 46282
rect 4272 46230 4324 46282
rect 4396 46230 4448 46282
rect 4520 46230 4572 46282
rect 4644 46230 4696 46282
rect 4768 46230 4820 46282
rect 4892 46230 4944 46282
rect 5016 46230 5068 46282
rect 5140 46230 5192 46282
rect 24024 46230 24076 46282
rect 24148 46230 24200 46282
rect 24272 46230 24324 46282
rect 24396 46230 24448 46282
rect 24520 46230 24572 46282
rect 24644 46230 24696 46282
rect 24768 46230 24820 46282
rect 24892 46230 24944 46282
rect 25016 46230 25068 46282
rect 25140 46230 25192 46282
rect 2718 45950 2770 46002
rect 13582 45950 13634 46002
rect 28814 45950 28866 46002
rect 37886 45950 37938 46002
rect 3502 45838 3554 45890
rect 14142 45838 14194 45890
rect 14814 45838 14866 45890
rect 2046 45726 2098 45778
rect 7870 45726 7922 45778
rect 17726 45726 17778 45778
rect 22654 45726 22706 45778
rect 32510 45726 32562 45778
rect 27918 45614 27970 45666
rect 28366 45614 28418 45666
rect 37214 45614 37266 45666
rect 37438 45614 37490 45666
rect 14024 45446 14076 45498
rect 14148 45446 14200 45498
rect 14272 45446 14324 45498
rect 14396 45446 14448 45498
rect 14520 45446 14572 45498
rect 14644 45446 14696 45498
rect 14768 45446 14820 45498
rect 14892 45446 14944 45498
rect 15016 45446 15068 45498
rect 15140 45446 15192 45498
rect 34024 45446 34076 45498
rect 34148 45446 34200 45498
rect 34272 45446 34324 45498
rect 34396 45446 34448 45498
rect 34520 45446 34572 45498
rect 34644 45446 34696 45498
rect 34768 45446 34820 45498
rect 34892 45446 34944 45498
rect 35016 45446 35068 45498
rect 35140 45446 35192 45498
rect 2158 45278 2210 45330
rect 1710 45166 1762 45218
rect 2718 44942 2770 44994
rect 4024 44662 4076 44714
rect 4148 44662 4200 44714
rect 4272 44662 4324 44714
rect 4396 44662 4448 44714
rect 4520 44662 4572 44714
rect 4644 44662 4696 44714
rect 4768 44662 4820 44714
rect 4892 44662 4944 44714
rect 5016 44662 5068 44714
rect 5140 44662 5192 44714
rect 24024 44662 24076 44714
rect 24148 44662 24200 44714
rect 24272 44662 24324 44714
rect 24396 44662 24448 44714
rect 24520 44662 24572 44714
rect 24644 44662 24696 44714
rect 24768 44662 24820 44714
rect 24892 44662 24944 44714
rect 25016 44662 25068 44714
rect 25140 44662 25192 44714
rect 14024 43878 14076 43930
rect 14148 43878 14200 43930
rect 14272 43878 14324 43930
rect 14396 43878 14448 43930
rect 14520 43878 14572 43930
rect 14644 43878 14696 43930
rect 14768 43878 14820 43930
rect 14892 43878 14944 43930
rect 15016 43878 15068 43930
rect 15140 43878 15192 43930
rect 34024 43878 34076 43930
rect 34148 43878 34200 43930
rect 34272 43878 34324 43930
rect 34396 43878 34448 43930
rect 34520 43878 34572 43930
rect 34644 43878 34696 43930
rect 34768 43878 34820 43930
rect 34892 43878 34944 43930
rect 35016 43878 35068 43930
rect 35140 43878 35192 43930
rect 1710 43598 1762 43650
rect 38222 43262 38274 43314
rect 4024 43094 4076 43146
rect 4148 43094 4200 43146
rect 4272 43094 4324 43146
rect 4396 43094 4448 43146
rect 4520 43094 4572 43146
rect 4644 43094 4696 43146
rect 4768 43094 4820 43146
rect 4892 43094 4944 43146
rect 5016 43094 5068 43146
rect 5140 43094 5192 43146
rect 24024 43094 24076 43146
rect 24148 43094 24200 43146
rect 24272 43094 24324 43146
rect 24396 43094 24448 43146
rect 24520 43094 24572 43146
rect 24644 43094 24696 43146
rect 24768 43094 24820 43146
rect 24892 43094 24944 43146
rect 25016 43094 25068 43146
rect 25140 43094 25192 43146
rect 14024 42310 14076 42362
rect 14148 42310 14200 42362
rect 14272 42310 14324 42362
rect 14396 42310 14448 42362
rect 14520 42310 14572 42362
rect 14644 42310 14696 42362
rect 14768 42310 14820 42362
rect 14892 42310 14944 42362
rect 15016 42310 15068 42362
rect 15140 42310 15192 42362
rect 34024 42310 34076 42362
rect 34148 42310 34200 42362
rect 34272 42310 34324 42362
rect 34396 42310 34448 42362
rect 34520 42310 34572 42362
rect 34644 42310 34696 42362
rect 34768 42310 34820 42362
rect 34892 42310 34944 42362
rect 35016 42310 35068 42362
rect 35140 42310 35192 42362
rect 1710 42030 1762 42082
rect 4024 41526 4076 41578
rect 4148 41526 4200 41578
rect 4272 41526 4324 41578
rect 4396 41526 4448 41578
rect 4520 41526 4572 41578
rect 4644 41526 4696 41578
rect 4768 41526 4820 41578
rect 4892 41526 4944 41578
rect 5016 41526 5068 41578
rect 5140 41526 5192 41578
rect 24024 41526 24076 41578
rect 24148 41526 24200 41578
rect 24272 41526 24324 41578
rect 24396 41526 24448 41578
rect 24520 41526 24572 41578
rect 24644 41526 24696 41578
rect 24768 41526 24820 41578
rect 24892 41526 24944 41578
rect 25016 41526 25068 41578
rect 25140 41526 25192 41578
rect 1710 40910 1762 40962
rect 14024 40742 14076 40794
rect 14148 40742 14200 40794
rect 14272 40742 14324 40794
rect 14396 40742 14448 40794
rect 14520 40742 14572 40794
rect 14644 40742 14696 40794
rect 14768 40742 14820 40794
rect 14892 40742 14944 40794
rect 15016 40742 15068 40794
rect 15140 40742 15192 40794
rect 34024 40742 34076 40794
rect 34148 40742 34200 40794
rect 34272 40742 34324 40794
rect 34396 40742 34448 40794
rect 34520 40742 34572 40794
rect 34644 40742 34696 40794
rect 34768 40742 34820 40794
rect 34892 40742 34944 40794
rect 35016 40742 35068 40794
rect 35140 40742 35192 40794
rect 4024 39958 4076 40010
rect 4148 39958 4200 40010
rect 4272 39958 4324 40010
rect 4396 39958 4448 40010
rect 4520 39958 4572 40010
rect 4644 39958 4696 40010
rect 4768 39958 4820 40010
rect 4892 39958 4944 40010
rect 5016 39958 5068 40010
rect 5140 39958 5192 40010
rect 24024 39958 24076 40010
rect 24148 39958 24200 40010
rect 24272 39958 24324 40010
rect 24396 39958 24448 40010
rect 24520 39958 24572 40010
rect 24644 39958 24696 40010
rect 24768 39958 24820 40010
rect 24892 39958 24944 40010
rect 25016 39958 25068 40010
rect 25140 39958 25192 40010
rect 1710 39342 1762 39394
rect 14024 39174 14076 39226
rect 14148 39174 14200 39226
rect 14272 39174 14324 39226
rect 14396 39174 14448 39226
rect 14520 39174 14572 39226
rect 14644 39174 14696 39226
rect 14768 39174 14820 39226
rect 14892 39174 14944 39226
rect 15016 39174 15068 39226
rect 15140 39174 15192 39226
rect 34024 39174 34076 39226
rect 34148 39174 34200 39226
rect 34272 39174 34324 39226
rect 34396 39174 34448 39226
rect 34520 39174 34572 39226
rect 34644 39174 34696 39226
rect 34768 39174 34820 39226
rect 34892 39174 34944 39226
rect 35016 39174 35068 39226
rect 35140 39174 35192 39226
rect 4024 38390 4076 38442
rect 4148 38390 4200 38442
rect 4272 38390 4324 38442
rect 4396 38390 4448 38442
rect 4520 38390 4572 38442
rect 4644 38390 4696 38442
rect 4768 38390 4820 38442
rect 4892 38390 4944 38442
rect 5016 38390 5068 38442
rect 5140 38390 5192 38442
rect 24024 38390 24076 38442
rect 24148 38390 24200 38442
rect 24272 38390 24324 38442
rect 24396 38390 24448 38442
rect 24520 38390 24572 38442
rect 24644 38390 24696 38442
rect 24768 38390 24820 38442
rect 24892 38390 24944 38442
rect 25016 38390 25068 38442
rect 25140 38390 25192 38442
rect 1710 37774 1762 37826
rect 14024 37606 14076 37658
rect 14148 37606 14200 37658
rect 14272 37606 14324 37658
rect 14396 37606 14448 37658
rect 14520 37606 14572 37658
rect 14644 37606 14696 37658
rect 14768 37606 14820 37658
rect 14892 37606 14944 37658
rect 15016 37606 15068 37658
rect 15140 37606 15192 37658
rect 34024 37606 34076 37658
rect 34148 37606 34200 37658
rect 34272 37606 34324 37658
rect 34396 37606 34448 37658
rect 34520 37606 34572 37658
rect 34644 37606 34696 37658
rect 34768 37606 34820 37658
rect 34892 37606 34944 37658
rect 35016 37606 35068 37658
rect 35140 37606 35192 37658
rect 4024 36822 4076 36874
rect 4148 36822 4200 36874
rect 4272 36822 4324 36874
rect 4396 36822 4448 36874
rect 4520 36822 4572 36874
rect 4644 36822 4696 36874
rect 4768 36822 4820 36874
rect 4892 36822 4944 36874
rect 5016 36822 5068 36874
rect 5140 36822 5192 36874
rect 24024 36822 24076 36874
rect 24148 36822 24200 36874
rect 24272 36822 24324 36874
rect 24396 36822 24448 36874
rect 24520 36822 24572 36874
rect 24644 36822 24696 36874
rect 24768 36822 24820 36874
rect 24892 36822 24944 36874
rect 25016 36822 25068 36874
rect 25140 36822 25192 36874
rect 1710 36318 1762 36370
rect 14024 36038 14076 36090
rect 14148 36038 14200 36090
rect 14272 36038 14324 36090
rect 14396 36038 14448 36090
rect 14520 36038 14572 36090
rect 14644 36038 14696 36090
rect 14768 36038 14820 36090
rect 14892 36038 14944 36090
rect 15016 36038 15068 36090
rect 15140 36038 15192 36090
rect 34024 36038 34076 36090
rect 34148 36038 34200 36090
rect 34272 36038 34324 36090
rect 34396 36038 34448 36090
rect 34520 36038 34572 36090
rect 34644 36038 34696 36090
rect 34768 36038 34820 36090
rect 34892 36038 34944 36090
rect 35016 36038 35068 36090
rect 35140 36038 35192 36090
rect 1710 35758 1762 35810
rect 4024 35254 4076 35306
rect 4148 35254 4200 35306
rect 4272 35254 4324 35306
rect 4396 35254 4448 35306
rect 4520 35254 4572 35306
rect 4644 35254 4696 35306
rect 4768 35254 4820 35306
rect 4892 35254 4944 35306
rect 5016 35254 5068 35306
rect 5140 35254 5192 35306
rect 24024 35254 24076 35306
rect 24148 35254 24200 35306
rect 24272 35254 24324 35306
rect 24396 35254 24448 35306
rect 24520 35254 24572 35306
rect 24644 35254 24696 35306
rect 24768 35254 24820 35306
rect 24892 35254 24944 35306
rect 25016 35254 25068 35306
rect 25140 35254 25192 35306
rect 14024 34470 14076 34522
rect 14148 34470 14200 34522
rect 14272 34470 14324 34522
rect 14396 34470 14448 34522
rect 14520 34470 14572 34522
rect 14644 34470 14696 34522
rect 14768 34470 14820 34522
rect 14892 34470 14944 34522
rect 15016 34470 15068 34522
rect 15140 34470 15192 34522
rect 34024 34470 34076 34522
rect 34148 34470 34200 34522
rect 34272 34470 34324 34522
rect 34396 34470 34448 34522
rect 34520 34470 34572 34522
rect 34644 34470 34696 34522
rect 34768 34470 34820 34522
rect 34892 34470 34944 34522
rect 35016 34470 35068 34522
rect 35140 34470 35192 34522
rect 1710 34190 1762 34242
rect 4024 33686 4076 33738
rect 4148 33686 4200 33738
rect 4272 33686 4324 33738
rect 4396 33686 4448 33738
rect 4520 33686 4572 33738
rect 4644 33686 4696 33738
rect 4768 33686 4820 33738
rect 4892 33686 4944 33738
rect 5016 33686 5068 33738
rect 5140 33686 5192 33738
rect 24024 33686 24076 33738
rect 24148 33686 24200 33738
rect 24272 33686 24324 33738
rect 24396 33686 24448 33738
rect 24520 33686 24572 33738
rect 24644 33686 24696 33738
rect 24768 33686 24820 33738
rect 24892 33686 24944 33738
rect 25016 33686 25068 33738
rect 25140 33686 25192 33738
rect 14024 32902 14076 32954
rect 14148 32902 14200 32954
rect 14272 32902 14324 32954
rect 14396 32902 14448 32954
rect 14520 32902 14572 32954
rect 14644 32902 14696 32954
rect 14768 32902 14820 32954
rect 14892 32902 14944 32954
rect 15016 32902 15068 32954
rect 15140 32902 15192 32954
rect 34024 32902 34076 32954
rect 34148 32902 34200 32954
rect 34272 32902 34324 32954
rect 34396 32902 34448 32954
rect 34520 32902 34572 32954
rect 34644 32902 34696 32954
rect 34768 32902 34820 32954
rect 34892 32902 34944 32954
rect 35016 32902 35068 32954
rect 35140 32902 35192 32954
rect 1710 32622 1762 32674
rect 4024 32118 4076 32170
rect 4148 32118 4200 32170
rect 4272 32118 4324 32170
rect 4396 32118 4448 32170
rect 4520 32118 4572 32170
rect 4644 32118 4696 32170
rect 4768 32118 4820 32170
rect 4892 32118 4944 32170
rect 5016 32118 5068 32170
rect 5140 32118 5192 32170
rect 24024 32118 24076 32170
rect 24148 32118 24200 32170
rect 24272 32118 24324 32170
rect 24396 32118 24448 32170
rect 24520 32118 24572 32170
rect 24644 32118 24696 32170
rect 24768 32118 24820 32170
rect 24892 32118 24944 32170
rect 25016 32118 25068 32170
rect 25140 32118 25192 32170
rect 1710 31502 1762 31554
rect 37662 31502 37714 31554
rect 37886 31502 37938 31554
rect 38222 31502 38274 31554
rect 14024 31334 14076 31386
rect 14148 31334 14200 31386
rect 14272 31334 14324 31386
rect 14396 31334 14448 31386
rect 14520 31334 14572 31386
rect 14644 31334 14696 31386
rect 14768 31334 14820 31386
rect 14892 31334 14944 31386
rect 15016 31334 15068 31386
rect 15140 31334 15192 31386
rect 34024 31334 34076 31386
rect 34148 31334 34200 31386
rect 34272 31334 34324 31386
rect 34396 31334 34448 31386
rect 34520 31334 34572 31386
rect 34644 31334 34696 31386
rect 34768 31334 34820 31386
rect 34892 31334 34944 31386
rect 35016 31334 35068 31386
rect 35140 31334 35192 31386
rect 4024 30550 4076 30602
rect 4148 30550 4200 30602
rect 4272 30550 4324 30602
rect 4396 30550 4448 30602
rect 4520 30550 4572 30602
rect 4644 30550 4696 30602
rect 4768 30550 4820 30602
rect 4892 30550 4944 30602
rect 5016 30550 5068 30602
rect 5140 30550 5192 30602
rect 24024 30550 24076 30602
rect 24148 30550 24200 30602
rect 24272 30550 24324 30602
rect 24396 30550 24448 30602
rect 24520 30550 24572 30602
rect 24644 30550 24696 30602
rect 24768 30550 24820 30602
rect 24892 30550 24944 30602
rect 25016 30550 25068 30602
rect 25140 30550 25192 30602
rect 1710 29934 1762 29986
rect 14024 29766 14076 29818
rect 14148 29766 14200 29818
rect 14272 29766 14324 29818
rect 14396 29766 14448 29818
rect 14520 29766 14572 29818
rect 14644 29766 14696 29818
rect 14768 29766 14820 29818
rect 14892 29766 14944 29818
rect 15016 29766 15068 29818
rect 15140 29766 15192 29818
rect 34024 29766 34076 29818
rect 34148 29766 34200 29818
rect 34272 29766 34324 29818
rect 34396 29766 34448 29818
rect 34520 29766 34572 29818
rect 34644 29766 34696 29818
rect 34768 29766 34820 29818
rect 34892 29766 34944 29818
rect 35016 29766 35068 29818
rect 35140 29766 35192 29818
rect 4024 28982 4076 29034
rect 4148 28982 4200 29034
rect 4272 28982 4324 29034
rect 4396 28982 4448 29034
rect 4520 28982 4572 29034
rect 4644 28982 4696 29034
rect 4768 28982 4820 29034
rect 4892 28982 4944 29034
rect 5016 28982 5068 29034
rect 5140 28982 5192 29034
rect 24024 28982 24076 29034
rect 24148 28982 24200 29034
rect 24272 28982 24324 29034
rect 24396 28982 24448 29034
rect 24520 28982 24572 29034
rect 24644 28982 24696 29034
rect 24768 28982 24820 29034
rect 24892 28982 24944 29034
rect 25016 28982 25068 29034
rect 25140 28982 25192 29034
rect 1710 28366 1762 28418
rect 14024 28198 14076 28250
rect 14148 28198 14200 28250
rect 14272 28198 14324 28250
rect 14396 28198 14448 28250
rect 14520 28198 14572 28250
rect 14644 28198 14696 28250
rect 14768 28198 14820 28250
rect 14892 28198 14944 28250
rect 15016 28198 15068 28250
rect 15140 28198 15192 28250
rect 34024 28198 34076 28250
rect 34148 28198 34200 28250
rect 34272 28198 34324 28250
rect 34396 28198 34448 28250
rect 34520 28198 34572 28250
rect 34644 28198 34696 28250
rect 34768 28198 34820 28250
rect 34892 28198 34944 28250
rect 35016 28198 35068 28250
rect 35140 28198 35192 28250
rect 4024 27414 4076 27466
rect 4148 27414 4200 27466
rect 4272 27414 4324 27466
rect 4396 27414 4448 27466
rect 4520 27414 4572 27466
rect 4644 27414 4696 27466
rect 4768 27414 4820 27466
rect 4892 27414 4944 27466
rect 5016 27414 5068 27466
rect 5140 27414 5192 27466
rect 24024 27414 24076 27466
rect 24148 27414 24200 27466
rect 24272 27414 24324 27466
rect 24396 27414 24448 27466
rect 24520 27414 24572 27466
rect 24644 27414 24696 27466
rect 24768 27414 24820 27466
rect 24892 27414 24944 27466
rect 25016 27414 25068 27466
rect 25140 27414 25192 27466
rect 1710 26798 1762 26850
rect 14024 26630 14076 26682
rect 14148 26630 14200 26682
rect 14272 26630 14324 26682
rect 14396 26630 14448 26682
rect 14520 26630 14572 26682
rect 14644 26630 14696 26682
rect 14768 26630 14820 26682
rect 14892 26630 14944 26682
rect 15016 26630 15068 26682
rect 15140 26630 15192 26682
rect 34024 26630 34076 26682
rect 34148 26630 34200 26682
rect 34272 26630 34324 26682
rect 34396 26630 34448 26682
rect 34520 26630 34572 26682
rect 34644 26630 34696 26682
rect 34768 26630 34820 26682
rect 34892 26630 34944 26682
rect 35016 26630 35068 26682
rect 35140 26630 35192 26682
rect 1710 26350 1762 26402
rect 4024 25846 4076 25898
rect 4148 25846 4200 25898
rect 4272 25846 4324 25898
rect 4396 25846 4448 25898
rect 4520 25846 4572 25898
rect 4644 25846 4696 25898
rect 4768 25846 4820 25898
rect 4892 25846 4944 25898
rect 5016 25846 5068 25898
rect 5140 25846 5192 25898
rect 24024 25846 24076 25898
rect 24148 25846 24200 25898
rect 24272 25846 24324 25898
rect 24396 25846 24448 25898
rect 24520 25846 24572 25898
rect 24644 25846 24696 25898
rect 24768 25846 24820 25898
rect 24892 25846 24944 25898
rect 25016 25846 25068 25898
rect 25140 25846 25192 25898
rect 14024 25062 14076 25114
rect 14148 25062 14200 25114
rect 14272 25062 14324 25114
rect 14396 25062 14448 25114
rect 14520 25062 14572 25114
rect 14644 25062 14696 25114
rect 14768 25062 14820 25114
rect 14892 25062 14944 25114
rect 15016 25062 15068 25114
rect 15140 25062 15192 25114
rect 34024 25062 34076 25114
rect 34148 25062 34200 25114
rect 34272 25062 34324 25114
rect 34396 25062 34448 25114
rect 34520 25062 34572 25114
rect 34644 25062 34696 25114
rect 34768 25062 34820 25114
rect 34892 25062 34944 25114
rect 35016 25062 35068 25114
rect 35140 25062 35192 25114
rect 1710 24782 1762 24834
rect 4024 24278 4076 24330
rect 4148 24278 4200 24330
rect 4272 24278 4324 24330
rect 4396 24278 4448 24330
rect 4520 24278 4572 24330
rect 4644 24278 4696 24330
rect 4768 24278 4820 24330
rect 4892 24278 4944 24330
rect 5016 24278 5068 24330
rect 5140 24278 5192 24330
rect 24024 24278 24076 24330
rect 24148 24278 24200 24330
rect 24272 24278 24324 24330
rect 24396 24278 24448 24330
rect 24520 24278 24572 24330
rect 24644 24278 24696 24330
rect 24768 24278 24820 24330
rect 24892 24278 24944 24330
rect 25016 24278 25068 24330
rect 25140 24278 25192 24330
rect 14024 23494 14076 23546
rect 14148 23494 14200 23546
rect 14272 23494 14324 23546
rect 14396 23494 14448 23546
rect 14520 23494 14572 23546
rect 14644 23494 14696 23546
rect 14768 23494 14820 23546
rect 14892 23494 14944 23546
rect 15016 23494 15068 23546
rect 15140 23494 15192 23546
rect 34024 23494 34076 23546
rect 34148 23494 34200 23546
rect 34272 23494 34324 23546
rect 34396 23494 34448 23546
rect 34520 23494 34572 23546
rect 34644 23494 34696 23546
rect 34768 23494 34820 23546
rect 34892 23494 34944 23546
rect 35016 23494 35068 23546
rect 35140 23494 35192 23546
rect 1710 23214 1762 23266
rect 4024 22710 4076 22762
rect 4148 22710 4200 22762
rect 4272 22710 4324 22762
rect 4396 22710 4448 22762
rect 4520 22710 4572 22762
rect 4644 22710 4696 22762
rect 4768 22710 4820 22762
rect 4892 22710 4944 22762
rect 5016 22710 5068 22762
rect 5140 22710 5192 22762
rect 24024 22710 24076 22762
rect 24148 22710 24200 22762
rect 24272 22710 24324 22762
rect 24396 22710 24448 22762
rect 24520 22710 24572 22762
rect 24644 22710 24696 22762
rect 24768 22710 24820 22762
rect 24892 22710 24944 22762
rect 25016 22710 25068 22762
rect 25140 22710 25192 22762
rect 1710 22094 1762 22146
rect 14024 21926 14076 21978
rect 14148 21926 14200 21978
rect 14272 21926 14324 21978
rect 14396 21926 14448 21978
rect 14520 21926 14572 21978
rect 14644 21926 14696 21978
rect 14768 21926 14820 21978
rect 14892 21926 14944 21978
rect 15016 21926 15068 21978
rect 15140 21926 15192 21978
rect 34024 21926 34076 21978
rect 34148 21926 34200 21978
rect 34272 21926 34324 21978
rect 34396 21926 34448 21978
rect 34520 21926 34572 21978
rect 34644 21926 34696 21978
rect 34768 21926 34820 21978
rect 34892 21926 34944 21978
rect 35016 21926 35068 21978
rect 35140 21926 35192 21978
rect 4024 21142 4076 21194
rect 4148 21142 4200 21194
rect 4272 21142 4324 21194
rect 4396 21142 4448 21194
rect 4520 21142 4572 21194
rect 4644 21142 4696 21194
rect 4768 21142 4820 21194
rect 4892 21142 4944 21194
rect 5016 21142 5068 21194
rect 5140 21142 5192 21194
rect 24024 21142 24076 21194
rect 24148 21142 24200 21194
rect 24272 21142 24324 21194
rect 24396 21142 24448 21194
rect 24520 21142 24572 21194
rect 24644 21142 24696 21194
rect 24768 21142 24820 21194
rect 24892 21142 24944 21194
rect 25016 21142 25068 21194
rect 25140 21142 25192 21194
rect 1710 20526 1762 20578
rect 14024 20358 14076 20410
rect 14148 20358 14200 20410
rect 14272 20358 14324 20410
rect 14396 20358 14448 20410
rect 14520 20358 14572 20410
rect 14644 20358 14696 20410
rect 14768 20358 14820 20410
rect 14892 20358 14944 20410
rect 15016 20358 15068 20410
rect 15140 20358 15192 20410
rect 34024 20358 34076 20410
rect 34148 20358 34200 20410
rect 34272 20358 34324 20410
rect 34396 20358 34448 20410
rect 34520 20358 34572 20410
rect 34644 20358 34696 20410
rect 34768 20358 34820 20410
rect 34892 20358 34944 20410
rect 35016 20358 35068 20410
rect 35140 20358 35192 20410
rect 4024 19574 4076 19626
rect 4148 19574 4200 19626
rect 4272 19574 4324 19626
rect 4396 19574 4448 19626
rect 4520 19574 4572 19626
rect 4644 19574 4696 19626
rect 4768 19574 4820 19626
rect 4892 19574 4944 19626
rect 5016 19574 5068 19626
rect 5140 19574 5192 19626
rect 24024 19574 24076 19626
rect 24148 19574 24200 19626
rect 24272 19574 24324 19626
rect 24396 19574 24448 19626
rect 24520 19574 24572 19626
rect 24644 19574 24696 19626
rect 24768 19574 24820 19626
rect 24892 19574 24944 19626
rect 25016 19574 25068 19626
rect 25140 19574 25192 19626
rect 1710 18958 1762 19010
rect 38222 18958 38274 19010
rect 14024 18790 14076 18842
rect 14148 18790 14200 18842
rect 14272 18790 14324 18842
rect 14396 18790 14448 18842
rect 14520 18790 14572 18842
rect 14644 18790 14696 18842
rect 14768 18790 14820 18842
rect 14892 18790 14944 18842
rect 15016 18790 15068 18842
rect 15140 18790 15192 18842
rect 34024 18790 34076 18842
rect 34148 18790 34200 18842
rect 34272 18790 34324 18842
rect 34396 18790 34448 18842
rect 34520 18790 34572 18842
rect 34644 18790 34696 18842
rect 34768 18790 34820 18842
rect 34892 18790 34944 18842
rect 35016 18790 35068 18842
rect 35140 18790 35192 18842
rect 4024 18006 4076 18058
rect 4148 18006 4200 18058
rect 4272 18006 4324 18058
rect 4396 18006 4448 18058
rect 4520 18006 4572 18058
rect 4644 18006 4696 18058
rect 4768 18006 4820 18058
rect 4892 18006 4944 18058
rect 5016 18006 5068 18058
rect 5140 18006 5192 18058
rect 24024 18006 24076 18058
rect 24148 18006 24200 18058
rect 24272 18006 24324 18058
rect 24396 18006 24448 18058
rect 24520 18006 24572 18058
rect 24644 18006 24696 18058
rect 24768 18006 24820 18058
rect 24892 18006 24944 18058
rect 25016 18006 25068 18058
rect 25140 18006 25192 18058
rect 1710 17502 1762 17554
rect 14024 17222 14076 17274
rect 14148 17222 14200 17274
rect 14272 17222 14324 17274
rect 14396 17222 14448 17274
rect 14520 17222 14572 17274
rect 14644 17222 14696 17274
rect 14768 17222 14820 17274
rect 14892 17222 14944 17274
rect 15016 17222 15068 17274
rect 15140 17222 15192 17274
rect 34024 17222 34076 17274
rect 34148 17222 34200 17274
rect 34272 17222 34324 17274
rect 34396 17222 34448 17274
rect 34520 17222 34572 17274
rect 34644 17222 34696 17274
rect 34768 17222 34820 17274
rect 34892 17222 34944 17274
rect 35016 17222 35068 17274
rect 35140 17222 35192 17274
rect 1710 16942 1762 16994
rect 4024 16438 4076 16490
rect 4148 16438 4200 16490
rect 4272 16438 4324 16490
rect 4396 16438 4448 16490
rect 4520 16438 4572 16490
rect 4644 16438 4696 16490
rect 4768 16438 4820 16490
rect 4892 16438 4944 16490
rect 5016 16438 5068 16490
rect 5140 16438 5192 16490
rect 24024 16438 24076 16490
rect 24148 16438 24200 16490
rect 24272 16438 24324 16490
rect 24396 16438 24448 16490
rect 24520 16438 24572 16490
rect 24644 16438 24696 16490
rect 24768 16438 24820 16490
rect 24892 16438 24944 16490
rect 25016 16438 25068 16490
rect 25140 16438 25192 16490
rect 14024 15654 14076 15706
rect 14148 15654 14200 15706
rect 14272 15654 14324 15706
rect 14396 15654 14448 15706
rect 14520 15654 14572 15706
rect 14644 15654 14696 15706
rect 14768 15654 14820 15706
rect 14892 15654 14944 15706
rect 15016 15654 15068 15706
rect 15140 15654 15192 15706
rect 34024 15654 34076 15706
rect 34148 15654 34200 15706
rect 34272 15654 34324 15706
rect 34396 15654 34448 15706
rect 34520 15654 34572 15706
rect 34644 15654 34696 15706
rect 34768 15654 34820 15706
rect 34892 15654 34944 15706
rect 35016 15654 35068 15706
rect 35140 15654 35192 15706
rect 1710 15374 1762 15426
rect 4024 14870 4076 14922
rect 4148 14870 4200 14922
rect 4272 14870 4324 14922
rect 4396 14870 4448 14922
rect 4520 14870 4572 14922
rect 4644 14870 4696 14922
rect 4768 14870 4820 14922
rect 4892 14870 4944 14922
rect 5016 14870 5068 14922
rect 5140 14870 5192 14922
rect 24024 14870 24076 14922
rect 24148 14870 24200 14922
rect 24272 14870 24324 14922
rect 24396 14870 24448 14922
rect 24520 14870 24572 14922
rect 24644 14870 24696 14922
rect 24768 14870 24820 14922
rect 24892 14870 24944 14922
rect 25016 14870 25068 14922
rect 25140 14870 25192 14922
rect 14024 14086 14076 14138
rect 14148 14086 14200 14138
rect 14272 14086 14324 14138
rect 14396 14086 14448 14138
rect 14520 14086 14572 14138
rect 14644 14086 14696 14138
rect 14768 14086 14820 14138
rect 14892 14086 14944 14138
rect 15016 14086 15068 14138
rect 15140 14086 15192 14138
rect 34024 14086 34076 14138
rect 34148 14086 34200 14138
rect 34272 14086 34324 14138
rect 34396 14086 34448 14138
rect 34520 14086 34572 14138
rect 34644 14086 34696 14138
rect 34768 14086 34820 14138
rect 34892 14086 34944 14138
rect 35016 14086 35068 14138
rect 35140 14086 35192 14138
rect 1710 13806 1762 13858
rect 4024 13302 4076 13354
rect 4148 13302 4200 13354
rect 4272 13302 4324 13354
rect 4396 13302 4448 13354
rect 4520 13302 4572 13354
rect 4644 13302 4696 13354
rect 4768 13302 4820 13354
rect 4892 13302 4944 13354
rect 5016 13302 5068 13354
rect 5140 13302 5192 13354
rect 24024 13302 24076 13354
rect 24148 13302 24200 13354
rect 24272 13302 24324 13354
rect 24396 13302 24448 13354
rect 24520 13302 24572 13354
rect 24644 13302 24696 13354
rect 24768 13302 24820 13354
rect 24892 13302 24944 13354
rect 25016 13302 25068 13354
rect 25140 13302 25192 13354
rect 1710 12686 1762 12738
rect 14024 12518 14076 12570
rect 14148 12518 14200 12570
rect 14272 12518 14324 12570
rect 14396 12518 14448 12570
rect 14520 12518 14572 12570
rect 14644 12518 14696 12570
rect 14768 12518 14820 12570
rect 14892 12518 14944 12570
rect 15016 12518 15068 12570
rect 15140 12518 15192 12570
rect 34024 12518 34076 12570
rect 34148 12518 34200 12570
rect 34272 12518 34324 12570
rect 34396 12518 34448 12570
rect 34520 12518 34572 12570
rect 34644 12518 34696 12570
rect 34768 12518 34820 12570
rect 34892 12518 34944 12570
rect 35016 12518 35068 12570
rect 35140 12518 35192 12570
rect 4024 11734 4076 11786
rect 4148 11734 4200 11786
rect 4272 11734 4324 11786
rect 4396 11734 4448 11786
rect 4520 11734 4572 11786
rect 4644 11734 4696 11786
rect 4768 11734 4820 11786
rect 4892 11734 4944 11786
rect 5016 11734 5068 11786
rect 5140 11734 5192 11786
rect 24024 11734 24076 11786
rect 24148 11734 24200 11786
rect 24272 11734 24324 11786
rect 24396 11734 24448 11786
rect 24520 11734 24572 11786
rect 24644 11734 24696 11786
rect 24768 11734 24820 11786
rect 24892 11734 24944 11786
rect 25016 11734 25068 11786
rect 25140 11734 25192 11786
rect 1710 11118 1762 11170
rect 14024 10950 14076 11002
rect 14148 10950 14200 11002
rect 14272 10950 14324 11002
rect 14396 10950 14448 11002
rect 14520 10950 14572 11002
rect 14644 10950 14696 11002
rect 14768 10950 14820 11002
rect 14892 10950 14944 11002
rect 15016 10950 15068 11002
rect 15140 10950 15192 11002
rect 34024 10950 34076 11002
rect 34148 10950 34200 11002
rect 34272 10950 34324 11002
rect 34396 10950 34448 11002
rect 34520 10950 34572 11002
rect 34644 10950 34696 11002
rect 34768 10950 34820 11002
rect 34892 10950 34944 11002
rect 35016 10950 35068 11002
rect 35140 10950 35192 11002
rect 11902 10558 11954 10610
rect 12126 10558 12178 10610
rect 12574 10558 12626 10610
rect 12910 10558 12962 10610
rect 12014 10446 12066 10498
rect 13358 10446 13410 10498
rect 12686 10334 12738 10386
rect 13358 10334 13410 10386
rect 4024 10166 4076 10218
rect 4148 10166 4200 10218
rect 4272 10166 4324 10218
rect 4396 10166 4448 10218
rect 4520 10166 4572 10218
rect 4644 10166 4696 10218
rect 4768 10166 4820 10218
rect 4892 10166 4944 10218
rect 5016 10166 5068 10218
rect 5140 10166 5192 10218
rect 24024 10166 24076 10218
rect 24148 10166 24200 10218
rect 24272 10166 24324 10218
rect 24396 10166 24448 10218
rect 24520 10166 24572 10218
rect 24644 10166 24696 10218
rect 24768 10166 24820 10218
rect 24892 10166 24944 10218
rect 25016 10166 25068 10218
rect 25140 10166 25192 10218
rect 12686 9886 12738 9938
rect 9774 9774 9826 9826
rect 7758 9662 7810 9714
rect 8318 9662 8370 9714
rect 10558 9662 10610 9714
rect 1710 9550 1762 9602
rect 7646 9550 7698 9602
rect 13694 9550 13746 9602
rect 14024 9382 14076 9434
rect 14148 9382 14200 9434
rect 14272 9382 14324 9434
rect 14396 9382 14448 9434
rect 14520 9382 14572 9434
rect 14644 9382 14696 9434
rect 14768 9382 14820 9434
rect 14892 9382 14944 9434
rect 15016 9382 15068 9434
rect 15140 9382 15192 9434
rect 34024 9382 34076 9434
rect 34148 9382 34200 9434
rect 34272 9382 34324 9434
rect 34396 9382 34448 9434
rect 34520 9382 34572 9434
rect 34644 9382 34696 9434
rect 34768 9382 34820 9434
rect 34892 9382 34944 9434
rect 35016 9382 35068 9434
rect 35140 9382 35192 9434
rect 10446 9214 10498 9266
rect 10782 9102 10834 9154
rect 10222 8990 10274 9042
rect 10446 8990 10498 9042
rect 11342 8990 11394 9042
rect 6414 8878 6466 8930
rect 7422 8878 7474 8930
rect 7870 8878 7922 8930
rect 8430 8878 8482 8930
rect 8766 8878 8818 8930
rect 9662 8878 9714 8930
rect 13470 8878 13522 8930
rect 4024 8598 4076 8650
rect 4148 8598 4200 8650
rect 4272 8598 4324 8650
rect 4396 8598 4448 8650
rect 4520 8598 4572 8650
rect 4644 8598 4696 8650
rect 4768 8598 4820 8650
rect 4892 8598 4944 8650
rect 5016 8598 5068 8650
rect 5140 8598 5192 8650
rect 24024 8598 24076 8650
rect 24148 8598 24200 8650
rect 24272 8598 24324 8650
rect 24396 8598 24448 8650
rect 24520 8598 24572 8650
rect 24644 8598 24696 8650
rect 24768 8598 24820 8650
rect 24892 8598 24944 8650
rect 25016 8598 25068 8650
rect 25140 8598 25192 8650
rect 7422 8318 7474 8370
rect 7758 8318 7810 8370
rect 5966 8206 6018 8258
rect 10782 8206 10834 8258
rect 12798 8206 12850 8258
rect 13470 8206 13522 8258
rect 1710 8094 1762 8146
rect 5630 8094 5682 8146
rect 8206 8094 8258 8146
rect 8318 8094 8370 8146
rect 9662 8094 9714 8146
rect 12910 8094 12962 8146
rect 14254 8094 14306 8146
rect 3054 7982 3106 8034
rect 3390 7982 3442 8034
rect 3950 7982 4002 8034
rect 4622 7982 4674 8034
rect 5182 7982 5234 8034
rect 5742 7982 5794 8034
rect 6526 7982 6578 8034
rect 6974 7982 7026 8034
rect 7646 7982 7698 8034
rect 7982 7982 8034 8034
rect 8766 7982 8818 8034
rect 9214 7982 9266 8034
rect 16494 7982 16546 8034
rect 14024 7814 14076 7866
rect 14148 7814 14200 7866
rect 14272 7814 14324 7866
rect 14396 7814 14448 7866
rect 14520 7814 14572 7866
rect 14644 7814 14696 7866
rect 14768 7814 14820 7866
rect 14892 7814 14944 7866
rect 15016 7814 15068 7866
rect 15140 7814 15192 7866
rect 34024 7814 34076 7866
rect 34148 7814 34200 7866
rect 34272 7814 34324 7866
rect 34396 7814 34448 7866
rect 34520 7814 34572 7866
rect 34644 7814 34696 7866
rect 34768 7814 34820 7866
rect 34892 7814 34944 7866
rect 35016 7814 35068 7866
rect 35140 7814 35192 7866
rect 8878 7646 8930 7698
rect 8990 7534 9042 7586
rect 10110 7534 10162 7586
rect 13134 7534 13186 7586
rect 2942 7422 2994 7474
rect 7198 7422 7250 7474
rect 7534 7422 7586 7474
rect 7758 7422 7810 7474
rect 8206 7422 8258 7474
rect 8654 7422 8706 7474
rect 11678 7422 11730 7474
rect 13694 7422 13746 7474
rect 14702 7422 14754 7474
rect 1934 7310 1986 7362
rect 3502 7310 3554 7362
rect 3950 7310 4002 7362
rect 4286 7310 4338 7362
rect 6414 7310 6466 7362
rect 7982 7310 8034 7362
rect 9774 7310 9826 7362
rect 11790 7310 11842 7362
rect 14254 7310 14306 7362
rect 15150 7310 15202 7362
rect 15598 7310 15650 7362
rect 3502 7198 3554 7250
rect 3950 7198 4002 7250
rect 14030 7198 14082 7250
rect 14254 7198 14306 7250
rect 15598 7198 15650 7250
rect 4024 7030 4076 7082
rect 4148 7030 4200 7082
rect 4272 7030 4324 7082
rect 4396 7030 4448 7082
rect 4520 7030 4572 7082
rect 4644 7030 4696 7082
rect 4768 7030 4820 7082
rect 4892 7030 4944 7082
rect 5016 7030 5068 7082
rect 5140 7030 5192 7082
rect 24024 7030 24076 7082
rect 24148 7030 24200 7082
rect 24272 7030 24324 7082
rect 24396 7030 24448 7082
rect 24520 7030 24572 7082
rect 24644 7030 24696 7082
rect 24768 7030 24820 7082
rect 24892 7030 24944 7082
rect 25016 7030 25068 7082
rect 25140 7030 25192 7082
rect 1822 6750 1874 6802
rect 7198 6750 7250 6802
rect 17614 6750 17666 6802
rect 4734 6638 4786 6690
rect 6526 6638 6578 6690
rect 6750 6638 6802 6690
rect 10222 6638 10274 6690
rect 10670 6638 10722 6690
rect 13470 6638 13522 6690
rect 15486 6638 15538 6690
rect 20526 6638 20578 6690
rect 21422 6638 21474 6690
rect 3950 6526 4002 6578
rect 5742 6526 5794 6578
rect 5854 6526 5906 6578
rect 5518 6414 5570 6466
rect 6190 6470 6242 6522
rect 7310 6526 7362 6578
rect 8654 6526 8706 6578
rect 11230 6526 11282 6578
rect 13582 6526 13634 6578
rect 16046 6526 16098 6578
rect 19742 6526 19794 6578
rect 37886 6526 37938 6578
rect 38222 6526 38274 6578
rect 6302 6414 6354 6466
rect 7086 6414 7138 6466
rect 7758 6414 7810 6466
rect 7870 6414 7922 6466
rect 7982 6414 8034 6466
rect 8206 6414 8258 6466
rect 11118 6414 11170 6466
rect 13022 6414 13074 6466
rect 15486 6414 15538 6466
rect 37662 6414 37714 6466
rect 14024 6246 14076 6298
rect 14148 6246 14200 6298
rect 14272 6246 14324 6298
rect 14396 6246 14448 6298
rect 14520 6246 14572 6298
rect 14644 6246 14696 6298
rect 14768 6246 14820 6298
rect 14892 6246 14944 6298
rect 15016 6246 15068 6298
rect 15140 6246 15192 6298
rect 34024 6246 34076 6298
rect 34148 6246 34200 6298
rect 34272 6246 34324 6298
rect 34396 6246 34448 6298
rect 34520 6246 34572 6298
rect 34644 6246 34696 6298
rect 34768 6246 34820 6298
rect 34892 6246 34944 6298
rect 35016 6246 35068 6298
rect 35140 6246 35192 6298
rect 6862 6078 6914 6130
rect 20750 6078 20802 6130
rect 2270 5966 2322 6018
rect 5966 5966 6018 6018
rect 6526 5966 6578 6018
rect 7422 5966 7474 6018
rect 7646 5966 7698 6018
rect 8094 5966 8146 6018
rect 8990 5966 9042 6018
rect 11342 5966 11394 6018
rect 1934 5854 1986 5906
rect 5518 5854 5570 5906
rect 6302 5854 6354 5906
rect 6974 5854 7026 5906
rect 8542 5854 8594 5906
rect 8654 5854 8706 5906
rect 14814 5854 14866 5906
rect 15374 5854 15426 5906
rect 2046 5742 2098 5794
rect 2606 5742 2658 5794
rect 4734 5742 4786 5794
rect 6078 5742 6130 5794
rect 7982 5742 8034 5794
rect 8878 5742 8930 5794
rect 15822 5742 15874 5794
rect 16158 5742 16210 5794
rect 16830 5742 16882 5794
rect 17502 5742 17554 5794
rect 17950 5742 18002 5794
rect 24334 5742 24386 5794
rect 7086 5630 7138 5682
rect 4024 5462 4076 5514
rect 4148 5462 4200 5514
rect 4272 5462 4324 5514
rect 4396 5462 4448 5514
rect 4520 5462 4572 5514
rect 4644 5462 4696 5514
rect 4768 5462 4820 5514
rect 4892 5462 4944 5514
rect 5016 5462 5068 5514
rect 5140 5462 5192 5514
rect 24024 5462 24076 5514
rect 24148 5462 24200 5514
rect 24272 5462 24324 5514
rect 24396 5462 24448 5514
rect 24520 5462 24572 5514
rect 24644 5462 24696 5514
rect 24768 5462 24820 5514
rect 24892 5462 24944 5514
rect 25016 5462 25068 5514
rect 25140 5462 25192 5514
rect 2158 5294 2210 5346
rect 6078 5182 6130 5234
rect 11566 5182 11618 5234
rect 2830 5070 2882 5122
rect 3390 5070 3442 5122
rect 4062 5070 4114 5122
rect 11118 5070 11170 5122
rect 12126 5070 12178 5122
rect 12238 5070 12290 5122
rect 13806 5070 13858 5122
rect 14366 5070 14418 5122
rect 16606 5070 16658 5122
rect 22206 5070 22258 5122
rect 26014 5070 26066 5122
rect 28142 5070 28194 5122
rect 30158 5070 30210 5122
rect 32286 5070 32338 5122
rect 34974 5070 35026 5122
rect 3726 4958 3778 5010
rect 4398 4958 4450 5010
rect 5070 4958 5122 5010
rect 11678 4958 11730 5010
rect 12574 4958 12626 5010
rect 14030 4958 14082 5010
rect 15598 4958 15650 5010
rect 17054 4958 17106 5010
rect 22878 4958 22930 5010
rect 24894 4958 24946 5010
rect 30270 4958 30322 5010
rect 32846 4958 32898 5010
rect 1710 4846 1762 4898
rect 4846 4846 4898 4898
rect 4958 4846 5010 4898
rect 11454 4846 11506 4898
rect 12462 4846 12514 4898
rect 15150 4846 15202 4898
rect 18734 4846 18786 4898
rect 19518 4846 19570 4898
rect 20526 4846 20578 4898
rect 21534 4846 21586 4898
rect 21982 4846 22034 4898
rect 23774 4846 23826 4898
rect 26462 4846 26514 4898
rect 26910 4846 26962 4898
rect 33854 4846 33906 4898
rect 34414 4846 34466 4898
rect 14024 4678 14076 4730
rect 14148 4678 14200 4730
rect 14272 4678 14324 4730
rect 14396 4678 14448 4730
rect 14520 4678 14572 4730
rect 14644 4678 14696 4730
rect 14768 4678 14820 4730
rect 14892 4678 14944 4730
rect 15016 4678 15068 4730
rect 15140 4678 15192 4730
rect 34024 4678 34076 4730
rect 34148 4678 34200 4730
rect 34272 4678 34324 4730
rect 34396 4678 34448 4730
rect 34520 4678 34572 4730
rect 34644 4678 34696 4730
rect 34768 4678 34820 4730
rect 34892 4678 34944 4730
rect 35016 4678 35068 4730
rect 35140 4678 35192 4730
rect 6862 4510 6914 4562
rect 8206 4510 8258 4562
rect 8990 4510 9042 4562
rect 9886 4510 9938 4562
rect 11118 4510 11170 4562
rect 11678 4510 11730 4562
rect 16382 4510 16434 4562
rect 25342 4510 25394 4562
rect 3838 4398 3890 4450
rect 5406 4398 5458 4450
rect 6078 4398 6130 4450
rect 7422 4398 7474 4450
rect 7646 4398 7698 4450
rect 8094 4398 8146 4450
rect 12126 4398 12178 4450
rect 14702 4398 14754 4450
rect 17390 4398 17442 4450
rect 19406 4398 19458 4450
rect 20862 4398 20914 4450
rect 23774 4398 23826 4450
rect 25902 4398 25954 4450
rect 27918 4398 27970 4450
rect 33070 4398 33122 4450
rect 33742 4398 33794 4450
rect 34750 4398 34802 4450
rect 35086 4398 35138 4450
rect 4622 4286 4674 4338
rect 5294 4286 5346 4338
rect 6414 4286 6466 4338
rect 6862 4286 6914 4338
rect 7982 4286 8034 4338
rect 8766 4286 8818 4338
rect 9886 4286 9938 4338
rect 10110 4286 10162 4338
rect 11566 4286 11618 4338
rect 13582 4286 13634 4338
rect 16046 4286 16098 4338
rect 18286 4286 18338 4338
rect 20414 4286 20466 4338
rect 24110 4286 24162 4338
rect 25342 4286 25394 4338
rect 27470 4286 27522 4338
rect 33294 4286 33346 4338
rect 33966 4286 34018 4338
rect 34414 4286 34466 4338
rect 35310 4286 35362 4338
rect 1710 4174 1762 4226
rect 9998 4174 10050 4226
rect 11230 4174 11282 4226
rect 16942 4174 16994 4226
rect 17726 4174 17778 4226
rect 18622 4174 18674 4226
rect 24558 4174 24610 4226
rect 29486 4174 29538 4226
rect 29934 4174 29986 4226
rect 30158 4174 30210 4226
rect 30494 4174 30546 4226
rect 7086 4062 7138 4114
rect 22766 4062 22818 4114
rect 29374 4062 29426 4114
rect 31838 4174 31890 4226
rect 32510 4174 32562 4226
rect 35982 4174 36034 4226
rect 36542 4174 36594 4226
rect 37438 4174 37490 4226
rect 31502 4062 31554 4114
rect 31838 4062 31890 4114
rect 34414 4062 34466 4114
rect 4024 3894 4076 3946
rect 4148 3894 4200 3946
rect 4272 3894 4324 3946
rect 4396 3894 4448 3946
rect 4520 3894 4572 3946
rect 4644 3894 4696 3946
rect 4768 3894 4820 3946
rect 4892 3894 4944 3946
rect 5016 3894 5068 3946
rect 5140 3894 5192 3946
rect 24024 3894 24076 3946
rect 24148 3894 24200 3946
rect 24272 3894 24324 3946
rect 24396 3894 24448 3946
rect 24520 3894 24572 3946
rect 24644 3894 24696 3946
rect 24768 3894 24820 3946
rect 24892 3894 24944 3946
rect 25016 3894 25068 3946
rect 25140 3894 25192 3946
rect 9438 3726 9490 3778
rect 11454 3726 11506 3778
rect 2158 3614 2210 3666
rect 3054 3614 3106 3666
rect 9326 3614 9378 3666
rect 13470 3614 13522 3666
rect 27694 3614 27746 3666
rect 32062 3614 32114 3666
rect 1710 3502 1762 3554
rect 3278 3502 3330 3554
rect 3950 3502 4002 3554
rect 4734 3502 4786 3554
rect 5742 3502 5794 3554
rect 6526 3502 6578 3554
rect 7870 3502 7922 3554
rect 8430 3502 8482 3554
rect 9774 3502 9826 3554
rect 10558 3502 10610 3554
rect 11118 3502 11170 3554
rect 11678 3502 11730 3554
rect 12574 3502 12626 3554
rect 14030 3502 14082 3554
rect 15262 3502 15314 3554
rect 16158 3502 16210 3554
rect 17278 3502 17330 3554
rect 17950 3502 18002 3554
rect 18846 3502 18898 3554
rect 19742 3502 19794 3554
rect 21534 3502 21586 3554
rect 22430 3502 22482 3554
rect 23438 3502 23490 3554
rect 26350 3502 26402 3554
rect 27134 3502 27186 3554
rect 28590 3502 28642 3554
rect 32286 3502 32338 3554
rect 34414 3502 34466 3554
rect 36206 3502 36258 3554
rect 36990 3502 37042 3554
rect 37886 3502 37938 3554
rect 3614 3390 3666 3442
rect 4286 3390 4338 3442
rect 4958 3390 5010 3442
rect 6078 3390 6130 3442
rect 6750 3390 6802 3442
rect 7422 3390 7474 3442
rect 8094 3390 8146 3442
rect 8766 3390 8818 3442
rect 10110 3390 10162 3442
rect 10782 3390 10834 3442
rect 12462 3390 12514 3442
rect 14814 3390 14866 3442
rect 16382 3390 16434 3442
rect 17054 3390 17106 3442
rect 18286 3390 18338 3442
rect 19182 3390 19234 3442
rect 20078 3390 20130 3442
rect 20750 3390 20802 3442
rect 21086 3390 21138 3442
rect 21870 3390 21922 3442
rect 22766 3390 22818 3442
rect 23662 3390 23714 3442
rect 24558 3390 24610 3442
rect 24894 3390 24946 3442
rect 25230 3390 25282 3442
rect 25566 3390 25618 3442
rect 26014 3390 26066 3442
rect 26910 3390 26962 3442
rect 28366 3390 28418 3442
rect 29038 3390 29090 3442
rect 29374 3390 29426 3442
rect 29710 3390 29762 3442
rect 30046 3390 30098 3442
rect 30494 3390 30546 3442
rect 30830 3390 30882 3442
rect 31278 3390 31330 3442
rect 33742 3390 33794 3442
rect 34526 3390 34578 3442
rect 7086 3278 7138 3330
rect 31614 3278 31666 3330
rect 35982 3278 36034 3330
rect 36766 3278 36818 3330
rect 37662 3278 37714 3330
rect 14024 3110 14076 3162
rect 14148 3110 14200 3162
rect 14272 3110 14324 3162
rect 14396 3110 14448 3162
rect 14520 3110 14572 3162
rect 14644 3110 14696 3162
rect 14768 3110 14820 3162
rect 14892 3110 14944 3162
rect 15016 3110 15068 3162
rect 15140 3110 15192 3162
rect 34024 3110 34076 3162
rect 34148 3110 34200 3162
rect 34272 3110 34324 3162
rect 34396 3110 34448 3162
rect 34520 3110 34572 3162
rect 34644 3110 34696 3162
rect 34768 3110 34820 3162
rect 34892 3110 34944 3162
rect 35016 3110 35068 3162
rect 35140 3110 35192 3162
rect 7086 2942 7138 2994
rect 9662 2942 9714 2994
<< metal2 >>
rect 2688 49200 2800 50000
rect 7616 49200 7728 50000
rect 12544 49200 12656 50000
rect 17472 49200 17584 50000
rect 22400 49200 22512 50000
rect 27328 49200 27440 50000
rect 32256 49200 32368 50000
rect 37184 49200 37296 50000
rect 2044 47012 2100 47022
rect 2044 45778 2100 46956
rect 2716 46002 2772 49200
rect 4008 46284 5208 46294
rect 4064 46282 4112 46284
rect 4168 46282 4216 46284
rect 4076 46230 4112 46282
rect 4200 46230 4216 46282
rect 4064 46228 4112 46230
rect 4168 46228 4216 46230
rect 4272 46282 4320 46284
rect 4376 46282 4424 46284
rect 4480 46282 4528 46284
rect 4376 46230 4396 46282
rect 4480 46230 4520 46282
rect 4272 46228 4320 46230
rect 4376 46228 4424 46230
rect 4480 46228 4528 46230
rect 4584 46228 4632 46284
rect 4688 46282 4736 46284
rect 4792 46282 4840 46284
rect 4896 46282 4944 46284
rect 4696 46230 4736 46282
rect 4820 46230 4840 46282
rect 4688 46228 4736 46230
rect 4792 46228 4840 46230
rect 4896 46228 4944 46230
rect 5000 46282 5048 46284
rect 5104 46282 5152 46284
rect 5000 46230 5016 46282
rect 5104 46230 5140 46282
rect 5000 46228 5048 46230
rect 5104 46228 5152 46230
rect 4008 46218 5208 46228
rect 2716 45950 2718 46002
rect 2770 45950 2772 46002
rect 2716 45938 2772 45950
rect 3500 45890 3556 45902
rect 3500 45838 3502 45890
rect 3554 45838 3556 45890
rect 2044 45726 2046 45778
rect 2098 45726 2100 45778
rect 2044 45714 2100 45726
rect 2156 45780 2212 45790
rect 2156 45330 2212 45724
rect 2156 45278 2158 45330
rect 2210 45278 2212 45330
rect 2156 45266 2212 45278
rect 1708 45218 1764 45230
rect 1708 45166 1710 45218
rect 1762 45166 1764 45218
rect 1708 44436 1764 45166
rect 1708 44370 1764 44380
rect 1820 44996 1876 45006
rect 1708 43650 1764 43662
rect 1708 43598 1710 43650
rect 1762 43598 1764 43650
rect 1708 43092 1764 43598
rect 1708 43026 1764 43036
rect 1708 42082 1764 42094
rect 1708 42030 1710 42082
rect 1762 42030 1764 42082
rect 1708 41748 1764 42030
rect 1708 41682 1764 41692
rect 1708 40962 1764 40974
rect 1708 40910 1710 40962
rect 1762 40910 1764 40962
rect 1708 40404 1764 40910
rect 1708 40338 1764 40348
rect 1708 39394 1764 39406
rect 1708 39342 1710 39394
rect 1762 39342 1764 39394
rect 1708 39060 1764 39342
rect 1708 38994 1764 39004
rect 1708 37828 1764 37838
rect 1708 37734 1764 37772
rect 1708 36372 1764 36382
rect 1708 36278 1764 36316
rect 1708 35810 1764 35822
rect 1708 35758 1710 35810
rect 1762 35758 1764 35810
rect 1708 35028 1764 35758
rect 1708 34962 1764 34972
rect 1708 34242 1764 34254
rect 1708 34190 1710 34242
rect 1762 34190 1764 34242
rect 1708 33684 1764 34190
rect 1708 33618 1764 33628
rect 1708 32674 1764 32686
rect 1708 32622 1710 32674
rect 1762 32622 1764 32674
rect 1708 32340 1764 32622
rect 1708 32274 1764 32284
rect 1708 31554 1764 31566
rect 1708 31502 1710 31554
rect 1762 31502 1764 31554
rect 1708 30996 1764 31502
rect 1708 30930 1764 30940
rect 1708 29986 1764 29998
rect 1708 29934 1710 29986
rect 1762 29934 1764 29986
rect 1708 29652 1764 29934
rect 1708 29586 1764 29596
rect 1708 28420 1764 28430
rect 1708 28326 1764 28364
rect 1708 26964 1764 26974
rect 1708 26850 1764 26908
rect 1708 26798 1710 26850
rect 1762 26798 1764 26850
rect 1708 26786 1764 26798
rect 1708 26402 1764 26414
rect 1708 26350 1710 26402
rect 1762 26350 1764 26402
rect 1708 25620 1764 26350
rect 1708 25554 1764 25564
rect 1708 24834 1764 24846
rect 1708 24782 1710 24834
rect 1762 24782 1764 24834
rect 1708 24276 1764 24782
rect 1708 24210 1764 24220
rect 1708 23266 1764 23278
rect 1708 23214 1710 23266
rect 1762 23214 1764 23266
rect 1708 22932 1764 23214
rect 1708 22866 1764 22876
rect 1708 22146 1764 22158
rect 1708 22094 1710 22146
rect 1762 22094 1764 22146
rect 1708 21588 1764 22094
rect 1708 21522 1764 21532
rect 1708 20578 1764 20590
rect 1708 20526 1710 20578
rect 1762 20526 1764 20578
rect 1708 20244 1764 20526
rect 1708 20178 1764 20188
rect 1708 19012 1764 19022
rect 1708 18918 1764 18956
rect 1708 17556 1764 17566
rect 1708 17462 1764 17500
rect 1708 16994 1764 17006
rect 1708 16942 1710 16994
rect 1762 16942 1764 16994
rect 1708 16212 1764 16942
rect 1708 16146 1764 16156
rect 1708 15426 1764 15438
rect 1708 15374 1710 15426
rect 1762 15374 1764 15426
rect 1708 14868 1764 15374
rect 1708 14802 1764 14812
rect 1708 13858 1764 13870
rect 1708 13806 1710 13858
rect 1762 13806 1764 13858
rect 1708 13524 1764 13806
rect 1708 13458 1764 13468
rect 1708 12738 1764 12750
rect 1708 12686 1710 12738
rect 1762 12686 1764 12738
rect 1708 12180 1764 12686
rect 1708 12114 1764 12124
rect 1708 11170 1764 11182
rect 1708 11118 1710 11170
rect 1762 11118 1764 11170
rect 1708 10836 1764 11118
rect 1708 10770 1764 10780
rect 1708 9604 1764 9614
rect 1708 9510 1764 9548
rect 1708 8148 1764 8158
rect 1708 8054 1764 8092
rect 1820 6802 1876 44940
rect 2716 44996 2772 45006
rect 2716 44902 2772 44940
rect 3500 44996 3556 45838
rect 7644 45780 7700 49200
rect 12572 46004 12628 49200
rect 12572 45938 12628 45948
rect 13580 46004 13636 46014
rect 13580 45910 13636 45948
rect 14140 45892 14196 45902
rect 14812 45892 14868 45902
rect 13804 45890 14868 45892
rect 13804 45838 14142 45890
rect 14194 45838 14814 45890
rect 14866 45838 14868 45890
rect 13804 45836 14868 45838
rect 7868 45780 7924 45790
rect 7644 45778 7924 45780
rect 7644 45726 7870 45778
rect 7922 45726 7924 45778
rect 7644 45724 7924 45726
rect 7868 45714 7924 45724
rect 3500 44930 3556 44940
rect 4008 44716 5208 44726
rect 4064 44714 4112 44716
rect 4168 44714 4216 44716
rect 4076 44662 4112 44714
rect 4200 44662 4216 44714
rect 4064 44660 4112 44662
rect 4168 44660 4216 44662
rect 4272 44714 4320 44716
rect 4376 44714 4424 44716
rect 4480 44714 4528 44716
rect 4376 44662 4396 44714
rect 4480 44662 4520 44714
rect 4272 44660 4320 44662
rect 4376 44660 4424 44662
rect 4480 44660 4528 44662
rect 4584 44660 4632 44716
rect 4688 44714 4736 44716
rect 4792 44714 4840 44716
rect 4896 44714 4944 44716
rect 4696 44662 4736 44714
rect 4820 44662 4840 44714
rect 4688 44660 4736 44662
rect 4792 44660 4840 44662
rect 4896 44660 4944 44662
rect 5000 44714 5048 44716
rect 5104 44714 5152 44716
rect 5000 44662 5016 44714
rect 5104 44662 5140 44714
rect 5000 44660 5048 44662
rect 5104 44660 5152 44662
rect 4008 44650 5208 44660
rect 4008 43148 5208 43158
rect 4064 43146 4112 43148
rect 4168 43146 4216 43148
rect 4076 43094 4112 43146
rect 4200 43094 4216 43146
rect 4064 43092 4112 43094
rect 4168 43092 4216 43094
rect 4272 43146 4320 43148
rect 4376 43146 4424 43148
rect 4480 43146 4528 43148
rect 4376 43094 4396 43146
rect 4480 43094 4520 43146
rect 4272 43092 4320 43094
rect 4376 43092 4424 43094
rect 4480 43092 4528 43094
rect 4584 43092 4632 43148
rect 4688 43146 4736 43148
rect 4792 43146 4840 43148
rect 4896 43146 4944 43148
rect 4696 43094 4736 43146
rect 4820 43094 4840 43146
rect 4688 43092 4736 43094
rect 4792 43092 4840 43094
rect 4896 43092 4944 43094
rect 5000 43146 5048 43148
rect 5104 43146 5152 43148
rect 5000 43094 5016 43146
rect 5104 43094 5140 43146
rect 5000 43092 5048 43094
rect 5104 43092 5152 43094
rect 4008 43082 5208 43092
rect 4008 41580 5208 41590
rect 4064 41578 4112 41580
rect 4168 41578 4216 41580
rect 4076 41526 4112 41578
rect 4200 41526 4216 41578
rect 4064 41524 4112 41526
rect 4168 41524 4216 41526
rect 4272 41578 4320 41580
rect 4376 41578 4424 41580
rect 4480 41578 4528 41580
rect 4376 41526 4396 41578
rect 4480 41526 4520 41578
rect 4272 41524 4320 41526
rect 4376 41524 4424 41526
rect 4480 41524 4528 41526
rect 4584 41524 4632 41580
rect 4688 41578 4736 41580
rect 4792 41578 4840 41580
rect 4896 41578 4944 41580
rect 4696 41526 4736 41578
rect 4820 41526 4840 41578
rect 4688 41524 4736 41526
rect 4792 41524 4840 41526
rect 4896 41524 4944 41526
rect 5000 41578 5048 41580
rect 5104 41578 5152 41580
rect 5000 41526 5016 41578
rect 5104 41526 5140 41578
rect 5000 41524 5048 41526
rect 5104 41524 5152 41526
rect 4008 41514 5208 41524
rect 4008 40012 5208 40022
rect 4064 40010 4112 40012
rect 4168 40010 4216 40012
rect 4076 39958 4112 40010
rect 4200 39958 4216 40010
rect 4064 39956 4112 39958
rect 4168 39956 4216 39958
rect 4272 40010 4320 40012
rect 4376 40010 4424 40012
rect 4480 40010 4528 40012
rect 4376 39958 4396 40010
rect 4480 39958 4520 40010
rect 4272 39956 4320 39958
rect 4376 39956 4424 39958
rect 4480 39956 4528 39958
rect 4584 39956 4632 40012
rect 4688 40010 4736 40012
rect 4792 40010 4840 40012
rect 4896 40010 4944 40012
rect 4696 39958 4736 40010
rect 4820 39958 4840 40010
rect 4688 39956 4736 39958
rect 4792 39956 4840 39958
rect 4896 39956 4944 39958
rect 5000 40010 5048 40012
rect 5104 40010 5152 40012
rect 5000 39958 5016 40010
rect 5104 39958 5140 40010
rect 5000 39956 5048 39958
rect 5104 39956 5152 39958
rect 4008 39946 5208 39956
rect 4008 38444 5208 38454
rect 4064 38442 4112 38444
rect 4168 38442 4216 38444
rect 4076 38390 4112 38442
rect 4200 38390 4216 38442
rect 4064 38388 4112 38390
rect 4168 38388 4216 38390
rect 4272 38442 4320 38444
rect 4376 38442 4424 38444
rect 4480 38442 4528 38444
rect 4376 38390 4396 38442
rect 4480 38390 4520 38442
rect 4272 38388 4320 38390
rect 4376 38388 4424 38390
rect 4480 38388 4528 38390
rect 4584 38388 4632 38444
rect 4688 38442 4736 38444
rect 4792 38442 4840 38444
rect 4896 38442 4944 38444
rect 4696 38390 4736 38442
rect 4820 38390 4840 38442
rect 4688 38388 4736 38390
rect 4792 38388 4840 38390
rect 4896 38388 4944 38390
rect 5000 38442 5048 38444
rect 5104 38442 5152 38444
rect 5000 38390 5016 38442
rect 5104 38390 5140 38442
rect 5000 38388 5048 38390
rect 5104 38388 5152 38390
rect 4008 38378 5208 38388
rect 4008 36876 5208 36886
rect 4064 36874 4112 36876
rect 4168 36874 4216 36876
rect 4076 36822 4112 36874
rect 4200 36822 4216 36874
rect 4064 36820 4112 36822
rect 4168 36820 4216 36822
rect 4272 36874 4320 36876
rect 4376 36874 4424 36876
rect 4480 36874 4528 36876
rect 4376 36822 4396 36874
rect 4480 36822 4520 36874
rect 4272 36820 4320 36822
rect 4376 36820 4424 36822
rect 4480 36820 4528 36822
rect 4584 36820 4632 36876
rect 4688 36874 4736 36876
rect 4792 36874 4840 36876
rect 4896 36874 4944 36876
rect 4696 36822 4736 36874
rect 4820 36822 4840 36874
rect 4688 36820 4736 36822
rect 4792 36820 4840 36822
rect 4896 36820 4944 36822
rect 5000 36874 5048 36876
rect 5104 36874 5152 36876
rect 5000 36822 5016 36874
rect 5104 36822 5140 36874
rect 5000 36820 5048 36822
rect 5104 36820 5152 36822
rect 4008 36810 5208 36820
rect 4008 35308 5208 35318
rect 4064 35306 4112 35308
rect 4168 35306 4216 35308
rect 4076 35254 4112 35306
rect 4200 35254 4216 35306
rect 4064 35252 4112 35254
rect 4168 35252 4216 35254
rect 4272 35306 4320 35308
rect 4376 35306 4424 35308
rect 4480 35306 4528 35308
rect 4376 35254 4396 35306
rect 4480 35254 4520 35306
rect 4272 35252 4320 35254
rect 4376 35252 4424 35254
rect 4480 35252 4528 35254
rect 4584 35252 4632 35308
rect 4688 35306 4736 35308
rect 4792 35306 4840 35308
rect 4896 35306 4944 35308
rect 4696 35254 4736 35306
rect 4820 35254 4840 35306
rect 4688 35252 4736 35254
rect 4792 35252 4840 35254
rect 4896 35252 4944 35254
rect 5000 35306 5048 35308
rect 5104 35306 5152 35308
rect 5000 35254 5016 35306
rect 5104 35254 5140 35306
rect 5000 35252 5048 35254
rect 5104 35252 5152 35254
rect 4008 35242 5208 35252
rect 4008 33740 5208 33750
rect 4064 33738 4112 33740
rect 4168 33738 4216 33740
rect 4076 33686 4112 33738
rect 4200 33686 4216 33738
rect 4064 33684 4112 33686
rect 4168 33684 4216 33686
rect 4272 33738 4320 33740
rect 4376 33738 4424 33740
rect 4480 33738 4528 33740
rect 4376 33686 4396 33738
rect 4480 33686 4520 33738
rect 4272 33684 4320 33686
rect 4376 33684 4424 33686
rect 4480 33684 4528 33686
rect 4584 33684 4632 33740
rect 4688 33738 4736 33740
rect 4792 33738 4840 33740
rect 4896 33738 4944 33740
rect 4696 33686 4736 33738
rect 4820 33686 4840 33738
rect 4688 33684 4736 33686
rect 4792 33684 4840 33686
rect 4896 33684 4944 33686
rect 5000 33738 5048 33740
rect 5104 33738 5152 33740
rect 5000 33686 5016 33738
rect 5104 33686 5140 33738
rect 5000 33684 5048 33686
rect 5104 33684 5152 33686
rect 4008 33674 5208 33684
rect 4008 32172 5208 32182
rect 4064 32170 4112 32172
rect 4168 32170 4216 32172
rect 4076 32118 4112 32170
rect 4200 32118 4216 32170
rect 4064 32116 4112 32118
rect 4168 32116 4216 32118
rect 4272 32170 4320 32172
rect 4376 32170 4424 32172
rect 4480 32170 4528 32172
rect 4376 32118 4396 32170
rect 4480 32118 4520 32170
rect 4272 32116 4320 32118
rect 4376 32116 4424 32118
rect 4480 32116 4528 32118
rect 4584 32116 4632 32172
rect 4688 32170 4736 32172
rect 4792 32170 4840 32172
rect 4896 32170 4944 32172
rect 4696 32118 4736 32170
rect 4820 32118 4840 32170
rect 4688 32116 4736 32118
rect 4792 32116 4840 32118
rect 4896 32116 4944 32118
rect 5000 32170 5048 32172
rect 5104 32170 5152 32172
rect 5000 32118 5016 32170
rect 5104 32118 5140 32170
rect 5000 32116 5048 32118
rect 5104 32116 5152 32118
rect 4008 32106 5208 32116
rect 4008 30604 5208 30614
rect 4064 30602 4112 30604
rect 4168 30602 4216 30604
rect 4076 30550 4112 30602
rect 4200 30550 4216 30602
rect 4064 30548 4112 30550
rect 4168 30548 4216 30550
rect 4272 30602 4320 30604
rect 4376 30602 4424 30604
rect 4480 30602 4528 30604
rect 4376 30550 4396 30602
rect 4480 30550 4520 30602
rect 4272 30548 4320 30550
rect 4376 30548 4424 30550
rect 4480 30548 4528 30550
rect 4584 30548 4632 30604
rect 4688 30602 4736 30604
rect 4792 30602 4840 30604
rect 4896 30602 4944 30604
rect 4696 30550 4736 30602
rect 4820 30550 4840 30602
rect 4688 30548 4736 30550
rect 4792 30548 4840 30550
rect 4896 30548 4944 30550
rect 5000 30602 5048 30604
rect 5104 30602 5152 30604
rect 5000 30550 5016 30602
rect 5104 30550 5140 30602
rect 5000 30548 5048 30550
rect 5104 30548 5152 30550
rect 4008 30538 5208 30548
rect 4008 29036 5208 29046
rect 4064 29034 4112 29036
rect 4168 29034 4216 29036
rect 4076 28982 4112 29034
rect 4200 28982 4216 29034
rect 4064 28980 4112 28982
rect 4168 28980 4216 28982
rect 4272 29034 4320 29036
rect 4376 29034 4424 29036
rect 4480 29034 4528 29036
rect 4376 28982 4396 29034
rect 4480 28982 4520 29034
rect 4272 28980 4320 28982
rect 4376 28980 4424 28982
rect 4480 28980 4528 28982
rect 4584 28980 4632 29036
rect 4688 29034 4736 29036
rect 4792 29034 4840 29036
rect 4896 29034 4944 29036
rect 4696 28982 4736 29034
rect 4820 28982 4840 29034
rect 4688 28980 4736 28982
rect 4792 28980 4840 28982
rect 4896 28980 4944 28982
rect 5000 29034 5048 29036
rect 5104 29034 5152 29036
rect 5000 28982 5016 29034
rect 5104 28982 5140 29034
rect 5000 28980 5048 28982
rect 5104 28980 5152 28982
rect 4008 28970 5208 28980
rect 4008 27468 5208 27478
rect 4064 27466 4112 27468
rect 4168 27466 4216 27468
rect 4076 27414 4112 27466
rect 4200 27414 4216 27466
rect 4064 27412 4112 27414
rect 4168 27412 4216 27414
rect 4272 27466 4320 27468
rect 4376 27466 4424 27468
rect 4480 27466 4528 27468
rect 4376 27414 4396 27466
rect 4480 27414 4520 27466
rect 4272 27412 4320 27414
rect 4376 27412 4424 27414
rect 4480 27412 4528 27414
rect 4584 27412 4632 27468
rect 4688 27466 4736 27468
rect 4792 27466 4840 27468
rect 4896 27466 4944 27468
rect 4696 27414 4736 27466
rect 4820 27414 4840 27466
rect 4688 27412 4736 27414
rect 4792 27412 4840 27414
rect 4896 27412 4944 27414
rect 5000 27466 5048 27468
rect 5104 27466 5152 27468
rect 5000 27414 5016 27466
rect 5104 27414 5140 27466
rect 5000 27412 5048 27414
rect 5104 27412 5152 27414
rect 4008 27402 5208 27412
rect 4008 25900 5208 25910
rect 4064 25898 4112 25900
rect 4168 25898 4216 25900
rect 4076 25846 4112 25898
rect 4200 25846 4216 25898
rect 4064 25844 4112 25846
rect 4168 25844 4216 25846
rect 4272 25898 4320 25900
rect 4376 25898 4424 25900
rect 4480 25898 4528 25900
rect 4376 25846 4396 25898
rect 4480 25846 4520 25898
rect 4272 25844 4320 25846
rect 4376 25844 4424 25846
rect 4480 25844 4528 25846
rect 4584 25844 4632 25900
rect 4688 25898 4736 25900
rect 4792 25898 4840 25900
rect 4896 25898 4944 25900
rect 4696 25846 4736 25898
rect 4820 25846 4840 25898
rect 4688 25844 4736 25846
rect 4792 25844 4840 25846
rect 4896 25844 4944 25846
rect 5000 25898 5048 25900
rect 5104 25898 5152 25900
rect 5000 25846 5016 25898
rect 5104 25846 5140 25898
rect 5000 25844 5048 25846
rect 5104 25844 5152 25846
rect 4008 25834 5208 25844
rect 4008 24332 5208 24342
rect 4064 24330 4112 24332
rect 4168 24330 4216 24332
rect 4076 24278 4112 24330
rect 4200 24278 4216 24330
rect 4064 24276 4112 24278
rect 4168 24276 4216 24278
rect 4272 24330 4320 24332
rect 4376 24330 4424 24332
rect 4480 24330 4528 24332
rect 4376 24278 4396 24330
rect 4480 24278 4520 24330
rect 4272 24276 4320 24278
rect 4376 24276 4424 24278
rect 4480 24276 4528 24278
rect 4584 24276 4632 24332
rect 4688 24330 4736 24332
rect 4792 24330 4840 24332
rect 4896 24330 4944 24332
rect 4696 24278 4736 24330
rect 4820 24278 4840 24330
rect 4688 24276 4736 24278
rect 4792 24276 4840 24278
rect 4896 24276 4944 24278
rect 5000 24330 5048 24332
rect 5104 24330 5152 24332
rect 5000 24278 5016 24330
rect 5104 24278 5140 24330
rect 5000 24276 5048 24278
rect 5104 24276 5152 24278
rect 4008 24266 5208 24276
rect 4008 22764 5208 22774
rect 4064 22762 4112 22764
rect 4168 22762 4216 22764
rect 4076 22710 4112 22762
rect 4200 22710 4216 22762
rect 4064 22708 4112 22710
rect 4168 22708 4216 22710
rect 4272 22762 4320 22764
rect 4376 22762 4424 22764
rect 4480 22762 4528 22764
rect 4376 22710 4396 22762
rect 4480 22710 4520 22762
rect 4272 22708 4320 22710
rect 4376 22708 4424 22710
rect 4480 22708 4528 22710
rect 4584 22708 4632 22764
rect 4688 22762 4736 22764
rect 4792 22762 4840 22764
rect 4896 22762 4944 22764
rect 4696 22710 4736 22762
rect 4820 22710 4840 22762
rect 4688 22708 4736 22710
rect 4792 22708 4840 22710
rect 4896 22708 4944 22710
rect 5000 22762 5048 22764
rect 5104 22762 5152 22764
rect 5000 22710 5016 22762
rect 5104 22710 5140 22762
rect 5000 22708 5048 22710
rect 5104 22708 5152 22710
rect 4008 22698 5208 22708
rect 4008 21196 5208 21206
rect 4064 21194 4112 21196
rect 4168 21194 4216 21196
rect 4076 21142 4112 21194
rect 4200 21142 4216 21194
rect 4064 21140 4112 21142
rect 4168 21140 4216 21142
rect 4272 21194 4320 21196
rect 4376 21194 4424 21196
rect 4480 21194 4528 21196
rect 4376 21142 4396 21194
rect 4480 21142 4520 21194
rect 4272 21140 4320 21142
rect 4376 21140 4424 21142
rect 4480 21140 4528 21142
rect 4584 21140 4632 21196
rect 4688 21194 4736 21196
rect 4792 21194 4840 21196
rect 4896 21194 4944 21196
rect 4696 21142 4736 21194
rect 4820 21142 4840 21194
rect 4688 21140 4736 21142
rect 4792 21140 4840 21142
rect 4896 21140 4944 21142
rect 5000 21194 5048 21196
rect 5104 21194 5152 21196
rect 5000 21142 5016 21194
rect 5104 21142 5140 21194
rect 5000 21140 5048 21142
rect 5104 21140 5152 21142
rect 4008 21130 5208 21140
rect 4008 19628 5208 19638
rect 4064 19626 4112 19628
rect 4168 19626 4216 19628
rect 4076 19574 4112 19626
rect 4200 19574 4216 19626
rect 4064 19572 4112 19574
rect 4168 19572 4216 19574
rect 4272 19626 4320 19628
rect 4376 19626 4424 19628
rect 4480 19626 4528 19628
rect 4376 19574 4396 19626
rect 4480 19574 4520 19626
rect 4272 19572 4320 19574
rect 4376 19572 4424 19574
rect 4480 19572 4528 19574
rect 4584 19572 4632 19628
rect 4688 19626 4736 19628
rect 4792 19626 4840 19628
rect 4896 19626 4944 19628
rect 4696 19574 4736 19626
rect 4820 19574 4840 19626
rect 4688 19572 4736 19574
rect 4792 19572 4840 19574
rect 4896 19572 4944 19574
rect 5000 19626 5048 19628
rect 5104 19626 5152 19628
rect 5000 19574 5016 19626
rect 5104 19574 5140 19626
rect 5000 19572 5048 19574
rect 5104 19572 5152 19574
rect 4008 19562 5208 19572
rect 4008 18060 5208 18070
rect 4064 18058 4112 18060
rect 4168 18058 4216 18060
rect 4076 18006 4112 18058
rect 4200 18006 4216 18058
rect 4064 18004 4112 18006
rect 4168 18004 4216 18006
rect 4272 18058 4320 18060
rect 4376 18058 4424 18060
rect 4480 18058 4528 18060
rect 4376 18006 4396 18058
rect 4480 18006 4520 18058
rect 4272 18004 4320 18006
rect 4376 18004 4424 18006
rect 4480 18004 4528 18006
rect 4584 18004 4632 18060
rect 4688 18058 4736 18060
rect 4792 18058 4840 18060
rect 4896 18058 4944 18060
rect 4696 18006 4736 18058
rect 4820 18006 4840 18058
rect 4688 18004 4736 18006
rect 4792 18004 4840 18006
rect 4896 18004 4944 18006
rect 5000 18058 5048 18060
rect 5104 18058 5152 18060
rect 5000 18006 5016 18058
rect 5104 18006 5140 18058
rect 5000 18004 5048 18006
rect 5104 18004 5152 18006
rect 4008 17994 5208 18004
rect 4008 16492 5208 16502
rect 4064 16490 4112 16492
rect 4168 16490 4216 16492
rect 4076 16438 4112 16490
rect 4200 16438 4216 16490
rect 4064 16436 4112 16438
rect 4168 16436 4216 16438
rect 4272 16490 4320 16492
rect 4376 16490 4424 16492
rect 4480 16490 4528 16492
rect 4376 16438 4396 16490
rect 4480 16438 4520 16490
rect 4272 16436 4320 16438
rect 4376 16436 4424 16438
rect 4480 16436 4528 16438
rect 4584 16436 4632 16492
rect 4688 16490 4736 16492
rect 4792 16490 4840 16492
rect 4896 16490 4944 16492
rect 4696 16438 4736 16490
rect 4820 16438 4840 16490
rect 4688 16436 4736 16438
rect 4792 16436 4840 16438
rect 4896 16436 4944 16438
rect 5000 16490 5048 16492
rect 5104 16490 5152 16492
rect 5000 16438 5016 16490
rect 5104 16438 5140 16490
rect 5000 16436 5048 16438
rect 5104 16436 5152 16438
rect 4008 16426 5208 16436
rect 4008 14924 5208 14934
rect 4064 14922 4112 14924
rect 4168 14922 4216 14924
rect 4076 14870 4112 14922
rect 4200 14870 4216 14922
rect 4064 14868 4112 14870
rect 4168 14868 4216 14870
rect 4272 14922 4320 14924
rect 4376 14922 4424 14924
rect 4480 14922 4528 14924
rect 4376 14870 4396 14922
rect 4480 14870 4520 14922
rect 4272 14868 4320 14870
rect 4376 14868 4424 14870
rect 4480 14868 4528 14870
rect 4584 14868 4632 14924
rect 4688 14922 4736 14924
rect 4792 14922 4840 14924
rect 4896 14922 4944 14924
rect 4696 14870 4736 14922
rect 4820 14870 4840 14922
rect 4688 14868 4736 14870
rect 4792 14868 4840 14870
rect 4896 14868 4944 14870
rect 5000 14922 5048 14924
rect 5104 14922 5152 14924
rect 5000 14870 5016 14922
rect 5104 14870 5140 14922
rect 5000 14868 5048 14870
rect 5104 14868 5152 14870
rect 4008 14858 5208 14868
rect 4008 13356 5208 13366
rect 4064 13354 4112 13356
rect 4168 13354 4216 13356
rect 4076 13302 4112 13354
rect 4200 13302 4216 13354
rect 4064 13300 4112 13302
rect 4168 13300 4216 13302
rect 4272 13354 4320 13356
rect 4376 13354 4424 13356
rect 4480 13354 4528 13356
rect 4376 13302 4396 13354
rect 4480 13302 4520 13354
rect 4272 13300 4320 13302
rect 4376 13300 4424 13302
rect 4480 13300 4528 13302
rect 4584 13300 4632 13356
rect 4688 13354 4736 13356
rect 4792 13354 4840 13356
rect 4896 13354 4944 13356
rect 4696 13302 4736 13354
rect 4820 13302 4840 13354
rect 4688 13300 4736 13302
rect 4792 13300 4840 13302
rect 4896 13300 4944 13302
rect 5000 13354 5048 13356
rect 5104 13354 5152 13356
rect 5000 13302 5016 13354
rect 5104 13302 5140 13354
rect 5000 13300 5048 13302
rect 5104 13300 5152 13302
rect 4008 13290 5208 13300
rect 4008 11788 5208 11798
rect 4064 11786 4112 11788
rect 4168 11786 4216 11788
rect 4076 11734 4112 11786
rect 4200 11734 4216 11786
rect 4064 11732 4112 11734
rect 4168 11732 4216 11734
rect 4272 11786 4320 11788
rect 4376 11786 4424 11788
rect 4480 11786 4528 11788
rect 4376 11734 4396 11786
rect 4480 11734 4520 11786
rect 4272 11732 4320 11734
rect 4376 11732 4424 11734
rect 4480 11732 4528 11734
rect 4584 11732 4632 11788
rect 4688 11786 4736 11788
rect 4792 11786 4840 11788
rect 4896 11786 4944 11788
rect 4696 11734 4736 11786
rect 4820 11734 4840 11786
rect 4688 11732 4736 11734
rect 4792 11732 4840 11734
rect 4896 11732 4944 11734
rect 5000 11786 5048 11788
rect 5104 11786 5152 11788
rect 5000 11734 5016 11786
rect 5104 11734 5140 11786
rect 5000 11732 5048 11734
rect 5104 11732 5152 11734
rect 4008 11722 5208 11732
rect 10332 10612 10388 10622
rect 4008 10220 5208 10230
rect 4064 10218 4112 10220
rect 4168 10218 4216 10220
rect 4076 10166 4112 10218
rect 4200 10166 4216 10218
rect 4064 10164 4112 10166
rect 4168 10164 4216 10166
rect 4272 10218 4320 10220
rect 4376 10218 4424 10220
rect 4480 10218 4528 10220
rect 4376 10166 4396 10218
rect 4480 10166 4520 10218
rect 4272 10164 4320 10166
rect 4376 10164 4424 10166
rect 4480 10164 4528 10166
rect 4584 10164 4632 10220
rect 4688 10218 4736 10220
rect 4792 10218 4840 10220
rect 4896 10218 4944 10220
rect 4696 10166 4736 10218
rect 4820 10166 4840 10218
rect 4688 10164 4736 10166
rect 4792 10164 4840 10166
rect 4896 10164 4944 10166
rect 5000 10218 5048 10220
rect 5104 10218 5152 10220
rect 5000 10166 5016 10218
rect 5104 10166 5140 10218
rect 5000 10164 5048 10166
rect 5104 10164 5152 10166
rect 4008 10154 5208 10164
rect 9772 9826 9828 9838
rect 9772 9774 9774 9826
rect 9826 9774 9828 9826
rect 7756 9716 7812 9726
rect 7756 9622 7812 9660
rect 8316 9716 8372 9726
rect 8316 9622 8372 9660
rect 7644 9604 7700 9614
rect 7532 9602 7700 9604
rect 7532 9550 7646 9602
rect 7698 9550 7700 9602
rect 7532 9548 7700 9550
rect 6412 8932 6468 8942
rect 6300 8930 6468 8932
rect 6300 8878 6414 8930
rect 6466 8878 6468 8930
rect 6300 8876 6468 8878
rect 4008 8652 5208 8662
rect 4064 8650 4112 8652
rect 4168 8650 4216 8652
rect 4076 8598 4112 8650
rect 4200 8598 4216 8650
rect 4064 8596 4112 8598
rect 4168 8596 4216 8598
rect 4272 8650 4320 8652
rect 4376 8650 4424 8652
rect 4480 8650 4528 8652
rect 4376 8598 4396 8650
rect 4480 8598 4520 8650
rect 4272 8596 4320 8598
rect 4376 8596 4424 8598
rect 4480 8596 4528 8598
rect 4584 8596 4632 8652
rect 4688 8650 4736 8652
rect 4792 8650 4840 8652
rect 4896 8650 4944 8652
rect 4696 8598 4736 8650
rect 4820 8598 4840 8650
rect 4688 8596 4736 8598
rect 4792 8596 4840 8598
rect 4896 8596 4944 8598
rect 5000 8650 5048 8652
rect 5104 8650 5152 8652
rect 5000 8598 5016 8650
rect 5104 8598 5140 8650
rect 5000 8596 5048 8598
rect 5104 8596 5152 8598
rect 4008 8586 5208 8596
rect 5964 8260 6020 8270
rect 5964 8166 6020 8204
rect 5628 8146 5684 8158
rect 5628 8094 5630 8146
rect 5682 8094 5684 8146
rect 3052 8034 3108 8046
rect 3052 7982 3054 8034
rect 3106 7982 3108 8034
rect 2940 7474 2996 7486
rect 2940 7422 2942 7474
rect 2994 7422 2996 7474
rect 1820 6750 1822 6802
rect 1874 6750 1876 6802
rect 1820 6738 1876 6750
rect 1932 7362 1988 7374
rect 1932 7310 1934 7362
rect 1986 7310 1988 7362
rect 1932 6804 1988 7310
rect 2940 7252 2996 7422
rect 2940 7186 2996 7196
rect 1932 6738 1988 6748
rect 2268 6468 2324 6478
rect 2268 6018 2324 6412
rect 2268 5966 2270 6018
rect 2322 5966 2324 6018
rect 2268 5954 2324 5966
rect 2604 6132 2660 6142
rect 1932 5908 1988 5918
rect 1932 5814 1988 5852
rect 2044 5794 2100 5806
rect 2044 5742 2046 5794
rect 2098 5742 2100 5794
rect 1708 4898 1764 4910
rect 1708 4846 1710 4898
rect 1762 4846 1764 4898
rect 1708 4452 1764 4846
rect 1708 4386 1764 4396
rect 2044 4452 2100 5742
rect 2604 5796 2660 6076
rect 2604 5794 2884 5796
rect 2604 5742 2606 5794
rect 2658 5742 2884 5794
rect 2604 5740 2884 5742
rect 2604 5730 2660 5740
rect 2156 5348 2212 5358
rect 2156 5254 2212 5292
rect 2044 4386 2100 4396
rect 2492 5124 2548 5134
rect 1708 4226 1764 4238
rect 1708 4174 1710 4226
rect 1762 4174 1764 4226
rect 1708 3554 1764 4174
rect 1708 3502 1710 3554
rect 1762 3502 1764 3554
rect 1708 3490 1764 3502
rect 2156 3666 2212 3678
rect 2156 3614 2158 3666
rect 2210 3614 2212 3666
rect 2156 2772 2212 3614
rect 2156 2706 2212 2716
rect 2492 800 2548 5068
rect 2828 5122 2884 5740
rect 2828 5070 2830 5122
rect 2882 5070 2884 5122
rect 2828 5058 2884 5070
rect 3052 5124 3108 7982
rect 3052 5058 3108 5068
rect 3388 8034 3444 8046
rect 3948 8036 4004 8046
rect 4620 8036 4676 8046
rect 3388 7982 3390 8034
rect 3442 7982 3444 8034
rect 3388 5122 3444 7982
rect 3612 8034 4004 8036
rect 3612 7982 3950 8034
rect 4002 7982 4004 8034
rect 3612 7980 4004 7982
rect 3500 7362 3556 7374
rect 3500 7310 3502 7362
rect 3554 7310 3556 7362
rect 3500 7250 3556 7310
rect 3500 7198 3502 7250
rect 3554 7198 3556 7250
rect 3500 6356 3556 7198
rect 3500 6290 3556 6300
rect 3388 5070 3390 5122
rect 3442 5070 3444 5122
rect 3052 4116 3108 4126
rect 3052 3666 3108 4060
rect 3388 3780 3444 5070
rect 3612 4340 3668 7980
rect 3948 7970 4004 7980
rect 4060 8034 4676 8036
rect 4060 7982 4622 8034
rect 4674 7982 4676 8034
rect 4060 7980 4676 7982
rect 4060 7588 4116 7980
rect 4620 7970 4676 7980
rect 5180 8036 5236 8046
rect 5180 8034 5348 8036
rect 5180 7982 5182 8034
rect 5234 7982 5348 8034
rect 5180 7980 5348 7982
rect 5180 7970 5236 7980
rect 3836 7532 4116 7588
rect 3724 5348 3780 5358
rect 3724 5010 3780 5292
rect 3724 4958 3726 5010
rect 3778 4958 3780 5010
rect 3724 4946 3780 4958
rect 3836 4676 3892 7532
rect 3948 7362 4004 7374
rect 3948 7310 3950 7362
rect 4002 7310 4004 7362
rect 3948 7250 4004 7310
rect 3948 7198 3950 7250
rect 4002 7198 4004 7250
rect 3948 7186 4004 7198
rect 4284 7362 4340 7374
rect 4284 7310 4286 7362
rect 4338 7310 4340 7362
rect 4284 7252 4340 7310
rect 4284 7186 4340 7196
rect 4008 7084 5208 7094
rect 4064 7082 4112 7084
rect 4168 7082 4216 7084
rect 4076 7030 4112 7082
rect 4200 7030 4216 7082
rect 4064 7028 4112 7030
rect 4168 7028 4216 7030
rect 4272 7082 4320 7084
rect 4376 7082 4424 7084
rect 4480 7082 4528 7084
rect 4376 7030 4396 7082
rect 4480 7030 4520 7082
rect 4272 7028 4320 7030
rect 4376 7028 4424 7030
rect 4480 7028 4528 7030
rect 4584 7028 4632 7084
rect 4688 7082 4736 7084
rect 4792 7082 4840 7084
rect 4896 7082 4944 7084
rect 4696 7030 4736 7082
rect 4820 7030 4840 7082
rect 4688 7028 4736 7030
rect 4792 7028 4840 7030
rect 4896 7028 4944 7030
rect 5000 7082 5048 7084
rect 5104 7082 5152 7084
rect 5000 7030 5016 7082
rect 5104 7030 5140 7082
rect 5000 7028 5048 7030
rect 5104 7028 5152 7030
rect 4008 7018 5208 7028
rect 4732 6690 4788 6702
rect 4732 6638 4734 6690
rect 4786 6638 4788 6690
rect 3948 6578 4004 6590
rect 3948 6526 3950 6578
rect 4002 6526 4004 6578
rect 3948 6356 4004 6526
rect 3948 6290 4004 6300
rect 4732 6020 4788 6638
rect 4732 5954 4788 5964
rect 4732 5796 4788 5806
rect 4732 5702 4788 5740
rect 4008 5516 5208 5526
rect 4064 5514 4112 5516
rect 4168 5514 4216 5516
rect 4076 5462 4112 5514
rect 4200 5462 4216 5514
rect 4064 5460 4112 5462
rect 4168 5460 4216 5462
rect 4272 5514 4320 5516
rect 4376 5514 4424 5516
rect 4480 5514 4528 5516
rect 4376 5462 4396 5514
rect 4480 5462 4520 5514
rect 4272 5460 4320 5462
rect 4376 5460 4424 5462
rect 4480 5460 4528 5462
rect 4584 5460 4632 5516
rect 4688 5514 4736 5516
rect 4792 5514 4840 5516
rect 4896 5514 4944 5516
rect 4696 5462 4736 5514
rect 4820 5462 4840 5514
rect 4688 5460 4736 5462
rect 4792 5460 4840 5462
rect 4896 5460 4944 5462
rect 5000 5514 5048 5516
rect 5104 5514 5152 5516
rect 5000 5462 5016 5514
rect 5104 5462 5140 5514
rect 5000 5460 5048 5462
rect 5104 5460 5152 5462
rect 4008 5450 5208 5460
rect 4620 5236 4676 5246
rect 4060 5124 4116 5134
rect 4060 5030 4116 5068
rect 4396 5124 4452 5134
rect 4396 5010 4452 5068
rect 4396 4958 4398 5010
rect 4450 4958 4452 5010
rect 4396 4946 4452 4958
rect 3052 3614 3054 3666
rect 3106 3614 3108 3666
rect 3052 3602 3108 3614
rect 3164 3724 3444 3780
rect 3500 4284 3668 4340
rect 3724 4620 3892 4676
rect 3164 3332 3220 3724
rect 3500 3668 3556 4284
rect 3276 3612 3500 3668
rect 3276 3554 3332 3612
rect 3500 3574 3556 3612
rect 3612 4116 3668 4126
rect 3276 3502 3278 3554
rect 3330 3502 3332 3554
rect 3276 3490 3332 3502
rect 3612 3442 3668 4060
rect 3724 3556 3780 4620
rect 3836 4452 3892 4462
rect 3836 4358 3892 4396
rect 4620 4338 4676 5180
rect 5068 5010 5124 5022
rect 5068 4958 5070 5010
rect 5122 4958 5124 5010
rect 4620 4286 4622 4338
rect 4674 4286 4676 4338
rect 4620 4274 4676 4286
rect 4844 4898 4900 4910
rect 4844 4846 4846 4898
rect 4898 4846 4900 4898
rect 4844 4116 4900 4846
rect 4956 4898 5012 4910
rect 4956 4846 4958 4898
rect 5010 4846 5012 4898
rect 4956 4676 5012 4846
rect 5068 4900 5124 4958
rect 5068 4834 5124 4844
rect 4956 4610 5012 4620
rect 5292 4564 5348 7980
rect 5628 6580 5684 8094
rect 5740 8036 5796 8046
rect 5740 8034 6132 8036
rect 5740 7982 5742 8034
rect 5794 7982 6132 8034
rect 5740 7980 6132 7982
rect 5740 7970 5796 7980
rect 5964 7700 6020 7710
rect 5740 6580 5796 6590
rect 5628 6578 5796 6580
rect 5628 6526 5742 6578
rect 5794 6526 5796 6578
rect 5628 6524 5796 6526
rect 5516 6468 5572 6478
rect 5516 6374 5572 6412
rect 5628 6244 5684 6524
rect 5740 6514 5796 6524
rect 5852 6578 5908 6590
rect 5852 6526 5854 6578
rect 5906 6526 5908 6578
rect 5852 6356 5908 6526
rect 5852 6290 5908 6300
rect 5180 4508 5348 4564
rect 5404 6188 5684 6244
rect 5404 5348 5460 6188
rect 5180 4116 5236 4508
rect 5404 4450 5460 5292
rect 5516 6020 5572 6030
rect 5516 5906 5572 5964
rect 5964 6018 6020 7644
rect 5964 5966 5966 6018
rect 6018 5966 6020 6018
rect 5964 5954 6020 5966
rect 6076 6020 6132 7980
rect 6300 6692 6356 8876
rect 6412 8866 6468 8876
rect 7420 8930 7476 8942
rect 7420 8878 7422 8930
rect 7474 8878 7476 8930
rect 7420 8708 7476 8878
rect 7420 8642 7476 8652
rect 7196 8596 7252 8606
rect 6524 8036 6580 8046
rect 6524 7942 6580 7980
rect 6972 8036 7028 8046
rect 6972 7942 7028 7980
rect 6524 7588 6580 7598
rect 6412 7364 6468 7374
rect 6412 7270 6468 7308
rect 6300 6636 6468 6692
rect 6188 6522 6244 6534
rect 6188 6470 6190 6522
rect 6242 6470 6244 6522
rect 6188 6244 6244 6470
rect 6300 6468 6356 6478
rect 6300 6374 6356 6412
rect 6188 6178 6244 6188
rect 6076 5964 6244 6020
rect 5516 5854 5518 5906
rect 5570 5854 5572 5906
rect 5516 5236 5572 5854
rect 6076 5796 6132 5806
rect 6076 5702 6132 5740
rect 6076 5236 6132 5246
rect 5572 5234 6132 5236
rect 5572 5182 6078 5234
rect 6130 5182 6132 5234
rect 5572 5180 6132 5182
rect 5516 5142 5572 5180
rect 6076 5170 6132 5180
rect 6188 5124 6244 5964
rect 5852 5012 5908 5022
rect 5404 4398 5406 4450
rect 5458 4398 5460 4450
rect 5404 4386 5460 4398
rect 5740 4956 5852 5012
rect 5292 4338 5348 4350
rect 5292 4286 5294 4338
rect 5346 4286 5348 4338
rect 5292 4228 5348 4286
rect 5292 4172 5460 4228
rect 5404 4116 5460 4172
rect 5180 4060 5348 4116
rect 4844 4050 4900 4060
rect 4008 3948 5208 3958
rect 4064 3946 4112 3948
rect 4168 3946 4216 3948
rect 4076 3894 4112 3946
rect 4200 3894 4216 3946
rect 4064 3892 4112 3894
rect 4168 3892 4216 3894
rect 4272 3946 4320 3948
rect 4376 3946 4424 3948
rect 4480 3946 4528 3948
rect 4376 3894 4396 3946
rect 4480 3894 4520 3946
rect 4272 3892 4320 3894
rect 4376 3892 4424 3894
rect 4480 3892 4528 3894
rect 4584 3892 4632 3948
rect 4688 3946 4736 3948
rect 4792 3946 4840 3948
rect 4896 3946 4944 3948
rect 4696 3894 4736 3946
rect 4820 3894 4840 3946
rect 4688 3892 4736 3894
rect 4792 3892 4840 3894
rect 4896 3892 4944 3894
rect 5000 3946 5048 3948
rect 5104 3946 5152 3948
rect 5000 3894 5016 3946
rect 5104 3894 5140 3946
rect 5000 3892 5048 3894
rect 5104 3892 5152 3894
rect 4008 3882 5208 3892
rect 4284 3780 4340 3790
rect 5292 3780 5348 4060
rect 5404 4050 5460 4060
rect 4060 3668 4116 3678
rect 3948 3556 4004 3566
rect 3724 3500 3948 3556
rect 3948 3462 4004 3500
rect 3612 3390 3614 3442
rect 3666 3390 3668 3442
rect 3612 3378 3668 3390
rect 3164 3276 3444 3332
rect 3388 800 3444 3276
rect 4060 980 4116 3612
rect 4284 3442 4340 3724
rect 4732 3724 5348 3780
rect 4732 3554 4788 3724
rect 4732 3502 4734 3554
rect 4786 3502 4788 3554
rect 4732 3490 4788 3502
rect 5180 3556 5236 3566
rect 4284 3390 4286 3442
rect 4338 3390 4340 3442
rect 4284 3378 4340 3390
rect 4956 3444 5012 3482
rect 4956 3378 5012 3388
rect 4060 924 4340 980
rect 4284 800 4340 924
rect 5180 800 5236 3500
rect 5292 3388 5348 3724
rect 5740 3556 5796 4956
rect 5852 4946 5908 4956
rect 6076 4452 6132 4462
rect 6188 4452 6244 5068
rect 6300 5906 6356 5918
rect 6300 5854 6302 5906
rect 6354 5854 6356 5906
rect 6300 4564 6356 5854
rect 6412 5012 6468 6636
rect 6524 6690 6580 7532
rect 7196 7474 7252 8540
rect 7420 8372 7476 8382
rect 7420 8278 7476 8316
rect 7532 7700 7588 9548
rect 7644 9538 7700 9548
rect 7868 8930 7924 8942
rect 7868 8878 7870 8930
rect 7922 8878 7924 8930
rect 7868 8708 7924 8878
rect 7868 8642 7924 8652
rect 8428 8930 8484 8942
rect 8428 8878 8430 8930
rect 8482 8878 8484 8930
rect 7756 8372 7812 8382
rect 7756 8278 7812 8316
rect 8204 8260 8260 8270
rect 8204 8146 8260 8204
rect 8204 8094 8206 8146
rect 8258 8094 8260 8146
rect 8204 8082 8260 8094
rect 8316 8146 8372 8158
rect 8316 8094 8318 8146
rect 8370 8094 8372 8146
rect 7644 8036 7700 8046
rect 7644 8034 7924 8036
rect 7644 7982 7646 8034
rect 7698 7982 7924 8034
rect 7644 7980 7924 7982
rect 7644 7970 7700 7980
rect 7532 7644 7700 7700
rect 7532 7476 7588 7486
rect 7196 7422 7198 7474
rect 7250 7422 7252 7474
rect 7196 7410 7252 7422
rect 7308 7474 7588 7476
rect 7308 7422 7534 7474
rect 7586 7422 7588 7474
rect 7308 7420 7588 7422
rect 6524 6638 6526 6690
rect 6578 6638 6580 6690
rect 6524 6626 6580 6638
rect 6748 6916 6804 6926
rect 6748 6690 6804 6860
rect 7196 6804 7252 6814
rect 7308 6804 7364 7420
rect 7532 7410 7588 7420
rect 7644 7028 7700 7644
rect 7756 7476 7812 7486
rect 7756 7382 7812 7420
rect 7196 6802 7364 6804
rect 7196 6750 7198 6802
rect 7250 6750 7364 6802
rect 7196 6748 7364 6750
rect 7532 6972 7700 7028
rect 7196 6738 7252 6748
rect 6748 6638 6750 6690
rect 6802 6638 6804 6690
rect 6748 6626 6804 6638
rect 7308 6578 7364 6590
rect 7532 6580 7588 6972
rect 7868 6804 7924 7980
rect 7980 8034 8036 8046
rect 7980 7982 7982 8034
rect 8034 7982 8036 8034
rect 7980 7700 8036 7982
rect 8316 8036 8372 8094
rect 8316 7700 8372 7980
rect 7980 7634 8036 7644
rect 8092 7644 8372 7700
rect 7980 7364 8036 7374
rect 7980 7270 8036 7308
rect 7308 6526 7310 6578
rect 7362 6526 7364 6578
rect 6636 6468 6692 6478
rect 6524 6020 6580 6030
rect 6636 6020 6692 6412
rect 7084 6466 7140 6478
rect 7084 6414 7086 6466
rect 7138 6414 7140 6466
rect 6860 6244 6916 6254
rect 6860 6130 6916 6188
rect 6860 6078 6862 6130
rect 6914 6078 6916 6130
rect 6860 6066 6916 6078
rect 6524 6018 6692 6020
rect 6524 5966 6526 6018
rect 6578 5966 6692 6018
rect 6524 5964 6692 5966
rect 7084 6020 7140 6414
rect 6524 5954 6580 5964
rect 7084 5954 7140 5964
rect 7308 6244 7364 6526
rect 6412 4946 6468 4956
rect 6972 5906 7028 5918
rect 6972 5854 6974 5906
rect 7026 5854 7028 5906
rect 6860 4900 6916 4910
rect 6300 4498 6356 4508
rect 6748 4844 6860 4900
rect 6076 4450 6244 4452
rect 6076 4398 6078 4450
rect 6130 4398 6244 4450
rect 6076 4396 6244 4398
rect 6076 4386 6132 4396
rect 6412 4340 6468 4350
rect 6412 4246 6468 4284
rect 5740 3490 5796 3500
rect 6076 3892 6132 3902
rect 6076 3442 6132 3836
rect 6076 3390 6078 3442
rect 6130 3390 6132 3442
rect 5292 3332 6020 3388
rect 6076 3378 6132 3390
rect 6524 3780 6580 3790
rect 6524 3554 6580 3724
rect 6524 3502 6526 3554
rect 6578 3502 6580 3554
rect 5964 1764 6020 3332
rect 5964 1708 6132 1764
rect 6076 800 6132 1708
rect 6524 980 6580 3502
rect 6748 3442 6804 4844
rect 6860 4834 6916 4844
rect 6860 4564 6916 4602
rect 6860 4498 6916 4508
rect 6860 4340 6916 4350
rect 6972 4340 7028 5854
rect 6860 4338 7028 4340
rect 6860 4286 6862 4338
rect 6914 4286 7028 4338
rect 6860 4284 7028 4286
rect 7084 5684 7140 5694
rect 6860 4116 6916 4284
rect 6860 4050 6916 4060
rect 7084 4114 7140 5628
rect 7308 4676 7364 6188
rect 7420 6524 7588 6580
rect 7644 6748 7924 6804
rect 7420 6018 7476 6524
rect 7644 6244 7700 6748
rect 7980 6692 8036 6702
rect 7420 5966 7422 6018
rect 7474 5966 7476 6018
rect 7420 5954 7476 5966
rect 7532 6188 7700 6244
rect 7756 6466 7812 6478
rect 7756 6414 7758 6466
rect 7810 6414 7812 6466
rect 7756 6244 7812 6414
rect 7868 6468 7924 6478
rect 7868 6374 7924 6412
rect 7980 6466 8036 6636
rect 7980 6414 7982 6466
rect 8034 6414 8036 6466
rect 7980 6402 8036 6414
rect 8092 6244 8148 7644
rect 8204 7476 8260 7486
rect 8204 7382 8260 7420
rect 8316 7364 8372 7374
rect 8204 6468 8260 6478
rect 8204 6374 8260 6412
rect 7308 4610 7364 4620
rect 7420 4452 7476 4462
rect 7532 4452 7588 6188
rect 7756 6178 7812 6188
rect 7868 6188 8148 6244
rect 7420 4450 7588 4452
rect 7420 4398 7422 4450
rect 7474 4398 7588 4450
rect 7420 4396 7588 4398
rect 7644 6020 7700 6030
rect 7644 4452 7700 5964
rect 7756 5908 7812 5918
rect 7756 4564 7812 5852
rect 7868 4676 7924 6188
rect 8092 6020 8148 6030
rect 8092 6018 8260 6020
rect 8092 5966 8094 6018
rect 8146 5966 8260 6018
rect 8092 5964 8260 5966
rect 8092 5954 8148 5964
rect 8204 5908 8260 5964
rect 8316 5908 8372 7308
rect 8204 5852 8372 5908
rect 7980 5794 8036 5806
rect 7980 5742 7982 5794
rect 8034 5742 8036 5794
rect 7980 4900 8036 5742
rect 7980 4834 8036 4844
rect 7868 4620 8260 4676
rect 7756 4508 8148 4564
rect 7644 4450 8036 4452
rect 7644 4398 7646 4450
rect 7698 4398 8036 4450
rect 7644 4396 8036 4398
rect 7420 4386 7476 4396
rect 7644 4386 7700 4396
rect 7980 4338 8036 4396
rect 8092 4450 8148 4508
rect 8204 4562 8260 4620
rect 8204 4510 8206 4562
rect 8258 4510 8260 4562
rect 8204 4498 8260 4510
rect 8428 4452 8484 8878
rect 8764 8930 8820 8942
rect 8764 8878 8766 8930
rect 8818 8878 8820 8930
rect 8764 8260 8820 8878
rect 8764 8194 8820 8204
rect 8876 8932 8932 8942
rect 8764 8034 8820 8046
rect 8764 7982 8766 8034
rect 8818 7982 8820 8034
rect 8652 7476 8708 7486
rect 8652 7382 8708 7420
rect 8764 6804 8820 7982
rect 8876 7698 8932 8876
rect 9660 8932 9716 8942
rect 9660 8838 9716 8876
rect 9772 8596 9828 9774
rect 10220 9044 10276 9054
rect 10332 9044 10388 10556
rect 11900 10612 11956 10622
rect 11900 10518 11956 10556
rect 12124 10612 12180 10622
rect 12124 10518 12180 10556
rect 12572 10612 12628 10622
rect 12908 10612 12964 10622
rect 12572 10610 12740 10612
rect 12572 10558 12574 10610
rect 12626 10558 12740 10610
rect 12572 10556 12740 10558
rect 12572 10546 12628 10556
rect 10780 10500 10836 10510
rect 10556 9716 10612 9726
rect 10444 9714 10612 9716
rect 10444 9662 10558 9714
rect 10610 9662 10612 9714
rect 10444 9660 10612 9662
rect 10444 9266 10500 9660
rect 10556 9650 10612 9660
rect 10444 9214 10446 9266
rect 10498 9214 10500 9266
rect 10444 9202 10500 9214
rect 10780 9154 10836 10444
rect 12012 10500 12068 10510
rect 12012 10406 12068 10444
rect 12684 10386 12740 10556
rect 12684 10334 12686 10386
rect 12738 10334 12740 10386
rect 12684 10322 12740 10334
rect 10780 9102 10782 9154
rect 10834 9102 10836 9154
rect 10780 9090 10836 9102
rect 12684 9940 12740 9950
rect 12908 9940 12964 10556
rect 12684 9938 12964 9940
rect 12684 9886 12686 9938
rect 12738 9886 12964 9938
rect 12684 9884 12964 9886
rect 13356 10498 13412 10510
rect 13356 10446 13358 10498
rect 13410 10446 13412 10498
rect 13356 10386 13412 10446
rect 13356 10334 13358 10386
rect 13410 10334 13412 10386
rect 10220 9042 10388 9044
rect 10220 8990 10222 9042
rect 10274 8990 10388 9042
rect 10220 8988 10388 8990
rect 10220 8978 10276 8988
rect 9772 8530 9828 8540
rect 9324 8148 9380 8158
rect 8876 7646 8878 7698
rect 8930 7646 8932 7698
rect 8876 7634 8932 7646
rect 8988 8036 9044 8046
rect 9212 8036 9268 8046
rect 9044 8034 9268 8036
rect 9044 7982 9214 8034
rect 9266 7982 9268 8034
rect 9044 7980 9268 7982
rect 8988 7586 9044 7980
rect 9212 7970 9268 7980
rect 8988 7534 8990 7586
rect 9042 7534 9044 7586
rect 8988 7522 9044 7534
rect 8764 6748 8932 6804
rect 8652 6580 8708 6590
rect 8652 6486 8708 6524
rect 8876 6020 8932 6748
rect 8764 5964 8932 6020
rect 8988 6132 9044 6142
rect 8988 6018 9044 6076
rect 8988 5966 8990 6018
rect 9042 5966 9044 6018
rect 8540 5908 8596 5918
rect 8540 5814 8596 5852
rect 8652 5906 8708 5918
rect 8652 5854 8654 5906
rect 8706 5854 8708 5906
rect 8652 5124 8708 5854
rect 8652 5058 8708 5068
rect 8092 4398 8094 4450
rect 8146 4398 8148 4450
rect 8092 4386 8148 4398
rect 8316 4396 8484 4452
rect 7980 4286 7982 4338
rect 8034 4286 8036 4338
rect 7980 4274 8036 4286
rect 7084 4062 7086 4114
rect 7138 4062 7140 4114
rect 7084 4050 7140 4062
rect 8092 4004 8148 4014
rect 7868 3780 7924 3790
rect 6748 3390 6750 3442
rect 6802 3390 6804 3442
rect 6748 3378 6804 3390
rect 6972 3556 7028 3566
rect 6524 914 6580 924
rect 6972 800 7028 3500
rect 7420 3556 7476 3566
rect 7420 3442 7476 3500
rect 7868 3554 7924 3724
rect 7868 3502 7870 3554
rect 7922 3502 7924 3554
rect 7868 3490 7924 3502
rect 7420 3390 7422 3442
rect 7474 3390 7476 3442
rect 7420 3378 7476 3390
rect 8092 3442 8148 3948
rect 8316 3780 8372 4396
rect 8764 4340 8820 5964
rect 8988 5954 9044 5966
rect 8876 5794 8932 5806
rect 8876 5742 8878 5794
rect 8930 5742 8932 5794
rect 8876 5684 8932 5742
rect 9324 5684 9380 8092
rect 9660 8146 9716 8158
rect 9660 8094 9662 8146
rect 9714 8094 9716 8146
rect 8876 5628 9380 5684
rect 9436 6580 9492 6590
rect 8652 4338 8820 4340
rect 8652 4286 8766 4338
rect 8818 4286 8820 4338
rect 8652 4284 8820 4286
rect 8316 3714 8372 3724
rect 8428 4228 8484 4238
rect 8428 3554 8484 4172
rect 8428 3502 8430 3554
rect 8482 3502 8484 3554
rect 8428 3490 8484 3502
rect 8092 3390 8094 3442
rect 8146 3390 8148 3442
rect 8092 3378 8148 3390
rect 7084 3332 7140 3342
rect 7084 2994 7140 3276
rect 7084 2942 7086 2994
rect 7138 2942 7140 2994
rect 7084 2930 7140 2942
rect 8652 1764 8708 4284
rect 8764 4274 8820 4284
rect 8876 5236 8932 5246
rect 9436 5236 9492 6524
rect 9660 5348 9716 8094
rect 10108 7588 10164 7598
rect 10108 7494 10164 7532
rect 9660 5282 9716 5292
rect 9772 7362 9828 7374
rect 9772 7310 9774 7362
rect 9826 7310 9828 7362
rect 8764 3444 8820 3454
rect 8876 3444 8932 5180
rect 8988 5180 9492 5236
rect 8988 4562 9044 5180
rect 8988 4510 8990 4562
rect 9042 4510 9044 4562
rect 8988 4498 9044 4510
rect 9324 3666 9380 5180
rect 9436 4900 9492 4910
rect 9436 3778 9492 4844
rect 9436 3726 9438 3778
rect 9490 3726 9492 3778
rect 9436 3714 9492 3726
rect 9324 3614 9326 3666
rect 9378 3614 9380 3666
rect 9324 3602 9380 3614
rect 9772 3556 9828 7310
rect 10220 6692 10276 6702
rect 9996 6690 10276 6692
rect 9996 6638 10222 6690
rect 10274 6638 10276 6690
rect 9996 6636 10276 6638
rect 9884 4788 9940 4798
rect 9884 4562 9940 4732
rect 9884 4510 9886 4562
rect 9938 4510 9940 4562
rect 9884 4498 9940 4510
rect 9884 4338 9940 4350
rect 9884 4286 9886 4338
rect 9938 4286 9940 4338
rect 9884 4116 9940 4286
rect 9884 4050 9940 4060
rect 9996 4226 10052 6636
rect 10220 6626 10276 6636
rect 10220 6132 10276 6142
rect 10332 6132 10388 8988
rect 10444 9042 10500 9054
rect 10444 8990 10446 9042
rect 10498 8990 10500 9042
rect 10444 7364 10500 8990
rect 11340 9042 11396 9054
rect 11340 8990 11342 9042
rect 11394 8990 11396 9042
rect 10444 7298 10500 7308
rect 10780 8258 10836 8270
rect 10780 8206 10782 8258
rect 10834 8206 10836 8258
rect 10780 7140 10836 8206
rect 10780 7074 10836 7084
rect 10276 6076 10388 6132
rect 10668 6690 10724 6702
rect 10668 6638 10670 6690
rect 10722 6638 10724 6690
rect 10220 6066 10276 6076
rect 10220 5012 10276 5022
rect 9996 4174 9998 4226
rect 10050 4174 10052 4226
rect 9772 3462 9828 3500
rect 9884 3780 9940 3790
rect 8764 3442 8932 3444
rect 8764 3390 8766 3442
rect 8818 3390 8932 3442
rect 8764 3388 8932 3390
rect 9884 3388 9940 3724
rect 9996 3668 10052 4174
rect 10108 4956 10220 5012
rect 10108 4338 10164 4956
rect 10220 4946 10276 4956
rect 10108 4286 10110 4338
rect 10162 4286 10164 4338
rect 10108 3892 10164 4286
rect 10108 3826 10164 3836
rect 10220 4676 10276 4686
rect 9996 3602 10052 3612
rect 10108 3444 10164 3454
rect 10220 3444 10276 4620
rect 10668 4116 10724 6638
rect 10668 4050 10724 4060
rect 10780 6692 10836 6702
rect 10556 3668 10612 3678
rect 10556 3554 10612 3612
rect 10556 3502 10558 3554
rect 10610 3502 10612 3554
rect 10556 3490 10612 3502
rect 10108 3442 10276 3444
rect 10108 3390 10110 3442
rect 10162 3390 10276 3442
rect 10108 3388 10276 3390
rect 10780 3442 10836 6636
rect 10892 6636 11284 6692
rect 10892 5012 10948 6636
rect 11228 6578 11284 6636
rect 11228 6526 11230 6578
rect 11282 6526 11284 6578
rect 11228 6514 11284 6526
rect 11116 6468 11172 6478
rect 10892 4946 10948 4956
rect 11004 6466 11172 6468
rect 11004 6414 11118 6466
rect 11170 6414 11172 6466
rect 11004 6412 11172 6414
rect 11004 3556 11060 6412
rect 11116 6402 11172 6412
rect 11340 6020 11396 8990
rect 12684 8932 12740 9884
rect 12684 8866 12740 8876
rect 11564 8260 11620 8270
rect 11564 7476 11620 8204
rect 12796 8258 12852 8270
rect 12796 8206 12798 8258
rect 12850 8206 12852 8258
rect 11564 6916 11620 7420
rect 11676 7474 11732 7486
rect 11676 7422 11678 7474
rect 11730 7422 11732 7474
rect 11676 7140 11732 7422
rect 11676 7074 11732 7084
rect 11788 7362 11844 7374
rect 11788 7310 11790 7362
rect 11842 7310 11844 7362
rect 11564 6860 11732 6916
rect 11116 6018 11396 6020
rect 11116 5966 11342 6018
rect 11394 5966 11396 6018
rect 11116 5964 11396 5966
rect 11116 5122 11172 5964
rect 11340 5954 11396 5964
rect 11452 6132 11508 6142
rect 11116 5070 11118 5122
rect 11170 5070 11172 5122
rect 11116 5058 11172 5070
rect 11228 5124 11284 5134
rect 11116 4564 11172 4574
rect 11228 4564 11284 5068
rect 11116 4562 11284 4564
rect 11116 4510 11118 4562
rect 11170 4510 11284 4562
rect 11116 4508 11284 4510
rect 11452 4898 11508 6076
rect 11564 5908 11620 5918
rect 11564 5234 11620 5852
rect 11564 5182 11566 5234
rect 11618 5182 11620 5234
rect 11564 5170 11620 5182
rect 11676 5010 11732 6860
rect 11788 6020 11844 7310
rect 12796 7364 12852 8206
rect 12908 8146 12964 8158
rect 12908 8094 12910 8146
rect 12962 8094 12964 8146
rect 12908 7588 12964 8094
rect 13132 7588 13188 7598
rect 12908 7586 13188 7588
rect 12908 7534 13134 7586
rect 13186 7534 13188 7586
rect 12908 7532 13188 7534
rect 12908 7364 12964 7374
rect 12796 7308 12908 7364
rect 12908 7298 12964 7308
rect 11788 5954 11844 5964
rect 12124 6580 12180 6590
rect 12124 5122 12180 6524
rect 13020 6466 13076 6478
rect 13020 6414 13022 6466
rect 13074 6414 13076 6466
rect 12124 5070 12126 5122
rect 12178 5070 12180 5122
rect 12124 5058 12180 5070
rect 12236 5348 12292 5358
rect 12236 5122 12292 5292
rect 12236 5070 12238 5122
rect 12290 5070 12292 5122
rect 12236 5058 12292 5070
rect 11676 4958 11678 5010
rect 11730 4958 11732 5010
rect 11676 4946 11732 4958
rect 12572 5010 12628 5022
rect 12572 4958 12574 5010
rect 12626 4958 12628 5010
rect 11452 4846 11454 4898
rect 11506 4846 11508 4898
rect 11452 4564 11508 4846
rect 12460 4900 12516 4910
rect 12460 4806 12516 4844
rect 12572 4788 12628 4958
rect 12572 4722 12628 4732
rect 11676 4564 11732 4574
rect 11452 4562 11732 4564
rect 11452 4510 11678 4562
rect 11730 4510 11732 4562
rect 11452 4508 11732 4510
rect 11116 4498 11172 4508
rect 11676 4498 11732 4508
rect 12124 4450 12180 4462
rect 12124 4398 12126 4450
rect 12178 4398 12180 4450
rect 11564 4340 11620 4350
rect 11452 4338 11620 4340
rect 11452 4286 11566 4338
rect 11618 4286 11620 4338
rect 11452 4284 11620 4286
rect 11228 4226 11284 4238
rect 11228 4174 11230 4226
rect 11282 4174 11284 4226
rect 11116 3556 11172 3566
rect 11004 3554 11172 3556
rect 11004 3502 11118 3554
rect 11170 3502 11172 3554
rect 11004 3500 11172 3502
rect 11116 3490 11172 3500
rect 10780 3390 10782 3442
rect 10834 3390 10836 3442
rect 8764 3378 8820 3388
rect 9884 3332 10052 3388
rect 10108 3378 10164 3388
rect 10780 3378 10836 3390
rect 11228 3444 11284 4174
rect 11452 3778 11508 4284
rect 11564 4274 11620 4284
rect 12012 4340 12068 4350
rect 12124 4340 12180 4398
rect 12068 4284 12180 4340
rect 12012 4274 12068 4284
rect 11452 3726 11454 3778
rect 11506 3726 11508 3778
rect 11452 3714 11508 3726
rect 12348 4228 12404 4238
rect 11228 3378 11284 3388
rect 11452 3556 11508 3566
rect 9996 3220 10052 3332
rect 9996 3164 10612 3220
rect 9660 2994 9716 3006
rect 9660 2942 9662 2994
rect 9714 2942 9716 2994
rect 8652 1708 8820 1764
rect 7868 980 7924 990
rect 7868 800 7924 924
rect 8764 800 8820 1708
rect 9660 800 9716 2942
rect 10556 800 10612 3164
rect 11452 800 11508 3500
rect 11676 3556 11732 3566
rect 11676 3462 11732 3500
rect 12348 800 12404 4172
rect 12572 3780 12628 3790
rect 12572 3554 12628 3724
rect 12572 3502 12574 3554
rect 12626 3502 12628 3554
rect 12572 3490 12628 3502
rect 13020 3668 13076 6414
rect 13132 6356 13188 7532
rect 13356 6580 13412 10334
rect 13692 9604 13748 9614
rect 13580 9602 13748 9604
rect 13580 9550 13694 9602
rect 13746 9550 13748 9602
rect 13580 9548 13748 9550
rect 13468 8930 13524 8942
rect 13468 8878 13470 8930
rect 13522 8878 13524 8930
rect 13468 8596 13524 8878
rect 13468 8258 13524 8540
rect 13468 8206 13470 8258
rect 13522 8206 13524 8258
rect 13468 8194 13524 8206
rect 13580 7140 13636 9548
rect 13692 9538 13748 9548
rect 13804 7588 13860 45836
rect 14140 45826 14196 45836
rect 14812 45826 14868 45836
rect 17500 45780 17556 49200
rect 17724 45780 17780 45790
rect 17500 45778 17780 45780
rect 17500 45726 17726 45778
rect 17778 45726 17780 45778
rect 17500 45724 17780 45726
rect 22428 45780 22484 49200
rect 24008 46284 25208 46294
rect 24064 46282 24112 46284
rect 24168 46282 24216 46284
rect 24076 46230 24112 46282
rect 24200 46230 24216 46282
rect 24064 46228 24112 46230
rect 24168 46228 24216 46230
rect 24272 46282 24320 46284
rect 24376 46282 24424 46284
rect 24480 46282 24528 46284
rect 24376 46230 24396 46282
rect 24480 46230 24520 46282
rect 24272 46228 24320 46230
rect 24376 46228 24424 46230
rect 24480 46228 24528 46230
rect 24584 46228 24632 46284
rect 24688 46282 24736 46284
rect 24792 46282 24840 46284
rect 24896 46282 24944 46284
rect 24696 46230 24736 46282
rect 24820 46230 24840 46282
rect 24688 46228 24736 46230
rect 24792 46228 24840 46230
rect 24896 46228 24944 46230
rect 25000 46282 25048 46284
rect 25104 46282 25152 46284
rect 25000 46230 25016 46282
rect 25104 46230 25140 46282
rect 25000 46228 25048 46230
rect 25104 46228 25152 46230
rect 24008 46218 25208 46228
rect 27356 46116 27412 49200
rect 27356 46050 27412 46060
rect 28812 46116 28868 46126
rect 28812 46002 28868 46060
rect 28812 45950 28814 46002
rect 28866 45950 28868 46002
rect 28812 45938 28868 45950
rect 22652 45780 22708 45790
rect 22428 45778 22708 45780
rect 22428 45726 22654 45778
rect 22706 45726 22708 45778
rect 22428 45724 22708 45726
rect 32284 45780 32340 49200
rect 37212 46562 37268 49200
rect 37212 46510 37214 46562
rect 37266 46510 37268 46562
rect 37212 46498 37268 46510
rect 37884 46562 37940 46574
rect 37884 46510 37886 46562
rect 37938 46510 37940 46562
rect 37884 46002 37940 46510
rect 37884 45950 37886 46002
rect 37938 45950 37940 46002
rect 37884 45938 37940 45950
rect 32508 45780 32564 45790
rect 32284 45778 32564 45780
rect 32284 45726 32510 45778
rect 32562 45726 32564 45778
rect 32284 45724 32564 45726
rect 17724 45714 17780 45724
rect 22652 45714 22708 45724
rect 32508 45714 32564 45724
rect 27916 45668 27972 45678
rect 28364 45668 28420 45678
rect 27916 45666 28420 45668
rect 27916 45614 27918 45666
rect 27970 45614 28366 45666
rect 28418 45614 28420 45666
rect 27916 45612 28420 45614
rect 27916 45602 27972 45612
rect 14008 45500 15208 45510
rect 14064 45498 14112 45500
rect 14168 45498 14216 45500
rect 14076 45446 14112 45498
rect 14200 45446 14216 45498
rect 14064 45444 14112 45446
rect 14168 45444 14216 45446
rect 14272 45498 14320 45500
rect 14376 45498 14424 45500
rect 14480 45498 14528 45500
rect 14376 45446 14396 45498
rect 14480 45446 14520 45498
rect 14272 45444 14320 45446
rect 14376 45444 14424 45446
rect 14480 45444 14528 45446
rect 14584 45444 14632 45500
rect 14688 45498 14736 45500
rect 14792 45498 14840 45500
rect 14896 45498 14944 45500
rect 14696 45446 14736 45498
rect 14820 45446 14840 45498
rect 14688 45444 14736 45446
rect 14792 45444 14840 45446
rect 14896 45444 14944 45446
rect 15000 45498 15048 45500
rect 15104 45498 15152 45500
rect 15000 45446 15016 45498
rect 15104 45446 15140 45498
rect 15000 45444 15048 45446
rect 15104 45444 15152 45446
rect 14008 45434 15208 45444
rect 24008 44716 25208 44726
rect 24064 44714 24112 44716
rect 24168 44714 24216 44716
rect 24076 44662 24112 44714
rect 24200 44662 24216 44714
rect 24064 44660 24112 44662
rect 24168 44660 24216 44662
rect 24272 44714 24320 44716
rect 24376 44714 24424 44716
rect 24480 44714 24528 44716
rect 24376 44662 24396 44714
rect 24480 44662 24520 44714
rect 24272 44660 24320 44662
rect 24376 44660 24424 44662
rect 24480 44660 24528 44662
rect 24584 44660 24632 44716
rect 24688 44714 24736 44716
rect 24792 44714 24840 44716
rect 24896 44714 24944 44716
rect 24696 44662 24736 44714
rect 24820 44662 24840 44714
rect 24688 44660 24736 44662
rect 24792 44660 24840 44662
rect 24896 44660 24944 44662
rect 25000 44714 25048 44716
rect 25104 44714 25152 44716
rect 25000 44662 25016 44714
rect 25104 44662 25140 44714
rect 25000 44660 25048 44662
rect 25104 44660 25152 44662
rect 24008 44650 25208 44660
rect 14008 43932 15208 43942
rect 14064 43930 14112 43932
rect 14168 43930 14216 43932
rect 14076 43878 14112 43930
rect 14200 43878 14216 43930
rect 14064 43876 14112 43878
rect 14168 43876 14216 43878
rect 14272 43930 14320 43932
rect 14376 43930 14424 43932
rect 14480 43930 14528 43932
rect 14376 43878 14396 43930
rect 14480 43878 14520 43930
rect 14272 43876 14320 43878
rect 14376 43876 14424 43878
rect 14480 43876 14528 43878
rect 14584 43876 14632 43932
rect 14688 43930 14736 43932
rect 14792 43930 14840 43932
rect 14896 43930 14944 43932
rect 14696 43878 14736 43930
rect 14820 43878 14840 43930
rect 14688 43876 14736 43878
rect 14792 43876 14840 43878
rect 14896 43876 14944 43878
rect 15000 43930 15048 43932
rect 15104 43930 15152 43932
rect 15000 43878 15016 43930
rect 15104 43878 15140 43930
rect 15000 43876 15048 43878
rect 15104 43876 15152 43878
rect 14008 43866 15208 43876
rect 24008 43148 25208 43158
rect 24064 43146 24112 43148
rect 24168 43146 24216 43148
rect 24076 43094 24112 43146
rect 24200 43094 24216 43146
rect 24064 43092 24112 43094
rect 24168 43092 24216 43094
rect 24272 43146 24320 43148
rect 24376 43146 24424 43148
rect 24480 43146 24528 43148
rect 24376 43094 24396 43146
rect 24480 43094 24520 43146
rect 24272 43092 24320 43094
rect 24376 43092 24424 43094
rect 24480 43092 24528 43094
rect 24584 43092 24632 43148
rect 24688 43146 24736 43148
rect 24792 43146 24840 43148
rect 24896 43146 24944 43148
rect 24696 43094 24736 43146
rect 24820 43094 24840 43146
rect 24688 43092 24736 43094
rect 24792 43092 24840 43094
rect 24896 43092 24944 43094
rect 25000 43146 25048 43148
rect 25104 43146 25152 43148
rect 25000 43094 25016 43146
rect 25104 43094 25140 43146
rect 25000 43092 25048 43094
rect 25104 43092 25152 43094
rect 24008 43082 25208 43092
rect 14008 42364 15208 42374
rect 14064 42362 14112 42364
rect 14168 42362 14216 42364
rect 14076 42310 14112 42362
rect 14200 42310 14216 42362
rect 14064 42308 14112 42310
rect 14168 42308 14216 42310
rect 14272 42362 14320 42364
rect 14376 42362 14424 42364
rect 14480 42362 14528 42364
rect 14376 42310 14396 42362
rect 14480 42310 14520 42362
rect 14272 42308 14320 42310
rect 14376 42308 14424 42310
rect 14480 42308 14528 42310
rect 14584 42308 14632 42364
rect 14688 42362 14736 42364
rect 14792 42362 14840 42364
rect 14896 42362 14944 42364
rect 14696 42310 14736 42362
rect 14820 42310 14840 42362
rect 14688 42308 14736 42310
rect 14792 42308 14840 42310
rect 14896 42308 14944 42310
rect 15000 42362 15048 42364
rect 15104 42362 15152 42364
rect 15000 42310 15016 42362
rect 15104 42310 15140 42362
rect 15000 42308 15048 42310
rect 15104 42308 15152 42310
rect 14008 42298 15208 42308
rect 24008 41580 25208 41590
rect 24064 41578 24112 41580
rect 24168 41578 24216 41580
rect 24076 41526 24112 41578
rect 24200 41526 24216 41578
rect 24064 41524 24112 41526
rect 24168 41524 24216 41526
rect 24272 41578 24320 41580
rect 24376 41578 24424 41580
rect 24480 41578 24528 41580
rect 24376 41526 24396 41578
rect 24480 41526 24520 41578
rect 24272 41524 24320 41526
rect 24376 41524 24424 41526
rect 24480 41524 24528 41526
rect 24584 41524 24632 41580
rect 24688 41578 24736 41580
rect 24792 41578 24840 41580
rect 24896 41578 24944 41580
rect 24696 41526 24736 41578
rect 24820 41526 24840 41578
rect 24688 41524 24736 41526
rect 24792 41524 24840 41526
rect 24896 41524 24944 41526
rect 25000 41578 25048 41580
rect 25104 41578 25152 41580
rect 25000 41526 25016 41578
rect 25104 41526 25140 41578
rect 25000 41524 25048 41526
rect 25104 41524 25152 41526
rect 24008 41514 25208 41524
rect 14008 40796 15208 40806
rect 14064 40794 14112 40796
rect 14168 40794 14216 40796
rect 14076 40742 14112 40794
rect 14200 40742 14216 40794
rect 14064 40740 14112 40742
rect 14168 40740 14216 40742
rect 14272 40794 14320 40796
rect 14376 40794 14424 40796
rect 14480 40794 14528 40796
rect 14376 40742 14396 40794
rect 14480 40742 14520 40794
rect 14272 40740 14320 40742
rect 14376 40740 14424 40742
rect 14480 40740 14528 40742
rect 14584 40740 14632 40796
rect 14688 40794 14736 40796
rect 14792 40794 14840 40796
rect 14896 40794 14944 40796
rect 14696 40742 14736 40794
rect 14820 40742 14840 40794
rect 14688 40740 14736 40742
rect 14792 40740 14840 40742
rect 14896 40740 14944 40742
rect 15000 40794 15048 40796
rect 15104 40794 15152 40796
rect 15000 40742 15016 40794
rect 15104 40742 15140 40794
rect 15000 40740 15048 40742
rect 15104 40740 15152 40742
rect 14008 40730 15208 40740
rect 24008 40012 25208 40022
rect 24064 40010 24112 40012
rect 24168 40010 24216 40012
rect 24076 39958 24112 40010
rect 24200 39958 24216 40010
rect 24064 39956 24112 39958
rect 24168 39956 24216 39958
rect 24272 40010 24320 40012
rect 24376 40010 24424 40012
rect 24480 40010 24528 40012
rect 24376 39958 24396 40010
rect 24480 39958 24520 40010
rect 24272 39956 24320 39958
rect 24376 39956 24424 39958
rect 24480 39956 24528 39958
rect 24584 39956 24632 40012
rect 24688 40010 24736 40012
rect 24792 40010 24840 40012
rect 24896 40010 24944 40012
rect 24696 39958 24736 40010
rect 24820 39958 24840 40010
rect 24688 39956 24736 39958
rect 24792 39956 24840 39958
rect 24896 39956 24944 39958
rect 25000 40010 25048 40012
rect 25104 40010 25152 40012
rect 25000 39958 25016 40010
rect 25104 39958 25140 40010
rect 25000 39956 25048 39958
rect 25104 39956 25152 39958
rect 24008 39946 25208 39956
rect 14008 39228 15208 39238
rect 14064 39226 14112 39228
rect 14168 39226 14216 39228
rect 14076 39174 14112 39226
rect 14200 39174 14216 39226
rect 14064 39172 14112 39174
rect 14168 39172 14216 39174
rect 14272 39226 14320 39228
rect 14376 39226 14424 39228
rect 14480 39226 14528 39228
rect 14376 39174 14396 39226
rect 14480 39174 14520 39226
rect 14272 39172 14320 39174
rect 14376 39172 14424 39174
rect 14480 39172 14528 39174
rect 14584 39172 14632 39228
rect 14688 39226 14736 39228
rect 14792 39226 14840 39228
rect 14896 39226 14944 39228
rect 14696 39174 14736 39226
rect 14820 39174 14840 39226
rect 14688 39172 14736 39174
rect 14792 39172 14840 39174
rect 14896 39172 14944 39174
rect 15000 39226 15048 39228
rect 15104 39226 15152 39228
rect 15000 39174 15016 39226
rect 15104 39174 15140 39226
rect 15000 39172 15048 39174
rect 15104 39172 15152 39174
rect 14008 39162 15208 39172
rect 24008 38444 25208 38454
rect 24064 38442 24112 38444
rect 24168 38442 24216 38444
rect 24076 38390 24112 38442
rect 24200 38390 24216 38442
rect 24064 38388 24112 38390
rect 24168 38388 24216 38390
rect 24272 38442 24320 38444
rect 24376 38442 24424 38444
rect 24480 38442 24528 38444
rect 24376 38390 24396 38442
rect 24480 38390 24520 38442
rect 24272 38388 24320 38390
rect 24376 38388 24424 38390
rect 24480 38388 24528 38390
rect 24584 38388 24632 38444
rect 24688 38442 24736 38444
rect 24792 38442 24840 38444
rect 24896 38442 24944 38444
rect 24696 38390 24736 38442
rect 24820 38390 24840 38442
rect 24688 38388 24736 38390
rect 24792 38388 24840 38390
rect 24896 38388 24944 38390
rect 25000 38442 25048 38444
rect 25104 38442 25152 38444
rect 25000 38390 25016 38442
rect 25104 38390 25140 38442
rect 25000 38388 25048 38390
rect 25104 38388 25152 38390
rect 24008 38378 25208 38388
rect 14008 37660 15208 37670
rect 14064 37658 14112 37660
rect 14168 37658 14216 37660
rect 14076 37606 14112 37658
rect 14200 37606 14216 37658
rect 14064 37604 14112 37606
rect 14168 37604 14216 37606
rect 14272 37658 14320 37660
rect 14376 37658 14424 37660
rect 14480 37658 14528 37660
rect 14376 37606 14396 37658
rect 14480 37606 14520 37658
rect 14272 37604 14320 37606
rect 14376 37604 14424 37606
rect 14480 37604 14528 37606
rect 14584 37604 14632 37660
rect 14688 37658 14736 37660
rect 14792 37658 14840 37660
rect 14896 37658 14944 37660
rect 14696 37606 14736 37658
rect 14820 37606 14840 37658
rect 14688 37604 14736 37606
rect 14792 37604 14840 37606
rect 14896 37604 14944 37606
rect 15000 37658 15048 37660
rect 15104 37658 15152 37660
rect 15000 37606 15016 37658
rect 15104 37606 15140 37658
rect 15000 37604 15048 37606
rect 15104 37604 15152 37606
rect 14008 37594 15208 37604
rect 24008 36876 25208 36886
rect 24064 36874 24112 36876
rect 24168 36874 24216 36876
rect 24076 36822 24112 36874
rect 24200 36822 24216 36874
rect 24064 36820 24112 36822
rect 24168 36820 24216 36822
rect 24272 36874 24320 36876
rect 24376 36874 24424 36876
rect 24480 36874 24528 36876
rect 24376 36822 24396 36874
rect 24480 36822 24520 36874
rect 24272 36820 24320 36822
rect 24376 36820 24424 36822
rect 24480 36820 24528 36822
rect 24584 36820 24632 36876
rect 24688 36874 24736 36876
rect 24792 36874 24840 36876
rect 24896 36874 24944 36876
rect 24696 36822 24736 36874
rect 24820 36822 24840 36874
rect 24688 36820 24736 36822
rect 24792 36820 24840 36822
rect 24896 36820 24944 36822
rect 25000 36874 25048 36876
rect 25104 36874 25152 36876
rect 25000 36822 25016 36874
rect 25104 36822 25140 36874
rect 25000 36820 25048 36822
rect 25104 36820 25152 36822
rect 24008 36810 25208 36820
rect 14008 36092 15208 36102
rect 14064 36090 14112 36092
rect 14168 36090 14216 36092
rect 14076 36038 14112 36090
rect 14200 36038 14216 36090
rect 14064 36036 14112 36038
rect 14168 36036 14216 36038
rect 14272 36090 14320 36092
rect 14376 36090 14424 36092
rect 14480 36090 14528 36092
rect 14376 36038 14396 36090
rect 14480 36038 14520 36090
rect 14272 36036 14320 36038
rect 14376 36036 14424 36038
rect 14480 36036 14528 36038
rect 14584 36036 14632 36092
rect 14688 36090 14736 36092
rect 14792 36090 14840 36092
rect 14896 36090 14944 36092
rect 14696 36038 14736 36090
rect 14820 36038 14840 36090
rect 14688 36036 14736 36038
rect 14792 36036 14840 36038
rect 14896 36036 14944 36038
rect 15000 36090 15048 36092
rect 15104 36090 15152 36092
rect 15000 36038 15016 36090
rect 15104 36038 15140 36090
rect 15000 36036 15048 36038
rect 15104 36036 15152 36038
rect 14008 36026 15208 36036
rect 24008 35308 25208 35318
rect 24064 35306 24112 35308
rect 24168 35306 24216 35308
rect 24076 35254 24112 35306
rect 24200 35254 24216 35306
rect 24064 35252 24112 35254
rect 24168 35252 24216 35254
rect 24272 35306 24320 35308
rect 24376 35306 24424 35308
rect 24480 35306 24528 35308
rect 24376 35254 24396 35306
rect 24480 35254 24520 35306
rect 24272 35252 24320 35254
rect 24376 35252 24424 35254
rect 24480 35252 24528 35254
rect 24584 35252 24632 35308
rect 24688 35306 24736 35308
rect 24792 35306 24840 35308
rect 24896 35306 24944 35308
rect 24696 35254 24736 35306
rect 24820 35254 24840 35306
rect 24688 35252 24736 35254
rect 24792 35252 24840 35254
rect 24896 35252 24944 35254
rect 25000 35306 25048 35308
rect 25104 35306 25152 35308
rect 25000 35254 25016 35306
rect 25104 35254 25140 35306
rect 25000 35252 25048 35254
rect 25104 35252 25152 35254
rect 24008 35242 25208 35252
rect 14008 34524 15208 34534
rect 14064 34522 14112 34524
rect 14168 34522 14216 34524
rect 14076 34470 14112 34522
rect 14200 34470 14216 34522
rect 14064 34468 14112 34470
rect 14168 34468 14216 34470
rect 14272 34522 14320 34524
rect 14376 34522 14424 34524
rect 14480 34522 14528 34524
rect 14376 34470 14396 34522
rect 14480 34470 14520 34522
rect 14272 34468 14320 34470
rect 14376 34468 14424 34470
rect 14480 34468 14528 34470
rect 14584 34468 14632 34524
rect 14688 34522 14736 34524
rect 14792 34522 14840 34524
rect 14896 34522 14944 34524
rect 14696 34470 14736 34522
rect 14820 34470 14840 34522
rect 14688 34468 14736 34470
rect 14792 34468 14840 34470
rect 14896 34468 14944 34470
rect 15000 34522 15048 34524
rect 15104 34522 15152 34524
rect 15000 34470 15016 34522
rect 15104 34470 15140 34522
rect 15000 34468 15048 34470
rect 15104 34468 15152 34470
rect 14008 34458 15208 34468
rect 24008 33740 25208 33750
rect 24064 33738 24112 33740
rect 24168 33738 24216 33740
rect 24076 33686 24112 33738
rect 24200 33686 24216 33738
rect 24064 33684 24112 33686
rect 24168 33684 24216 33686
rect 24272 33738 24320 33740
rect 24376 33738 24424 33740
rect 24480 33738 24528 33740
rect 24376 33686 24396 33738
rect 24480 33686 24520 33738
rect 24272 33684 24320 33686
rect 24376 33684 24424 33686
rect 24480 33684 24528 33686
rect 24584 33684 24632 33740
rect 24688 33738 24736 33740
rect 24792 33738 24840 33740
rect 24896 33738 24944 33740
rect 24696 33686 24736 33738
rect 24820 33686 24840 33738
rect 24688 33684 24736 33686
rect 24792 33684 24840 33686
rect 24896 33684 24944 33686
rect 25000 33738 25048 33740
rect 25104 33738 25152 33740
rect 25000 33686 25016 33738
rect 25104 33686 25140 33738
rect 25000 33684 25048 33686
rect 25104 33684 25152 33686
rect 24008 33674 25208 33684
rect 14008 32956 15208 32966
rect 14064 32954 14112 32956
rect 14168 32954 14216 32956
rect 14076 32902 14112 32954
rect 14200 32902 14216 32954
rect 14064 32900 14112 32902
rect 14168 32900 14216 32902
rect 14272 32954 14320 32956
rect 14376 32954 14424 32956
rect 14480 32954 14528 32956
rect 14376 32902 14396 32954
rect 14480 32902 14520 32954
rect 14272 32900 14320 32902
rect 14376 32900 14424 32902
rect 14480 32900 14528 32902
rect 14584 32900 14632 32956
rect 14688 32954 14736 32956
rect 14792 32954 14840 32956
rect 14896 32954 14944 32956
rect 14696 32902 14736 32954
rect 14820 32902 14840 32954
rect 14688 32900 14736 32902
rect 14792 32900 14840 32902
rect 14896 32900 14944 32902
rect 15000 32954 15048 32956
rect 15104 32954 15152 32956
rect 15000 32902 15016 32954
rect 15104 32902 15140 32954
rect 15000 32900 15048 32902
rect 15104 32900 15152 32902
rect 14008 32890 15208 32900
rect 24008 32172 25208 32182
rect 24064 32170 24112 32172
rect 24168 32170 24216 32172
rect 24076 32118 24112 32170
rect 24200 32118 24216 32170
rect 24064 32116 24112 32118
rect 24168 32116 24216 32118
rect 24272 32170 24320 32172
rect 24376 32170 24424 32172
rect 24480 32170 24528 32172
rect 24376 32118 24396 32170
rect 24480 32118 24520 32170
rect 24272 32116 24320 32118
rect 24376 32116 24424 32118
rect 24480 32116 24528 32118
rect 24584 32116 24632 32172
rect 24688 32170 24736 32172
rect 24792 32170 24840 32172
rect 24896 32170 24944 32172
rect 24696 32118 24736 32170
rect 24820 32118 24840 32170
rect 24688 32116 24736 32118
rect 24792 32116 24840 32118
rect 24896 32116 24944 32118
rect 25000 32170 25048 32172
rect 25104 32170 25152 32172
rect 25000 32118 25016 32170
rect 25104 32118 25140 32170
rect 25000 32116 25048 32118
rect 25104 32116 25152 32118
rect 24008 32106 25208 32116
rect 14008 31388 15208 31398
rect 14064 31386 14112 31388
rect 14168 31386 14216 31388
rect 14076 31334 14112 31386
rect 14200 31334 14216 31386
rect 14064 31332 14112 31334
rect 14168 31332 14216 31334
rect 14272 31386 14320 31388
rect 14376 31386 14424 31388
rect 14480 31386 14528 31388
rect 14376 31334 14396 31386
rect 14480 31334 14520 31386
rect 14272 31332 14320 31334
rect 14376 31332 14424 31334
rect 14480 31332 14528 31334
rect 14584 31332 14632 31388
rect 14688 31386 14736 31388
rect 14792 31386 14840 31388
rect 14896 31386 14944 31388
rect 14696 31334 14736 31386
rect 14820 31334 14840 31386
rect 14688 31332 14736 31334
rect 14792 31332 14840 31334
rect 14896 31332 14944 31334
rect 15000 31386 15048 31388
rect 15104 31386 15152 31388
rect 15000 31334 15016 31386
rect 15104 31334 15140 31386
rect 15000 31332 15048 31334
rect 15104 31332 15152 31334
rect 14008 31322 15208 31332
rect 24008 30604 25208 30614
rect 24064 30602 24112 30604
rect 24168 30602 24216 30604
rect 24076 30550 24112 30602
rect 24200 30550 24216 30602
rect 24064 30548 24112 30550
rect 24168 30548 24216 30550
rect 24272 30602 24320 30604
rect 24376 30602 24424 30604
rect 24480 30602 24528 30604
rect 24376 30550 24396 30602
rect 24480 30550 24520 30602
rect 24272 30548 24320 30550
rect 24376 30548 24424 30550
rect 24480 30548 24528 30550
rect 24584 30548 24632 30604
rect 24688 30602 24736 30604
rect 24792 30602 24840 30604
rect 24896 30602 24944 30604
rect 24696 30550 24736 30602
rect 24820 30550 24840 30602
rect 24688 30548 24736 30550
rect 24792 30548 24840 30550
rect 24896 30548 24944 30550
rect 25000 30602 25048 30604
rect 25104 30602 25152 30604
rect 25000 30550 25016 30602
rect 25104 30550 25140 30602
rect 25000 30548 25048 30550
rect 25104 30548 25152 30550
rect 24008 30538 25208 30548
rect 14008 29820 15208 29830
rect 14064 29818 14112 29820
rect 14168 29818 14216 29820
rect 14076 29766 14112 29818
rect 14200 29766 14216 29818
rect 14064 29764 14112 29766
rect 14168 29764 14216 29766
rect 14272 29818 14320 29820
rect 14376 29818 14424 29820
rect 14480 29818 14528 29820
rect 14376 29766 14396 29818
rect 14480 29766 14520 29818
rect 14272 29764 14320 29766
rect 14376 29764 14424 29766
rect 14480 29764 14528 29766
rect 14584 29764 14632 29820
rect 14688 29818 14736 29820
rect 14792 29818 14840 29820
rect 14896 29818 14944 29820
rect 14696 29766 14736 29818
rect 14820 29766 14840 29818
rect 14688 29764 14736 29766
rect 14792 29764 14840 29766
rect 14896 29764 14944 29766
rect 15000 29818 15048 29820
rect 15104 29818 15152 29820
rect 15000 29766 15016 29818
rect 15104 29766 15140 29818
rect 15000 29764 15048 29766
rect 15104 29764 15152 29766
rect 14008 29754 15208 29764
rect 24008 29036 25208 29046
rect 24064 29034 24112 29036
rect 24168 29034 24216 29036
rect 24076 28982 24112 29034
rect 24200 28982 24216 29034
rect 24064 28980 24112 28982
rect 24168 28980 24216 28982
rect 24272 29034 24320 29036
rect 24376 29034 24424 29036
rect 24480 29034 24528 29036
rect 24376 28982 24396 29034
rect 24480 28982 24520 29034
rect 24272 28980 24320 28982
rect 24376 28980 24424 28982
rect 24480 28980 24528 28982
rect 24584 28980 24632 29036
rect 24688 29034 24736 29036
rect 24792 29034 24840 29036
rect 24896 29034 24944 29036
rect 24696 28982 24736 29034
rect 24820 28982 24840 29034
rect 24688 28980 24736 28982
rect 24792 28980 24840 28982
rect 24896 28980 24944 28982
rect 25000 29034 25048 29036
rect 25104 29034 25152 29036
rect 25000 28982 25016 29034
rect 25104 28982 25140 29034
rect 25000 28980 25048 28982
rect 25104 28980 25152 28982
rect 24008 28970 25208 28980
rect 14008 28252 15208 28262
rect 14064 28250 14112 28252
rect 14168 28250 14216 28252
rect 14076 28198 14112 28250
rect 14200 28198 14216 28250
rect 14064 28196 14112 28198
rect 14168 28196 14216 28198
rect 14272 28250 14320 28252
rect 14376 28250 14424 28252
rect 14480 28250 14528 28252
rect 14376 28198 14396 28250
rect 14480 28198 14520 28250
rect 14272 28196 14320 28198
rect 14376 28196 14424 28198
rect 14480 28196 14528 28198
rect 14584 28196 14632 28252
rect 14688 28250 14736 28252
rect 14792 28250 14840 28252
rect 14896 28250 14944 28252
rect 14696 28198 14736 28250
rect 14820 28198 14840 28250
rect 14688 28196 14736 28198
rect 14792 28196 14840 28198
rect 14896 28196 14944 28198
rect 15000 28250 15048 28252
rect 15104 28250 15152 28252
rect 15000 28198 15016 28250
rect 15104 28198 15140 28250
rect 15000 28196 15048 28198
rect 15104 28196 15152 28198
rect 14008 28186 15208 28196
rect 24008 27468 25208 27478
rect 24064 27466 24112 27468
rect 24168 27466 24216 27468
rect 24076 27414 24112 27466
rect 24200 27414 24216 27466
rect 24064 27412 24112 27414
rect 24168 27412 24216 27414
rect 24272 27466 24320 27468
rect 24376 27466 24424 27468
rect 24480 27466 24528 27468
rect 24376 27414 24396 27466
rect 24480 27414 24520 27466
rect 24272 27412 24320 27414
rect 24376 27412 24424 27414
rect 24480 27412 24528 27414
rect 24584 27412 24632 27468
rect 24688 27466 24736 27468
rect 24792 27466 24840 27468
rect 24896 27466 24944 27468
rect 24696 27414 24736 27466
rect 24820 27414 24840 27466
rect 24688 27412 24736 27414
rect 24792 27412 24840 27414
rect 24896 27412 24944 27414
rect 25000 27466 25048 27468
rect 25104 27466 25152 27468
rect 25000 27414 25016 27466
rect 25104 27414 25140 27466
rect 25000 27412 25048 27414
rect 25104 27412 25152 27414
rect 24008 27402 25208 27412
rect 14008 26684 15208 26694
rect 14064 26682 14112 26684
rect 14168 26682 14216 26684
rect 14076 26630 14112 26682
rect 14200 26630 14216 26682
rect 14064 26628 14112 26630
rect 14168 26628 14216 26630
rect 14272 26682 14320 26684
rect 14376 26682 14424 26684
rect 14480 26682 14528 26684
rect 14376 26630 14396 26682
rect 14480 26630 14520 26682
rect 14272 26628 14320 26630
rect 14376 26628 14424 26630
rect 14480 26628 14528 26630
rect 14584 26628 14632 26684
rect 14688 26682 14736 26684
rect 14792 26682 14840 26684
rect 14896 26682 14944 26684
rect 14696 26630 14736 26682
rect 14820 26630 14840 26682
rect 14688 26628 14736 26630
rect 14792 26628 14840 26630
rect 14896 26628 14944 26630
rect 15000 26682 15048 26684
rect 15104 26682 15152 26684
rect 15000 26630 15016 26682
rect 15104 26630 15140 26682
rect 15000 26628 15048 26630
rect 15104 26628 15152 26630
rect 14008 26618 15208 26628
rect 24008 25900 25208 25910
rect 24064 25898 24112 25900
rect 24168 25898 24216 25900
rect 24076 25846 24112 25898
rect 24200 25846 24216 25898
rect 24064 25844 24112 25846
rect 24168 25844 24216 25846
rect 24272 25898 24320 25900
rect 24376 25898 24424 25900
rect 24480 25898 24528 25900
rect 24376 25846 24396 25898
rect 24480 25846 24520 25898
rect 24272 25844 24320 25846
rect 24376 25844 24424 25846
rect 24480 25844 24528 25846
rect 24584 25844 24632 25900
rect 24688 25898 24736 25900
rect 24792 25898 24840 25900
rect 24896 25898 24944 25900
rect 24696 25846 24736 25898
rect 24820 25846 24840 25898
rect 24688 25844 24736 25846
rect 24792 25844 24840 25846
rect 24896 25844 24944 25846
rect 25000 25898 25048 25900
rect 25104 25898 25152 25900
rect 25000 25846 25016 25898
rect 25104 25846 25140 25898
rect 25000 25844 25048 25846
rect 25104 25844 25152 25846
rect 24008 25834 25208 25844
rect 14008 25116 15208 25126
rect 14064 25114 14112 25116
rect 14168 25114 14216 25116
rect 14076 25062 14112 25114
rect 14200 25062 14216 25114
rect 14064 25060 14112 25062
rect 14168 25060 14216 25062
rect 14272 25114 14320 25116
rect 14376 25114 14424 25116
rect 14480 25114 14528 25116
rect 14376 25062 14396 25114
rect 14480 25062 14520 25114
rect 14272 25060 14320 25062
rect 14376 25060 14424 25062
rect 14480 25060 14528 25062
rect 14584 25060 14632 25116
rect 14688 25114 14736 25116
rect 14792 25114 14840 25116
rect 14896 25114 14944 25116
rect 14696 25062 14736 25114
rect 14820 25062 14840 25114
rect 14688 25060 14736 25062
rect 14792 25060 14840 25062
rect 14896 25060 14944 25062
rect 15000 25114 15048 25116
rect 15104 25114 15152 25116
rect 15000 25062 15016 25114
rect 15104 25062 15140 25114
rect 15000 25060 15048 25062
rect 15104 25060 15152 25062
rect 14008 25050 15208 25060
rect 24008 24332 25208 24342
rect 24064 24330 24112 24332
rect 24168 24330 24216 24332
rect 24076 24278 24112 24330
rect 24200 24278 24216 24330
rect 24064 24276 24112 24278
rect 24168 24276 24216 24278
rect 24272 24330 24320 24332
rect 24376 24330 24424 24332
rect 24480 24330 24528 24332
rect 24376 24278 24396 24330
rect 24480 24278 24520 24330
rect 24272 24276 24320 24278
rect 24376 24276 24424 24278
rect 24480 24276 24528 24278
rect 24584 24276 24632 24332
rect 24688 24330 24736 24332
rect 24792 24330 24840 24332
rect 24896 24330 24944 24332
rect 24696 24278 24736 24330
rect 24820 24278 24840 24330
rect 24688 24276 24736 24278
rect 24792 24276 24840 24278
rect 24896 24276 24944 24278
rect 25000 24330 25048 24332
rect 25104 24330 25152 24332
rect 25000 24278 25016 24330
rect 25104 24278 25140 24330
rect 25000 24276 25048 24278
rect 25104 24276 25152 24278
rect 24008 24266 25208 24276
rect 14008 23548 15208 23558
rect 14064 23546 14112 23548
rect 14168 23546 14216 23548
rect 14076 23494 14112 23546
rect 14200 23494 14216 23546
rect 14064 23492 14112 23494
rect 14168 23492 14216 23494
rect 14272 23546 14320 23548
rect 14376 23546 14424 23548
rect 14480 23546 14528 23548
rect 14376 23494 14396 23546
rect 14480 23494 14520 23546
rect 14272 23492 14320 23494
rect 14376 23492 14424 23494
rect 14480 23492 14528 23494
rect 14584 23492 14632 23548
rect 14688 23546 14736 23548
rect 14792 23546 14840 23548
rect 14896 23546 14944 23548
rect 14696 23494 14736 23546
rect 14820 23494 14840 23546
rect 14688 23492 14736 23494
rect 14792 23492 14840 23494
rect 14896 23492 14944 23494
rect 15000 23546 15048 23548
rect 15104 23546 15152 23548
rect 15000 23494 15016 23546
rect 15104 23494 15140 23546
rect 15000 23492 15048 23494
rect 15104 23492 15152 23494
rect 14008 23482 15208 23492
rect 24008 22764 25208 22774
rect 24064 22762 24112 22764
rect 24168 22762 24216 22764
rect 24076 22710 24112 22762
rect 24200 22710 24216 22762
rect 24064 22708 24112 22710
rect 24168 22708 24216 22710
rect 24272 22762 24320 22764
rect 24376 22762 24424 22764
rect 24480 22762 24528 22764
rect 24376 22710 24396 22762
rect 24480 22710 24520 22762
rect 24272 22708 24320 22710
rect 24376 22708 24424 22710
rect 24480 22708 24528 22710
rect 24584 22708 24632 22764
rect 24688 22762 24736 22764
rect 24792 22762 24840 22764
rect 24896 22762 24944 22764
rect 24696 22710 24736 22762
rect 24820 22710 24840 22762
rect 24688 22708 24736 22710
rect 24792 22708 24840 22710
rect 24896 22708 24944 22710
rect 25000 22762 25048 22764
rect 25104 22762 25152 22764
rect 25000 22710 25016 22762
rect 25104 22710 25140 22762
rect 25000 22708 25048 22710
rect 25104 22708 25152 22710
rect 24008 22698 25208 22708
rect 14008 21980 15208 21990
rect 14064 21978 14112 21980
rect 14168 21978 14216 21980
rect 14076 21926 14112 21978
rect 14200 21926 14216 21978
rect 14064 21924 14112 21926
rect 14168 21924 14216 21926
rect 14272 21978 14320 21980
rect 14376 21978 14424 21980
rect 14480 21978 14528 21980
rect 14376 21926 14396 21978
rect 14480 21926 14520 21978
rect 14272 21924 14320 21926
rect 14376 21924 14424 21926
rect 14480 21924 14528 21926
rect 14584 21924 14632 21980
rect 14688 21978 14736 21980
rect 14792 21978 14840 21980
rect 14896 21978 14944 21980
rect 14696 21926 14736 21978
rect 14820 21926 14840 21978
rect 14688 21924 14736 21926
rect 14792 21924 14840 21926
rect 14896 21924 14944 21926
rect 15000 21978 15048 21980
rect 15104 21978 15152 21980
rect 15000 21926 15016 21978
rect 15104 21926 15140 21978
rect 15000 21924 15048 21926
rect 15104 21924 15152 21926
rect 14008 21914 15208 21924
rect 24008 21196 25208 21206
rect 24064 21194 24112 21196
rect 24168 21194 24216 21196
rect 24076 21142 24112 21194
rect 24200 21142 24216 21194
rect 24064 21140 24112 21142
rect 24168 21140 24216 21142
rect 24272 21194 24320 21196
rect 24376 21194 24424 21196
rect 24480 21194 24528 21196
rect 24376 21142 24396 21194
rect 24480 21142 24520 21194
rect 24272 21140 24320 21142
rect 24376 21140 24424 21142
rect 24480 21140 24528 21142
rect 24584 21140 24632 21196
rect 24688 21194 24736 21196
rect 24792 21194 24840 21196
rect 24896 21194 24944 21196
rect 24696 21142 24736 21194
rect 24820 21142 24840 21194
rect 24688 21140 24736 21142
rect 24792 21140 24840 21142
rect 24896 21140 24944 21142
rect 25000 21194 25048 21196
rect 25104 21194 25152 21196
rect 25000 21142 25016 21194
rect 25104 21142 25140 21194
rect 25000 21140 25048 21142
rect 25104 21140 25152 21142
rect 24008 21130 25208 21140
rect 14008 20412 15208 20422
rect 14064 20410 14112 20412
rect 14168 20410 14216 20412
rect 14076 20358 14112 20410
rect 14200 20358 14216 20410
rect 14064 20356 14112 20358
rect 14168 20356 14216 20358
rect 14272 20410 14320 20412
rect 14376 20410 14424 20412
rect 14480 20410 14528 20412
rect 14376 20358 14396 20410
rect 14480 20358 14520 20410
rect 14272 20356 14320 20358
rect 14376 20356 14424 20358
rect 14480 20356 14528 20358
rect 14584 20356 14632 20412
rect 14688 20410 14736 20412
rect 14792 20410 14840 20412
rect 14896 20410 14944 20412
rect 14696 20358 14736 20410
rect 14820 20358 14840 20410
rect 14688 20356 14736 20358
rect 14792 20356 14840 20358
rect 14896 20356 14944 20358
rect 15000 20410 15048 20412
rect 15104 20410 15152 20412
rect 15000 20358 15016 20410
rect 15104 20358 15140 20410
rect 15000 20356 15048 20358
rect 15104 20356 15152 20358
rect 14008 20346 15208 20356
rect 24008 19628 25208 19638
rect 24064 19626 24112 19628
rect 24168 19626 24216 19628
rect 24076 19574 24112 19626
rect 24200 19574 24216 19626
rect 24064 19572 24112 19574
rect 24168 19572 24216 19574
rect 24272 19626 24320 19628
rect 24376 19626 24424 19628
rect 24480 19626 24528 19628
rect 24376 19574 24396 19626
rect 24480 19574 24520 19626
rect 24272 19572 24320 19574
rect 24376 19572 24424 19574
rect 24480 19572 24528 19574
rect 24584 19572 24632 19628
rect 24688 19626 24736 19628
rect 24792 19626 24840 19628
rect 24896 19626 24944 19628
rect 24696 19574 24736 19626
rect 24820 19574 24840 19626
rect 24688 19572 24736 19574
rect 24792 19572 24840 19574
rect 24896 19572 24944 19574
rect 25000 19626 25048 19628
rect 25104 19626 25152 19628
rect 25000 19574 25016 19626
rect 25104 19574 25140 19626
rect 25000 19572 25048 19574
rect 25104 19572 25152 19574
rect 24008 19562 25208 19572
rect 14008 18844 15208 18854
rect 14064 18842 14112 18844
rect 14168 18842 14216 18844
rect 14076 18790 14112 18842
rect 14200 18790 14216 18842
rect 14064 18788 14112 18790
rect 14168 18788 14216 18790
rect 14272 18842 14320 18844
rect 14376 18842 14424 18844
rect 14480 18842 14528 18844
rect 14376 18790 14396 18842
rect 14480 18790 14520 18842
rect 14272 18788 14320 18790
rect 14376 18788 14424 18790
rect 14480 18788 14528 18790
rect 14584 18788 14632 18844
rect 14688 18842 14736 18844
rect 14792 18842 14840 18844
rect 14896 18842 14944 18844
rect 14696 18790 14736 18842
rect 14820 18790 14840 18842
rect 14688 18788 14736 18790
rect 14792 18788 14840 18790
rect 14896 18788 14944 18790
rect 15000 18842 15048 18844
rect 15104 18842 15152 18844
rect 15000 18790 15016 18842
rect 15104 18790 15140 18842
rect 15000 18788 15048 18790
rect 15104 18788 15152 18790
rect 14008 18778 15208 18788
rect 24008 18060 25208 18070
rect 24064 18058 24112 18060
rect 24168 18058 24216 18060
rect 24076 18006 24112 18058
rect 24200 18006 24216 18058
rect 24064 18004 24112 18006
rect 24168 18004 24216 18006
rect 24272 18058 24320 18060
rect 24376 18058 24424 18060
rect 24480 18058 24528 18060
rect 24376 18006 24396 18058
rect 24480 18006 24520 18058
rect 24272 18004 24320 18006
rect 24376 18004 24424 18006
rect 24480 18004 24528 18006
rect 24584 18004 24632 18060
rect 24688 18058 24736 18060
rect 24792 18058 24840 18060
rect 24896 18058 24944 18060
rect 24696 18006 24736 18058
rect 24820 18006 24840 18058
rect 24688 18004 24736 18006
rect 24792 18004 24840 18006
rect 24896 18004 24944 18006
rect 25000 18058 25048 18060
rect 25104 18058 25152 18060
rect 25000 18006 25016 18058
rect 25104 18006 25140 18058
rect 25000 18004 25048 18006
rect 25104 18004 25152 18006
rect 24008 17994 25208 18004
rect 14008 17276 15208 17286
rect 14064 17274 14112 17276
rect 14168 17274 14216 17276
rect 14076 17222 14112 17274
rect 14200 17222 14216 17274
rect 14064 17220 14112 17222
rect 14168 17220 14216 17222
rect 14272 17274 14320 17276
rect 14376 17274 14424 17276
rect 14480 17274 14528 17276
rect 14376 17222 14396 17274
rect 14480 17222 14520 17274
rect 14272 17220 14320 17222
rect 14376 17220 14424 17222
rect 14480 17220 14528 17222
rect 14584 17220 14632 17276
rect 14688 17274 14736 17276
rect 14792 17274 14840 17276
rect 14896 17274 14944 17276
rect 14696 17222 14736 17274
rect 14820 17222 14840 17274
rect 14688 17220 14736 17222
rect 14792 17220 14840 17222
rect 14896 17220 14944 17222
rect 15000 17274 15048 17276
rect 15104 17274 15152 17276
rect 15000 17222 15016 17274
rect 15104 17222 15140 17274
rect 15000 17220 15048 17222
rect 15104 17220 15152 17222
rect 14008 17210 15208 17220
rect 24008 16492 25208 16502
rect 24064 16490 24112 16492
rect 24168 16490 24216 16492
rect 24076 16438 24112 16490
rect 24200 16438 24216 16490
rect 24064 16436 24112 16438
rect 24168 16436 24216 16438
rect 24272 16490 24320 16492
rect 24376 16490 24424 16492
rect 24480 16490 24528 16492
rect 24376 16438 24396 16490
rect 24480 16438 24520 16490
rect 24272 16436 24320 16438
rect 24376 16436 24424 16438
rect 24480 16436 24528 16438
rect 24584 16436 24632 16492
rect 24688 16490 24736 16492
rect 24792 16490 24840 16492
rect 24896 16490 24944 16492
rect 24696 16438 24736 16490
rect 24820 16438 24840 16490
rect 24688 16436 24736 16438
rect 24792 16436 24840 16438
rect 24896 16436 24944 16438
rect 25000 16490 25048 16492
rect 25104 16490 25152 16492
rect 25000 16438 25016 16490
rect 25104 16438 25140 16490
rect 25000 16436 25048 16438
rect 25104 16436 25152 16438
rect 24008 16426 25208 16436
rect 14008 15708 15208 15718
rect 14064 15706 14112 15708
rect 14168 15706 14216 15708
rect 14076 15654 14112 15706
rect 14200 15654 14216 15706
rect 14064 15652 14112 15654
rect 14168 15652 14216 15654
rect 14272 15706 14320 15708
rect 14376 15706 14424 15708
rect 14480 15706 14528 15708
rect 14376 15654 14396 15706
rect 14480 15654 14520 15706
rect 14272 15652 14320 15654
rect 14376 15652 14424 15654
rect 14480 15652 14528 15654
rect 14584 15652 14632 15708
rect 14688 15706 14736 15708
rect 14792 15706 14840 15708
rect 14896 15706 14944 15708
rect 14696 15654 14736 15706
rect 14820 15654 14840 15706
rect 14688 15652 14736 15654
rect 14792 15652 14840 15654
rect 14896 15652 14944 15654
rect 15000 15706 15048 15708
rect 15104 15706 15152 15708
rect 15000 15654 15016 15706
rect 15104 15654 15140 15706
rect 15000 15652 15048 15654
rect 15104 15652 15152 15654
rect 14008 15642 15208 15652
rect 24008 14924 25208 14934
rect 24064 14922 24112 14924
rect 24168 14922 24216 14924
rect 24076 14870 24112 14922
rect 24200 14870 24216 14922
rect 24064 14868 24112 14870
rect 24168 14868 24216 14870
rect 24272 14922 24320 14924
rect 24376 14922 24424 14924
rect 24480 14922 24528 14924
rect 24376 14870 24396 14922
rect 24480 14870 24520 14922
rect 24272 14868 24320 14870
rect 24376 14868 24424 14870
rect 24480 14868 24528 14870
rect 24584 14868 24632 14924
rect 24688 14922 24736 14924
rect 24792 14922 24840 14924
rect 24896 14922 24944 14924
rect 24696 14870 24736 14922
rect 24820 14870 24840 14922
rect 24688 14868 24736 14870
rect 24792 14868 24840 14870
rect 24896 14868 24944 14870
rect 25000 14922 25048 14924
rect 25104 14922 25152 14924
rect 25000 14870 25016 14922
rect 25104 14870 25140 14922
rect 25000 14868 25048 14870
rect 25104 14868 25152 14870
rect 24008 14858 25208 14868
rect 14008 14140 15208 14150
rect 14064 14138 14112 14140
rect 14168 14138 14216 14140
rect 14076 14086 14112 14138
rect 14200 14086 14216 14138
rect 14064 14084 14112 14086
rect 14168 14084 14216 14086
rect 14272 14138 14320 14140
rect 14376 14138 14424 14140
rect 14480 14138 14528 14140
rect 14376 14086 14396 14138
rect 14480 14086 14520 14138
rect 14272 14084 14320 14086
rect 14376 14084 14424 14086
rect 14480 14084 14528 14086
rect 14584 14084 14632 14140
rect 14688 14138 14736 14140
rect 14792 14138 14840 14140
rect 14896 14138 14944 14140
rect 14696 14086 14736 14138
rect 14820 14086 14840 14138
rect 14688 14084 14736 14086
rect 14792 14084 14840 14086
rect 14896 14084 14944 14086
rect 15000 14138 15048 14140
rect 15104 14138 15152 14140
rect 15000 14086 15016 14138
rect 15104 14086 15140 14138
rect 15000 14084 15048 14086
rect 15104 14084 15152 14086
rect 14008 14074 15208 14084
rect 24008 13356 25208 13366
rect 24064 13354 24112 13356
rect 24168 13354 24216 13356
rect 24076 13302 24112 13354
rect 24200 13302 24216 13354
rect 24064 13300 24112 13302
rect 24168 13300 24216 13302
rect 24272 13354 24320 13356
rect 24376 13354 24424 13356
rect 24480 13354 24528 13356
rect 24376 13302 24396 13354
rect 24480 13302 24520 13354
rect 24272 13300 24320 13302
rect 24376 13300 24424 13302
rect 24480 13300 24528 13302
rect 24584 13300 24632 13356
rect 24688 13354 24736 13356
rect 24792 13354 24840 13356
rect 24896 13354 24944 13356
rect 24696 13302 24736 13354
rect 24820 13302 24840 13354
rect 24688 13300 24736 13302
rect 24792 13300 24840 13302
rect 24896 13300 24944 13302
rect 25000 13354 25048 13356
rect 25104 13354 25152 13356
rect 25000 13302 25016 13354
rect 25104 13302 25140 13354
rect 25000 13300 25048 13302
rect 25104 13300 25152 13302
rect 24008 13290 25208 13300
rect 14008 12572 15208 12582
rect 14064 12570 14112 12572
rect 14168 12570 14216 12572
rect 14076 12518 14112 12570
rect 14200 12518 14216 12570
rect 14064 12516 14112 12518
rect 14168 12516 14216 12518
rect 14272 12570 14320 12572
rect 14376 12570 14424 12572
rect 14480 12570 14528 12572
rect 14376 12518 14396 12570
rect 14480 12518 14520 12570
rect 14272 12516 14320 12518
rect 14376 12516 14424 12518
rect 14480 12516 14528 12518
rect 14584 12516 14632 12572
rect 14688 12570 14736 12572
rect 14792 12570 14840 12572
rect 14896 12570 14944 12572
rect 14696 12518 14736 12570
rect 14820 12518 14840 12570
rect 14688 12516 14736 12518
rect 14792 12516 14840 12518
rect 14896 12516 14944 12518
rect 15000 12570 15048 12572
rect 15104 12570 15152 12572
rect 15000 12518 15016 12570
rect 15104 12518 15140 12570
rect 15000 12516 15048 12518
rect 15104 12516 15152 12518
rect 14008 12506 15208 12516
rect 24008 11788 25208 11798
rect 24064 11786 24112 11788
rect 24168 11786 24216 11788
rect 24076 11734 24112 11786
rect 24200 11734 24216 11786
rect 24064 11732 24112 11734
rect 24168 11732 24216 11734
rect 24272 11786 24320 11788
rect 24376 11786 24424 11788
rect 24480 11786 24528 11788
rect 24376 11734 24396 11786
rect 24480 11734 24520 11786
rect 24272 11732 24320 11734
rect 24376 11732 24424 11734
rect 24480 11732 24528 11734
rect 24584 11732 24632 11788
rect 24688 11786 24736 11788
rect 24792 11786 24840 11788
rect 24896 11786 24944 11788
rect 24696 11734 24736 11786
rect 24820 11734 24840 11786
rect 24688 11732 24736 11734
rect 24792 11732 24840 11734
rect 24896 11732 24944 11734
rect 25000 11786 25048 11788
rect 25104 11786 25152 11788
rect 25000 11734 25016 11786
rect 25104 11734 25140 11786
rect 25000 11732 25048 11734
rect 25104 11732 25152 11734
rect 24008 11722 25208 11732
rect 14008 11004 15208 11014
rect 14064 11002 14112 11004
rect 14168 11002 14216 11004
rect 14076 10950 14112 11002
rect 14200 10950 14216 11002
rect 14064 10948 14112 10950
rect 14168 10948 14216 10950
rect 14272 11002 14320 11004
rect 14376 11002 14424 11004
rect 14480 11002 14528 11004
rect 14376 10950 14396 11002
rect 14480 10950 14520 11002
rect 14272 10948 14320 10950
rect 14376 10948 14424 10950
rect 14480 10948 14528 10950
rect 14584 10948 14632 11004
rect 14688 11002 14736 11004
rect 14792 11002 14840 11004
rect 14896 11002 14944 11004
rect 14696 10950 14736 11002
rect 14820 10950 14840 11002
rect 14688 10948 14736 10950
rect 14792 10948 14840 10950
rect 14896 10948 14944 10950
rect 15000 11002 15048 11004
rect 15104 11002 15152 11004
rect 15000 10950 15016 11002
rect 15104 10950 15140 11002
rect 15000 10948 15048 10950
rect 15104 10948 15152 10950
rect 14008 10938 15208 10948
rect 24008 10220 25208 10230
rect 24064 10218 24112 10220
rect 24168 10218 24216 10220
rect 24076 10166 24112 10218
rect 24200 10166 24216 10218
rect 24064 10164 24112 10166
rect 24168 10164 24216 10166
rect 24272 10218 24320 10220
rect 24376 10218 24424 10220
rect 24480 10218 24528 10220
rect 24376 10166 24396 10218
rect 24480 10166 24520 10218
rect 24272 10164 24320 10166
rect 24376 10164 24424 10166
rect 24480 10164 24528 10166
rect 24584 10164 24632 10220
rect 24688 10218 24736 10220
rect 24792 10218 24840 10220
rect 24896 10218 24944 10220
rect 24696 10166 24736 10218
rect 24820 10166 24840 10218
rect 24688 10164 24736 10166
rect 24792 10164 24840 10166
rect 24896 10164 24944 10166
rect 25000 10218 25048 10220
rect 25104 10218 25152 10220
rect 25000 10166 25016 10218
rect 25104 10166 25140 10218
rect 25000 10164 25048 10166
rect 25104 10164 25152 10166
rect 24008 10154 25208 10164
rect 14008 9436 15208 9446
rect 14064 9434 14112 9436
rect 14168 9434 14216 9436
rect 14076 9382 14112 9434
rect 14200 9382 14216 9434
rect 14064 9380 14112 9382
rect 14168 9380 14216 9382
rect 14272 9434 14320 9436
rect 14376 9434 14424 9436
rect 14480 9434 14528 9436
rect 14376 9382 14396 9434
rect 14480 9382 14520 9434
rect 14272 9380 14320 9382
rect 14376 9380 14424 9382
rect 14480 9380 14528 9382
rect 14584 9380 14632 9436
rect 14688 9434 14736 9436
rect 14792 9434 14840 9436
rect 14896 9434 14944 9436
rect 14696 9382 14736 9434
rect 14820 9382 14840 9434
rect 14688 9380 14736 9382
rect 14792 9380 14840 9382
rect 14896 9380 14944 9382
rect 15000 9434 15048 9436
rect 15104 9434 15152 9436
rect 15000 9382 15016 9434
rect 15104 9382 15140 9434
rect 15000 9380 15048 9382
rect 15104 9380 15152 9382
rect 14008 9370 15208 9380
rect 24008 8652 25208 8662
rect 24064 8650 24112 8652
rect 24168 8650 24216 8652
rect 24076 8598 24112 8650
rect 24200 8598 24216 8650
rect 24064 8596 24112 8598
rect 24168 8596 24216 8598
rect 24272 8650 24320 8652
rect 24376 8650 24424 8652
rect 24480 8650 24528 8652
rect 24376 8598 24396 8650
rect 24480 8598 24520 8650
rect 24272 8596 24320 8598
rect 24376 8596 24424 8598
rect 24480 8596 24528 8598
rect 24584 8596 24632 8652
rect 24688 8650 24736 8652
rect 24792 8650 24840 8652
rect 24896 8650 24944 8652
rect 24696 8598 24736 8650
rect 24820 8598 24840 8650
rect 24688 8596 24736 8598
rect 24792 8596 24840 8598
rect 24896 8596 24944 8598
rect 25000 8650 25048 8652
rect 25104 8650 25152 8652
rect 25000 8598 25016 8650
rect 25104 8598 25140 8650
rect 25000 8596 25048 8598
rect 25104 8596 25152 8598
rect 24008 8586 25208 8596
rect 14252 8148 14308 8158
rect 14252 8054 14308 8092
rect 16492 8036 16548 8046
rect 16492 7942 16548 7980
rect 28364 8036 28420 45612
rect 37212 45668 37268 45678
rect 37436 45668 37492 45678
rect 37212 45666 37492 45668
rect 37212 45614 37214 45666
rect 37266 45614 37438 45666
rect 37490 45614 37492 45666
rect 37212 45612 37492 45614
rect 37212 45602 37268 45612
rect 34008 45500 35208 45510
rect 34064 45498 34112 45500
rect 34168 45498 34216 45500
rect 34076 45446 34112 45498
rect 34200 45446 34216 45498
rect 34064 45444 34112 45446
rect 34168 45444 34216 45446
rect 34272 45498 34320 45500
rect 34376 45498 34424 45500
rect 34480 45498 34528 45500
rect 34376 45446 34396 45498
rect 34480 45446 34520 45498
rect 34272 45444 34320 45446
rect 34376 45444 34424 45446
rect 34480 45444 34528 45446
rect 34584 45444 34632 45500
rect 34688 45498 34736 45500
rect 34792 45498 34840 45500
rect 34896 45498 34944 45500
rect 34696 45446 34736 45498
rect 34820 45446 34840 45498
rect 34688 45444 34736 45446
rect 34792 45444 34840 45446
rect 34896 45444 34944 45446
rect 35000 45498 35048 45500
rect 35104 45498 35152 45500
rect 35000 45446 35016 45498
rect 35104 45446 35140 45498
rect 35000 45444 35048 45446
rect 35104 45444 35152 45446
rect 34008 45434 35208 45444
rect 34008 43932 35208 43942
rect 34064 43930 34112 43932
rect 34168 43930 34216 43932
rect 34076 43878 34112 43930
rect 34200 43878 34216 43930
rect 34064 43876 34112 43878
rect 34168 43876 34216 43878
rect 34272 43930 34320 43932
rect 34376 43930 34424 43932
rect 34480 43930 34528 43932
rect 34376 43878 34396 43930
rect 34480 43878 34520 43930
rect 34272 43876 34320 43878
rect 34376 43876 34424 43878
rect 34480 43876 34528 43878
rect 34584 43876 34632 43932
rect 34688 43930 34736 43932
rect 34792 43930 34840 43932
rect 34896 43930 34944 43932
rect 34696 43878 34736 43930
rect 34820 43878 34840 43930
rect 34688 43876 34736 43878
rect 34792 43876 34840 43878
rect 34896 43876 34944 43878
rect 35000 43930 35048 43932
rect 35104 43930 35152 43932
rect 35000 43878 35016 43930
rect 35104 43878 35140 43930
rect 35000 43876 35048 43878
rect 35104 43876 35152 43878
rect 34008 43866 35208 43876
rect 34008 42364 35208 42374
rect 34064 42362 34112 42364
rect 34168 42362 34216 42364
rect 34076 42310 34112 42362
rect 34200 42310 34216 42362
rect 34064 42308 34112 42310
rect 34168 42308 34216 42310
rect 34272 42362 34320 42364
rect 34376 42362 34424 42364
rect 34480 42362 34528 42364
rect 34376 42310 34396 42362
rect 34480 42310 34520 42362
rect 34272 42308 34320 42310
rect 34376 42308 34424 42310
rect 34480 42308 34528 42310
rect 34584 42308 34632 42364
rect 34688 42362 34736 42364
rect 34792 42362 34840 42364
rect 34896 42362 34944 42364
rect 34696 42310 34736 42362
rect 34820 42310 34840 42362
rect 34688 42308 34736 42310
rect 34792 42308 34840 42310
rect 34896 42308 34944 42310
rect 35000 42362 35048 42364
rect 35104 42362 35152 42364
rect 35000 42310 35016 42362
rect 35104 42310 35140 42362
rect 35000 42308 35048 42310
rect 35104 42308 35152 42310
rect 34008 42298 35208 42308
rect 34008 40796 35208 40806
rect 34064 40794 34112 40796
rect 34168 40794 34216 40796
rect 34076 40742 34112 40794
rect 34200 40742 34216 40794
rect 34064 40740 34112 40742
rect 34168 40740 34216 40742
rect 34272 40794 34320 40796
rect 34376 40794 34424 40796
rect 34480 40794 34528 40796
rect 34376 40742 34396 40794
rect 34480 40742 34520 40794
rect 34272 40740 34320 40742
rect 34376 40740 34424 40742
rect 34480 40740 34528 40742
rect 34584 40740 34632 40796
rect 34688 40794 34736 40796
rect 34792 40794 34840 40796
rect 34896 40794 34944 40796
rect 34696 40742 34736 40794
rect 34820 40742 34840 40794
rect 34688 40740 34736 40742
rect 34792 40740 34840 40742
rect 34896 40740 34944 40742
rect 35000 40794 35048 40796
rect 35104 40794 35152 40796
rect 35000 40742 35016 40794
rect 35104 40742 35140 40794
rect 35000 40740 35048 40742
rect 35104 40740 35152 40742
rect 34008 40730 35208 40740
rect 34008 39228 35208 39238
rect 34064 39226 34112 39228
rect 34168 39226 34216 39228
rect 34076 39174 34112 39226
rect 34200 39174 34216 39226
rect 34064 39172 34112 39174
rect 34168 39172 34216 39174
rect 34272 39226 34320 39228
rect 34376 39226 34424 39228
rect 34480 39226 34528 39228
rect 34376 39174 34396 39226
rect 34480 39174 34520 39226
rect 34272 39172 34320 39174
rect 34376 39172 34424 39174
rect 34480 39172 34528 39174
rect 34584 39172 34632 39228
rect 34688 39226 34736 39228
rect 34792 39226 34840 39228
rect 34896 39226 34944 39228
rect 34696 39174 34736 39226
rect 34820 39174 34840 39226
rect 34688 39172 34736 39174
rect 34792 39172 34840 39174
rect 34896 39172 34944 39174
rect 35000 39226 35048 39228
rect 35104 39226 35152 39228
rect 35000 39174 35016 39226
rect 35104 39174 35140 39226
rect 35000 39172 35048 39174
rect 35104 39172 35152 39174
rect 34008 39162 35208 39172
rect 34008 37660 35208 37670
rect 34064 37658 34112 37660
rect 34168 37658 34216 37660
rect 34076 37606 34112 37658
rect 34200 37606 34216 37658
rect 34064 37604 34112 37606
rect 34168 37604 34216 37606
rect 34272 37658 34320 37660
rect 34376 37658 34424 37660
rect 34480 37658 34528 37660
rect 34376 37606 34396 37658
rect 34480 37606 34520 37658
rect 34272 37604 34320 37606
rect 34376 37604 34424 37606
rect 34480 37604 34528 37606
rect 34584 37604 34632 37660
rect 34688 37658 34736 37660
rect 34792 37658 34840 37660
rect 34896 37658 34944 37660
rect 34696 37606 34736 37658
rect 34820 37606 34840 37658
rect 34688 37604 34736 37606
rect 34792 37604 34840 37606
rect 34896 37604 34944 37606
rect 35000 37658 35048 37660
rect 35104 37658 35152 37660
rect 35000 37606 35016 37658
rect 35104 37606 35140 37658
rect 35000 37604 35048 37606
rect 35104 37604 35152 37606
rect 34008 37594 35208 37604
rect 34008 36092 35208 36102
rect 34064 36090 34112 36092
rect 34168 36090 34216 36092
rect 34076 36038 34112 36090
rect 34200 36038 34216 36090
rect 34064 36036 34112 36038
rect 34168 36036 34216 36038
rect 34272 36090 34320 36092
rect 34376 36090 34424 36092
rect 34480 36090 34528 36092
rect 34376 36038 34396 36090
rect 34480 36038 34520 36090
rect 34272 36036 34320 36038
rect 34376 36036 34424 36038
rect 34480 36036 34528 36038
rect 34584 36036 34632 36092
rect 34688 36090 34736 36092
rect 34792 36090 34840 36092
rect 34896 36090 34944 36092
rect 34696 36038 34736 36090
rect 34820 36038 34840 36090
rect 34688 36036 34736 36038
rect 34792 36036 34840 36038
rect 34896 36036 34944 36038
rect 35000 36090 35048 36092
rect 35104 36090 35152 36092
rect 35000 36038 35016 36090
rect 35104 36038 35140 36090
rect 35000 36036 35048 36038
rect 35104 36036 35152 36038
rect 34008 36026 35208 36036
rect 34008 34524 35208 34534
rect 34064 34522 34112 34524
rect 34168 34522 34216 34524
rect 34076 34470 34112 34522
rect 34200 34470 34216 34522
rect 34064 34468 34112 34470
rect 34168 34468 34216 34470
rect 34272 34522 34320 34524
rect 34376 34522 34424 34524
rect 34480 34522 34528 34524
rect 34376 34470 34396 34522
rect 34480 34470 34520 34522
rect 34272 34468 34320 34470
rect 34376 34468 34424 34470
rect 34480 34468 34528 34470
rect 34584 34468 34632 34524
rect 34688 34522 34736 34524
rect 34792 34522 34840 34524
rect 34896 34522 34944 34524
rect 34696 34470 34736 34522
rect 34820 34470 34840 34522
rect 34688 34468 34736 34470
rect 34792 34468 34840 34470
rect 34896 34468 34944 34470
rect 35000 34522 35048 34524
rect 35104 34522 35152 34524
rect 35000 34470 35016 34522
rect 35104 34470 35140 34522
rect 35000 34468 35048 34470
rect 35104 34468 35152 34470
rect 34008 34458 35208 34468
rect 34008 32956 35208 32966
rect 34064 32954 34112 32956
rect 34168 32954 34216 32956
rect 34076 32902 34112 32954
rect 34200 32902 34216 32954
rect 34064 32900 34112 32902
rect 34168 32900 34216 32902
rect 34272 32954 34320 32956
rect 34376 32954 34424 32956
rect 34480 32954 34528 32956
rect 34376 32902 34396 32954
rect 34480 32902 34520 32954
rect 34272 32900 34320 32902
rect 34376 32900 34424 32902
rect 34480 32900 34528 32902
rect 34584 32900 34632 32956
rect 34688 32954 34736 32956
rect 34792 32954 34840 32956
rect 34896 32954 34944 32956
rect 34696 32902 34736 32954
rect 34820 32902 34840 32954
rect 34688 32900 34736 32902
rect 34792 32900 34840 32902
rect 34896 32900 34944 32902
rect 35000 32954 35048 32956
rect 35104 32954 35152 32956
rect 35000 32902 35016 32954
rect 35104 32902 35140 32954
rect 35000 32900 35048 32902
rect 35104 32900 35152 32902
rect 34008 32890 35208 32900
rect 34008 31388 35208 31398
rect 34064 31386 34112 31388
rect 34168 31386 34216 31388
rect 34076 31334 34112 31386
rect 34200 31334 34216 31386
rect 34064 31332 34112 31334
rect 34168 31332 34216 31334
rect 34272 31386 34320 31388
rect 34376 31386 34424 31388
rect 34480 31386 34528 31388
rect 34376 31334 34396 31386
rect 34480 31334 34520 31386
rect 34272 31332 34320 31334
rect 34376 31332 34424 31334
rect 34480 31332 34528 31334
rect 34584 31332 34632 31388
rect 34688 31386 34736 31388
rect 34792 31386 34840 31388
rect 34896 31386 34944 31388
rect 34696 31334 34736 31386
rect 34820 31334 34840 31386
rect 34688 31332 34736 31334
rect 34792 31332 34840 31334
rect 34896 31332 34944 31334
rect 35000 31386 35048 31388
rect 35104 31386 35152 31388
rect 35000 31334 35016 31386
rect 35104 31334 35140 31386
rect 35000 31332 35048 31334
rect 35104 31332 35152 31334
rect 34008 31322 35208 31332
rect 34008 29820 35208 29830
rect 34064 29818 34112 29820
rect 34168 29818 34216 29820
rect 34076 29766 34112 29818
rect 34200 29766 34216 29818
rect 34064 29764 34112 29766
rect 34168 29764 34216 29766
rect 34272 29818 34320 29820
rect 34376 29818 34424 29820
rect 34480 29818 34528 29820
rect 34376 29766 34396 29818
rect 34480 29766 34520 29818
rect 34272 29764 34320 29766
rect 34376 29764 34424 29766
rect 34480 29764 34528 29766
rect 34584 29764 34632 29820
rect 34688 29818 34736 29820
rect 34792 29818 34840 29820
rect 34896 29818 34944 29820
rect 34696 29766 34736 29818
rect 34820 29766 34840 29818
rect 34688 29764 34736 29766
rect 34792 29764 34840 29766
rect 34896 29764 34944 29766
rect 35000 29818 35048 29820
rect 35104 29818 35152 29820
rect 35000 29766 35016 29818
rect 35104 29766 35140 29818
rect 35000 29764 35048 29766
rect 35104 29764 35152 29766
rect 34008 29754 35208 29764
rect 34008 28252 35208 28262
rect 34064 28250 34112 28252
rect 34168 28250 34216 28252
rect 34076 28198 34112 28250
rect 34200 28198 34216 28250
rect 34064 28196 34112 28198
rect 34168 28196 34216 28198
rect 34272 28250 34320 28252
rect 34376 28250 34424 28252
rect 34480 28250 34528 28252
rect 34376 28198 34396 28250
rect 34480 28198 34520 28250
rect 34272 28196 34320 28198
rect 34376 28196 34424 28198
rect 34480 28196 34528 28198
rect 34584 28196 34632 28252
rect 34688 28250 34736 28252
rect 34792 28250 34840 28252
rect 34896 28250 34944 28252
rect 34696 28198 34736 28250
rect 34820 28198 34840 28250
rect 34688 28196 34736 28198
rect 34792 28196 34840 28198
rect 34896 28196 34944 28198
rect 35000 28250 35048 28252
rect 35104 28250 35152 28252
rect 35000 28198 35016 28250
rect 35104 28198 35140 28250
rect 35000 28196 35048 28198
rect 35104 28196 35152 28198
rect 34008 28186 35208 28196
rect 34008 26684 35208 26694
rect 34064 26682 34112 26684
rect 34168 26682 34216 26684
rect 34076 26630 34112 26682
rect 34200 26630 34216 26682
rect 34064 26628 34112 26630
rect 34168 26628 34216 26630
rect 34272 26682 34320 26684
rect 34376 26682 34424 26684
rect 34480 26682 34528 26684
rect 34376 26630 34396 26682
rect 34480 26630 34520 26682
rect 34272 26628 34320 26630
rect 34376 26628 34424 26630
rect 34480 26628 34528 26630
rect 34584 26628 34632 26684
rect 34688 26682 34736 26684
rect 34792 26682 34840 26684
rect 34896 26682 34944 26684
rect 34696 26630 34736 26682
rect 34820 26630 34840 26682
rect 34688 26628 34736 26630
rect 34792 26628 34840 26630
rect 34896 26628 34944 26630
rect 35000 26682 35048 26684
rect 35104 26682 35152 26684
rect 35000 26630 35016 26682
rect 35104 26630 35140 26682
rect 35000 26628 35048 26630
rect 35104 26628 35152 26630
rect 34008 26618 35208 26628
rect 34008 25116 35208 25126
rect 34064 25114 34112 25116
rect 34168 25114 34216 25116
rect 34076 25062 34112 25114
rect 34200 25062 34216 25114
rect 34064 25060 34112 25062
rect 34168 25060 34216 25062
rect 34272 25114 34320 25116
rect 34376 25114 34424 25116
rect 34480 25114 34528 25116
rect 34376 25062 34396 25114
rect 34480 25062 34520 25114
rect 34272 25060 34320 25062
rect 34376 25060 34424 25062
rect 34480 25060 34528 25062
rect 34584 25060 34632 25116
rect 34688 25114 34736 25116
rect 34792 25114 34840 25116
rect 34896 25114 34944 25116
rect 34696 25062 34736 25114
rect 34820 25062 34840 25114
rect 34688 25060 34736 25062
rect 34792 25060 34840 25062
rect 34896 25060 34944 25062
rect 35000 25114 35048 25116
rect 35104 25114 35152 25116
rect 35000 25062 35016 25114
rect 35104 25062 35140 25114
rect 35000 25060 35048 25062
rect 35104 25060 35152 25062
rect 34008 25050 35208 25060
rect 34008 23548 35208 23558
rect 34064 23546 34112 23548
rect 34168 23546 34216 23548
rect 34076 23494 34112 23546
rect 34200 23494 34216 23546
rect 34064 23492 34112 23494
rect 34168 23492 34216 23494
rect 34272 23546 34320 23548
rect 34376 23546 34424 23548
rect 34480 23546 34528 23548
rect 34376 23494 34396 23546
rect 34480 23494 34520 23546
rect 34272 23492 34320 23494
rect 34376 23492 34424 23494
rect 34480 23492 34528 23494
rect 34584 23492 34632 23548
rect 34688 23546 34736 23548
rect 34792 23546 34840 23548
rect 34896 23546 34944 23548
rect 34696 23494 34736 23546
rect 34820 23494 34840 23546
rect 34688 23492 34736 23494
rect 34792 23492 34840 23494
rect 34896 23492 34944 23494
rect 35000 23546 35048 23548
rect 35104 23546 35152 23548
rect 35000 23494 35016 23546
rect 35104 23494 35140 23546
rect 35000 23492 35048 23494
rect 35104 23492 35152 23494
rect 34008 23482 35208 23492
rect 34008 21980 35208 21990
rect 34064 21978 34112 21980
rect 34168 21978 34216 21980
rect 34076 21926 34112 21978
rect 34200 21926 34216 21978
rect 34064 21924 34112 21926
rect 34168 21924 34216 21926
rect 34272 21978 34320 21980
rect 34376 21978 34424 21980
rect 34480 21978 34528 21980
rect 34376 21926 34396 21978
rect 34480 21926 34520 21978
rect 34272 21924 34320 21926
rect 34376 21924 34424 21926
rect 34480 21924 34528 21926
rect 34584 21924 34632 21980
rect 34688 21978 34736 21980
rect 34792 21978 34840 21980
rect 34896 21978 34944 21980
rect 34696 21926 34736 21978
rect 34820 21926 34840 21978
rect 34688 21924 34736 21926
rect 34792 21924 34840 21926
rect 34896 21924 34944 21926
rect 35000 21978 35048 21980
rect 35104 21978 35152 21980
rect 35000 21926 35016 21978
rect 35104 21926 35140 21978
rect 35000 21924 35048 21926
rect 35104 21924 35152 21926
rect 34008 21914 35208 21924
rect 34008 20412 35208 20422
rect 34064 20410 34112 20412
rect 34168 20410 34216 20412
rect 34076 20358 34112 20410
rect 34200 20358 34216 20410
rect 34064 20356 34112 20358
rect 34168 20356 34216 20358
rect 34272 20410 34320 20412
rect 34376 20410 34424 20412
rect 34480 20410 34528 20412
rect 34376 20358 34396 20410
rect 34480 20358 34520 20410
rect 34272 20356 34320 20358
rect 34376 20356 34424 20358
rect 34480 20356 34528 20358
rect 34584 20356 34632 20412
rect 34688 20410 34736 20412
rect 34792 20410 34840 20412
rect 34896 20410 34944 20412
rect 34696 20358 34736 20410
rect 34820 20358 34840 20410
rect 34688 20356 34736 20358
rect 34792 20356 34840 20358
rect 34896 20356 34944 20358
rect 35000 20410 35048 20412
rect 35104 20410 35152 20412
rect 35000 20358 35016 20410
rect 35104 20358 35140 20410
rect 35000 20356 35048 20358
rect 35104 20356 35152 20358
rect 34008 20346 35208 20356
rect 34008 18844 35208 18854
rect 34064 18842 34112 18844
rect 34168 18842 34216 18844
rect 34076 18790 34112 18842
rect 34200 18790 34216 18842
rect 34064 18788 34112 18790
rect 34168 18788 34216 18790
rect 34272 18842 34320 18844
rect 34376 18842 34424 18844
rect 34480 18842 34528 18844
rect 34376 18790 34396 18842
rect 34480 18790 34520 18842
rect 34272 18788 34320 18790
rect 34376 18788 34424 18790
rect 34480 18788 34528 18790
rect 34584 18788 34632 18844
rect 34688 18842 34736 18844
rect 34792 18842 34840 18844
rect 34896 18842 34944 18844
rect 34696 18790 34736 18842
rect 34820 18790 34840 18842
rect 34688 18788 34736 18790
rect 34792 18788 34840 18790
rect 34896 18788 34944 18790
rect 35000 18842 35048 18844
rect 35104 18842 35152 18844
rect 35000 18790 35016 18842
rect 35104 18790 35140 18842
rect 35000 18788 35048 18790
rect 35104 18788 35152 18790
rect 34008 18778 35208 18788
rect 34008 17276 35208 17286
rect 34064 17274 34112 17276
rect 34168 17274 34216 17276
rect 34076 17222 34112 17274
rect 34200 17222 34216 17274
rect 34064 17220 34112 17222
rect 34168 17220 34216 17222
rect 34272 17274 34320 17276
rect 34376 17274 34424 17276
rect 34480 17274 34528 17276
rect 34376 17222 34396 17274
rect 34480 17222 34520 17274
rect 34272 17220 34320 17222
rect 34376 17220 34424 17222
rect 34480 17220 34528 17222
rect 34584 17220 34632 17276
rect 34688 17274 34736 17276
rect 34792 17274 34840 17276
rect 34896 17274 34944 17276
rect 34696 17222 34736 17274
rect 34820 17222 34840 17274
rect 34688 17220 34736 17222
rect 34792 17220 34840 17222
rect 34896 17220 34944 17222
rect 35000 17274 35048 17276
rect 35104 17274 35152 17276
rect 35000 17222 35016 17274
rect 35104 17222 35140 17274
rect 35000 17220 35048 17222
rect 35104 17220 35152 17222
rect 34008 17210 35208 17220
rect 34008 15708 35208 15718
rect 34064 15706 34112 15708
rect 34168 15706 34216 15708
rect 34076 15654 34112 15706
rect 34200 15654 34216 15706
rect 34064 15652 34112 15654
rect 34168 15652 34216 15654
rect 34272 15706 34320 15708
rect 34376 15706 34424 15708
rect 34480 15706 34528 15708
rect 34376 15654 34396 15706
rect 34480 15654 34520 15706
rect 34272 15652 34320 15654
rect 34376 15652 34424 15654
rect 34480 15652 34528 15654
rect 34584 15652 34632 15708
rect 34688 15706 34736 15708
rect 34792 15706 34840 15708
rect 34896 15706 34944 15708
rect 34696 15654 34736 15706
rect 34820 15654 34840 15706
rect 34688 15652 34736 15654
rect 34792 15652 34840 15654
rect 34896 15652 34944 15654
rect 35000 15706 35048 15708
rect 35104 15706 35152 15708
rect 35000 15654 35016 15706
rect 35104 15654 35140 15706
rect 35000 15652 35048 15654
rect 35104 15652 35152 15654
rect 34008 15642 35208 15652
rect 34008 14140 35208 14150
rect 34064 14138 34112 14140
rect 34168 14138 34216 14140
rect 34076 14086 34112 14138
rect 34200 14086 34216 14138
rect 34064 14084 34112 14086
rect 34168 14084 34216 14086
rect 34272 14138 34320 14140
rect 34376 14138 34424 14140
rect 34480 14138 34528 14140
rect 34376 14086 34396 14138
rect 34480 14086 34520 14138
rect 34272 14084 34320 14086
rect 34376 14084 34424 14086
rect 34480 14084 34528 14086
rect 34584 14084 34632 14140
rect 34688 14138 34736 14140
rect 34792 14138 34840 14140
rect 34896 14138 34944 14140
rect 34696 14086 34736 14138
rect 34820 14086 34840 14138
rect 34688 14084 34736 14086
rect 34792 14084 34840 14086
rect 34896 14084 34944 14086
rect 35000 14138 35048 14140
rect 35104 14138 35152 14140
rect 35000 14086 35016 14138
rect 35104 14086 35140 14138
rect 35000 14084 35048 14086
rect 35104 14084 35152 14086
rect 34008 14074 35208 14084
rect 34008 12572 35208 12582
rect 34064 12570 34112 12572
rect 34168 12570 34216 12572
rect 34076 12518 34112 12570
rect 34200 12518 34216 12570
rect 34064 12516 34112 12518
rect 34168 12516 34216 12518
rect 34272 12570 34320 12572
rect 34376 12570 34424 12572
rect 34480 12570 34528 12572
rect 34376 12518 34396 12570
rect 34480 12518 34520 12570
rect 34272 12516 34320 12518
rect 34376 12516 34424 12518
rect 34480 12516 34528 12518
rect 34584 12516 34632 12572
rect 34688 12570 34736 12572
rect 34792 12570 34840 12572
rect 34896 12570 34944 12572
rect 34696 12518 34736 12570
rect 34820 12518 34840 12570
rect 34688 12516 34736 12518
rect 34792 12516 34840 12518
rect 34896 12516 34944 12518
rect 35000 12570 35048 12572
rect 35104 12570 35152 12572
rect 35000 12518 35016 12570
rect 35104 12518 35140 12570
rect 35000 12516 35048 12518
rect 35104 12516 35152 12518
rect 34008 12506 35208 12516
rect 34008 11004 35208 11014
rect 34064 11002 34112 11004
rect 34168 11002 34216 11004
rect 34076 10950 34112 11002
rect 34200 10950 34216 11002
rect 34064 10948 34112 10950
rect 34168 10948 34216 10950
rect 34272 11002 34320 11004
rect 34376 11002 34424 11004
rect 34480 11002 34528 11004
rect 34376 10950 34396 11002
rect 34480 10950 34520 11002
rect 34272 10948 34320 10950
rect 34376 10948 34424 10950
rect 34480 10948 34528 10950
rect 34584 10948 34632 11004
rect 34688 11002 34736 11004
rect 34792 11002 34840 11004
rect 34896 11002 34944 11004
rect 34696 10950 34736 11002
rect 34820 10950 34840 11002
rect 34688 10948 34736 10950
rect 34792 10948 34840 10950
rect 34896 10948 34944 10950
rect 35000 11002 35048 11004
rect 35104 11002 35152 11004
rect 35000 10950 35016 11002
rect 35104 10950 35140 11002
rect 35000 10948 35048 10950
rect 35104 10948 35152 10950
rect 34008 10938 35208 10948
rect 37436 10500 37492 45612
rect 38220 43316 38276 43326
rect 38220 43222 38276 43260
rect 37660 31556 37716 31566
rect 37660 31462 37716 31500
rect 37884 31554 37940 31566
rect 37884 31502 37886 31554
rect 37938 31502 37940 31554
rect 37436 10434 37492 10444
rect 37884 9716 37940 31502
rect 38220 31556 38276 31566
rect 38220 30996 38276 31500
rect 38220 30930 38276 30940
rect 38220 19010 38276 19022
rect 38220 18958 38222 19010
rect 38274 18958 38276 19010
rect 38220 18676 38276 18958
rect 38220 18610 38276 18620
rect 37884 9650 37940 9660
rect 34008 9436 35208 9446
rect 34064 9434 34112 9436
rect 34168 9434 34216 9436
rect 34076 9382 34112 9434
rect 34200 9382 34216 9434
rect 34064 9380 34112 9382
rect 34168 9380 34216 9382
rect 34272 9434 34320 9436
rect 34376 9434 34424 9436
rect 34480 9434 34528 9436
rect 34376 9382 34396 9434
rect 34480 9382 34520 9434
rect 34272 9380 34320 9382
rect 34376 9380 34424 9382
rect 34480 9380 34528 9382
rect 34584 9380 34632 9436
rect 34688 9434 34736 9436
rect 34792 9434 34840 9436
rect 34896 9434 34944 9436
rect 34696 9382 34736 9434
rect 34820 9382 34840 9434
rect 34688 9380 34736 9382
rect 34792 9380 34840 9382
rect 34896 9380 34944 9382
rect 35000 9434 35048 9436
rect 35104 9434 35152 9436
rect 35000 9382 35016 9434
rect 35104 9382 35140 9434
rect 35000 9380 35048 9382
rect 35104 9380 35152 9382
rect 34008 9370 35208 9380
rect 28364 7970 28420 7980
rect 37884 8372 37940 8382
rect 14008 7868 15208 7878
rect 14064 7866 14112 7868
rect 14168 7866 14216 7868
rect 14076 7814 14112 7866
rect 14200 7814 14216 7866
rect 14064 7812 14112 7814
rect 14168 7812 14216 7814
rect 14272 7866 14320 7868
rect 14376 7866 14424 7868
rect 14480 7866 14528 7868
rect 14376 7814 14396 7866
rect 14480 7814 14520 7866
rect 14272 7812 14320 7814
rect 14376 7812 14424 7814
rect 14480 7812 14528 7814
rect 14584 7812 14632 7868
rect 14688 7866 14736 7868
rect 14792 7866 14840 7868
rect 14896 7866 14944 7868
rect 14696 7814 14736 7866
rect 14820 7814 14840 7866
rect 14688 7812 14736 7814
rect 14792 7812 14840 7814
rect 14896 7812 14944 7814
rect 15000 7866 15048 7868
rect 15104 7866 15152 7868
rect 15000 7814 15016 7866
rect 15104 7814 15140 7866
rect 15000 7812 15048 7814
rect 15104 7812 15152 7814
rect 14008 7802 15208 7812
rect 34008 7868 35208 7878
rect 34064 7866 34112 7868
rect 34168 7866 34216 7868
rect 34076 7814 34112 7866
rect 34200 7814 34216 7866
rect 34064 7812 34112 7814
rect 34168 7812 34216 7814
rect 34272 7866 34320 7868
rect 34376 7866 34424 7868
rect 34480 7866 34528 7868
rect 34376 7814 34396 7866
rect 34480 7814 34520 7866
rect 34272 7812 34320 7814
rect 34376 7812 34424 7814
rect 34480 7812 34528 7814
rect 34584 7812 34632 7868
rect 34688 7866 34736 7868
rect 34792 7866 34840 7868
rect 34896 7866 34944 7868
rect 34696 7814 34736 7866
rect 34820 7814 34840 7866
rect 34688 7812 34736 7814
rect 34792 7812 34840 7814
rect 34896 7812 34944 7814
rect 35000 7866 35048 7868
rect 35104 7866 35152 7868
rect 35000 7814 35016 7866
rect 35104 7814 35140 7866
rect 35000 7812 35048 7814
rect 35104 7812 35152 7814
rect 34008 7802 35208 7812
rect 13804 7522 13860 7532
rect 14700 7700 14756 7710
rect 13580 7074 13636 7084
rect 13692 7474 13748 7486
rect 13692 7422 13694 7474
rect 13746 7422 13748 7474
rect 13692 7364 13748 7422
rect 14700 7476 14756 7644
rect 14700 7382 14756 7420
rect 17612 7588 17668 7598
rect 13468 6692 13524 6702
rect 13468 6598 13524 6636
rect 13356 6514 13412 6524
rect 13580 6578 13636 6590
rect 13580 6526 13582 6578
rect 13634 6526 13636 6578
rect 13132 6300 13524 6356
rect 12460 3444 12516 3482
rect 12460 3378 12516 3388
rect 13020 3388 13076 3612
rect 13468 3666 13524 6300
rect 13580 5236 13636 6526
rect 13580 5170 13636 5180
rect 13580 5012 13636 5022
rect 13580 4452 13636 4956
rect 13580 4338 13636 4396
rect 13580 4286 13582 4338
rect 13634 4286 13636 4338
rect 13580 4274 13636 4286
rect 13692 4116 13748 7308
rect 14252 7362 14308 7374
rect 14252 7310 14254 7362
rect 14306 7310 14308 7362
rect 14028 7250 14084 7262
rect 14028 7198 14030 7250
rect 14082 7198 14084 7250
rect 13804 7140 13860 7150
rect 14028 7140 14084 7198
rect 14252 7250 14308 7310
rect 14252 7198 14254 7250
rect 14306 7198 14308 7250
rect 14252 7186 14308 7198
rect 15148 7362 15204 7374
rect 15148 7310 15150 7362
rect 15202 7310 15204 7362
rect 13860 7084 14084 7140
rect 13804 6132 13860 7084
rect 15148 6580 15204 7310
rect 15596 7362 15652 7374
rect 15596 7310 15598 7362
rect 15650 7310 15652 7362
rect 15596 7250 15652 7310
rect 15596 7198 15598 7250
rect 15650 7198 15652 7250
rect 15596 7186 15652 7198
rect 17612 6802 17668 7532
rect 24008 7084 25208 7094
rect 24064 7082 24112 7084
rect 24168 7082 24216 7084
rect 24076 7030 24112 7082
rect 24200 7030 24216 7082
rect 24064 7028 24112 7030
rect 24168 7028 24216 7030
rect 24272 7082 24320 7084
rect 24376 7082 24424 7084
rect 24480 7082 24528 7084
rect 24376 7030 24396 7082
rect 24480 7030 24520 7082
rect 24272 7028 24320 7030
rect 24376 7028 24424 7030
rect 24480 7028 24528 7030
rect 24584 7028 24632 7084
rect 24688 7082 24736 7084
rect 24792 7082 24840 7084
rect 24896 7082 24944 7084
rect 24696 7030 24736 7082
rect 24820 7030 24840 7082
rect 24688 7028 24736 7030
rect 24792 7028 24840 7030
rect 24896 7028 24944 7030
rect 25000 7082 25048 7084
rect 25104 7082 25152 7084
rect 25000 7030 25016 7082
rect 25104 7030 25140 7082
rect 25000 7028 25048 7030
rect 25104 7028 25152 7030
rect 24008 7018 25208 7028
rect 17612 6750 17614 6802
rect 17666 6750 17668 6802
rect 17612 6738 17668 6750
rect 15484 6692 15540 6702
rect 20524 6692 20580 6702
rect 15484 6690 15764 6692
rect 15484 6638 15486 6690
rect 15538 6638 15764 6690
rect 15484 6636 15764 6638
rect 15484 6626 15540 6636
rect 15148 6514 15204 6524
rect 15484 6466 15540 6478
rect 15484 6414 15486 6466
rect 15538 6414 15540 6466
rect 14008 6300 15208 6310
rect 14064 6298 14112 6300
rect 14168 6298 14216 6300
rect 14076 6246 14112 6298
rect 14200 6246 14216 6298
rect 14064 6244 14112 6246
rect 14168 6244 14216 6246
rect 14272 6298 14320 6300
rect 14376 6298 14424 6300
rect 14480 6298 14528 6300
rect 14376 6246 14396 6298
rect 14480 6246 14520 6298
rect 14272 6244 14320 6246
rect 14376 6244 14424 6246
rect 14480 6244 14528 6246
rect 14584 6244 14632 6300
rect 14688 6298 14736 6300
rect 14792 6298 14840 6300
rect 14896 6298 14944 6300
rect 14696 6246 14736 6298
rect 14820 6246 14840 6298
rect 14688 6244 14736 6246
rect 14792 6244 14840 6246
rect 14896 6244 14944 6246
rect 15000 6298 15048 6300
rect 15104 6298 15152 6300
rect 15000 6246 15016 6298
rect 15104 6246 15140 6298
rect 15000 6244 15048 6246
rect 15104 6244 15152 6246
rect 14008 6234 15208 6244
rect 13804 6076 13972 6132
rect 13692 4050 13748 4060
rect 13804 5796 13860 5806
rect 13804 5122 13860 5740
rect 13804 5070 13806 5122
rect 13858 5070 13860 5122
rect 13468 3614 13470 3666
rect 13522 3614 13524 3666
rect 13468 3602 13524 3614
rect 13020 3332 13300 3388
rect 13244 800 13300 3332
rect 13804 980 13860 5070
rect 13916 5012 13972 6076
rect 14812 5908 14868 5918
rect 14812 5814 14868 5852
rect 15372 5908 15428 5918
rect 15372 5814 15428 5852
rect 14364 5124 14420 5134
rect 13916 4946 13972 4956
rect 14028 5122 14420 5124
rect 14028 5070 14366 5122
rect 14418 5070 14420 5122
rect 14028 5068 14420 5070
rect 14028 5010 14084 5068
rect 14364 5058 14420 5068
rect 14028 4958 14030 5010
rect 14082 4958 14084 5010
rect 14028 4946 14084 4958
rect 15148 4900 15204 4910
rect 15148 4898 15428 4900
rect 15148 4846 15150 4898
rect 15202 4846 15428 4898
rect 15148 4844 15428 4846
rect 15148 4834 15204 4844
rect 14008 4732 15208 4742
rect 14064 4730 14112 4732
rect 14168 4730 14216 4732
rect 14076 4678 14112 4730
rect 14200 4678 14216 4730
rect 14064 4676 14112 4678
rect 14168 4676 14216 4678
rect 14272 4730 14320 4732
rect 14376 4730 14424 4732
rect 14480 4730 14528 4732
rect 14376 4678 14396 4730
rect 14480 4678 14520 4730
rect 14272 4676 14320 4678
rect 14376 4676 14424 4678
rect 14480 4676 14528 4678
rect 14584 4676 14632 4732
rect 14688 4730 14736 4732
rect 14792 4730 14840 4732
rect 14896 4730 14944 4732
rect 14696 4678 14736 4730
rect 14820 4678 14840 4730
rect 14688 4676 14736 4678
rect 14792 4676 14840 4678
rect 14896 4676 14944 4678
rect 15000 4730 15048 4732
rect 15104 4730 15152 4732
rect 15000 4678 15016 4730
rect 15104 4678 15140 4730
rect 15000 4676 15048 4678
rect 15104 4676 15152 4678
rect 14008 4666 15208 4676
rect 14812 4564 14868 4574
rect 14700 4450 14756 4462
rect 14700 4398 14702 4450
rect 14754 4398 14756 4450
rect 14700 4116 14756 4398
rect 14700 4050 14756 4060
rect 14028 3780 14084 3790
rect 14028 3554 14084 3724
rect 14028 3502 14030 3554
rect 14082 3502 14084 3554
rect 14028 3490 14084 3502
rect 14812 3444 14868 4508
rect 15372 4452 15428 4844
rect 15484 4564 15540 6414
rect 15596 5010 15652 5022
rect 15596 4958 15598 5010
rect 15650 4958 15652 5010
rect 15596 4564 15652 4958
rect 15708 4788 15764 6636
rect 20524 6598 20580 6636
rect 21420 6692 21476 6702
rect 21420 6598 21476 6636
rect 36428 6692 36484 6702
rect 16044 6578 16100 6590
rect 16044 6526 16046 6578
rect 16098 6526 16100 6578
rect 15708 4722 15764 4732
rect 15820 5794 15876 5806
rect 15820 5742 15822 5794
rect 15874 5742 15876 5794
rect 15820 4676 15876 5742
rect 16044 4900 16100 6526
rect 17388 6580 17444 6590
rect 16380 5908 16436 5918
rect 16156 5796 16212 5806
rect 16156 5702 16212 5740
rect 16044 4834 16100 4844
rect 16268 5124 16324 5134
rect 15820 4620 16100 4676
rect 15708 4564 15764 4574
rect 15596 4508 15708 4564
rect 15484 4498 15540 4508
rect 15708 4498 15764 4508
rect 15260 4396 15428 4452
rect 15260 3556 15316 4396
rect 16044 4340 16100 4620
rect 15260 3462 15316 3500
rect 15372 4338 16100 4340
rect 15372 4286 16046 4338
rect 16098 4286 16100 4338
rect 15372 4284 16100 4286
rect 14812 3378 14868 3388
rect 14008 3164 15208 3174
rect 14064 3162 14112 3164
rect 14168 3162 14216 3164
rect 14076 3110 14112 3162
rect 14200 3110 14216 3162
rect 14064 3108 14112 3110
rect 14168 3108 14216 3110
rect 14272 3162 14320 3164
rect 14376 3162 14424 3164
rect 14480 3162 14528 3164
rect 14376 3110 14396 3162
rect 14480 3110 14520 3162
rect 14272 3108 14320 3110
rect 14376 3108 14424 3110
rect 14480 3108 14528 3110
rect 14584 3108 14632 3164
rect 14688 3162 14736 3164
rect 14792 3162 14840 3164
rect 14896 3162 14944 3164
rect 14696 3110 14736 3162
rect 14820 3110 14840 3162
rect 14688 3108 14736 3110
rect 14792 3108 14840 3110
rect 14896 3108 14944 3110
rect 15000 3162 15048 3164
rect 15104 3162 15152 3164
rect 15000 3110 15016 3162
rect 15104 3110 15140 3162
rect 15000 3108 15048 3110
rect 15104 3108 15152 3110
rect 14008 3098 15208 3108
rect 15372 2996 15428 4284
rect 16044 4274 16100 4284
rect 16156 3556 16212 3566
rect 16268 3556 16324 5068
rect 16380 4900 16436 5852
rect 16828 5796 16884 5806
rect 16828 5794 17332 5796
rect 16828 5742 16830 5794
rect 16882 5742 17332 5794
rect 16828 5740 17332 5742
rect 16828 5730 16884 5740
rect 16604 5124 16660 5134
rect 16604 5122 16884 5124
rect 16604 5070 16606 5122
rect 16658 5070 16884 5122
rect 16604 5068 16884 5070
rect 16604 5058 16660 5068
rect 16380 4834 16436 4844
rect 16492 5012 16548 5022
rect 16380 4564 16436 4574
rect 16380 4470 16436 4508
rect 16156 3554 16324 3556
rect 16156 3502 16158 3554
rect 16210 3502 16324 3554
rect 16156 3500 16324 3502
rect 16156 3388 16212 3500
rect 15036 2940 15428 2996
rect 15932 3332 16212 3388
rect 16380 3444 16436 3454
rect 16492 3444 16548 4956
rect 16716 4900 16772 4910
rect 16716 4228 16772 4844
rect 16716 4162 16772 4172
rect 16380 3442 16548 3444
rect 16380 3390 16382 3442
rect 16434 3390 16548 3442
rect 16380 3388 16548 3390
rect 16828 3444 16884 5068
rect 17052 5012 17108 5022
rect 17052 4918 17108 4956
rect 16940 4226 16996 4238
rect 16940 4174 16942 4226
rect 16994 4174 16996 4226
rect 16940 3892 16996 4174
rect 16940 3826 16996 3836
rect 17276 3554 17332 5740
rect 17388 4450 17444 6524
rect 19740 6580 19796 6590
rect 19740 6486 19796 6524
rect 20748 6580 20804 6590
rect 20748 6130 20804 6524
rect 34008 6300 35208 6310
rect 34064 6298 34112 6300
rect 34168 6298 34216 6300
rect 34076 6246 34112 6298
rect 34200 6246 34216 6298
rect 34064 6244 34112 6246
rect 34168 6244 34216 6246
rect 34272 6298 34320 6300
rect 34376 6298 34424 6300
rect 34480 6298 34528 6300
rect 34376 6246 34396 6298
rect 34480 6246 34520 6298
rect 34272 6244 34320 6246
rect 34376 6244 34424 6246
rect 34480 6244 34528 6246
rect 34584 6244 34632 6300
rect 34688 6298 34736 6300
rect 34792 6298 34840 6300
rect 34896 6298 34944 6300
rect 34696 6246 34736 6298
rect 34820 6246 34840 6298
rect 34688 6244 34736 6246
rect 34792 6244 34840 6246
rect 34896 6244 34944 6246
rect 35000 6298 35048 6300
rect 35104 6298 35152 6300
rect 35000 6246 35016 6298
rect 35104 6246 35140 6298
rect 35000 6244 35048 6246
rect 35104 6244 35152 6246
rect 34008 6234 35208 6244
rect 20748 6078 20750 6130
rect 20802 6078 20804 6130
rect 20748 6066 20804 6078
rect 17500 5794 17556 5806
rect 17500 5742 17502 5794
rect 17554 5742 17556 5794
rect 17500 5124 17556 5742
rect 17500 5058 17556 5068
rect 17948 5794 18004 5806
rect 24332 5796 24388 5806
rect 17948 5742 17950 5794
rect 18002 5742 18004 5794
rect 17388 4398 17390 4450
rect 17442 4398 17444 4450
rect 17388 4386 17444 4398
rect 17724 4226 17780 4238
rect 17724 4174 17726 4226
rect 17778 4174 17780 4226
rect 17724 3892 17780 4174
rect 17724 3826 17780 3836
rect 17276 3502 17278 3554
rect 17330 3502 17332 3554
rect 17052 3444 17108 3454
rect 16828 3442 17108 3444
rect 16828 3390 17054 3442
rect 17106 3390 17108 3442
rect 16828 3388 17108 3390
rect 16380 3378 16436 3388
rect 17052 3378 17108 3388
rect 13804 924 14196 980
rect 14140 800 14196 924
rect 15036 800 15092 2940
rect 15932 800 15988 3332
rect 17276 3108 17332 3502
rect 17948 3554 18004 5742
rect 23884 5794 24388 5796
rect 23884 5742 24334 5794
rect 24386 5742 24388 5794
rect 23884 5740 24388 5742
rect 22204 5124 22260 5134
rect 21868 5122 22260 5124
rect 21868 5070 22206 5122
rect 22258 5070 22260 5122
rect 21868 5068 22260 5070
rect 18732 4898 18788 4910
rect 18732 4846 18734 4898
rect 18786 4846 18788 4898
rect 17948 3502 17950 3554
rect 18002 3502 18004 3554
rect 17948 3388 18004 3502
rect 16828 3052 17332 3108
rect 17724 3332 18004 3388
rect 18284 4338 18340 4350
rect 18284 4286 18286 4338
rect 18338 4286 18340 4338
rect 18284 3442 18340 4286
rect 18620 4226 18676 4238
rect 18620 4174 18622 4226
rect 18674 4174 18676 4226
rect 18620 3780 18676 4174
rect 18620 3714 18676 3724
rect 18284 3390 18286 3442
rect 18338 3390 18340 3442
rect 18284 3378 18340 3390
rect 18732 3556 18788 4846
rect 19516 4898 19572 4910
rect 20524 4900 20580 4910
rect 19516 4846 19518 4898
rect 19570 4846 19572 4898
rect 19404 4452 19460 4462
rect 19180 4450 19460 4452
rect 19180 4398 19406 4450
rect 19458 4398 19460 4450
rect 19180 4396 19460 4398
rect 18844 3556 18900 3566
rect 18732 3554 18900 3556
rect 18732 3502 18846 3554
rect 18898 3502 18900 3554
rect 18732 3500 18900 3502
rect 18732 3388 18788 3500
rect 18844 3490 18900 3500
rect 18620 3332 18788 3388
rect 19180 3442 19236 4396
rect 19404 4386 19460 4396
rect 19180 3390 19182 3442
rect 19234 3390 19236 3442
rect 19180 3378 19236 3390
rect 19516 3556 19572 4846
rect 20300 4898 20580 4900
rect 20300 4846 20526 4898
rect 20578 4846 20580 4898
rect 20300 4844 20580 4846
rect 20076 4452 20132 4462
rect 19740 3556 19796 3566
rect 19516 3554 19796 3556
rect 19516 3502 19742 3554
rect 19794 3502 19796 3554
rect 19516 3500 19796 3502
rect 16828 800 16884 3052
rect 17724 800 17780 3332
rect 18620 800 18676 3332
rect 19516 800 19572 3500
rect 19740 3490 19796 3500
rect 20076 3442 20132 4396
rect 20076 3390 20078 3442
rect 20130 3390 20132 3442
rect 20076 3378 20132 3390
rect 20300 3388 20356 4844
rect 20524 4834 20580 4844
rect 21532 4898 21588 4910
rect 21532 4846 21534 4898
rect 21586 4846 21588 4898
rect 20860 4452 20916 4462
rect 20860 4358 20916 4396
rect 20412 4340 20468 4350
rect 20412 4338 20804 4340
rect 20412 4286 20414 4338
rect 20466 4286 20804 4338
rect 20412 4284 20804 4286
rect 20412 4274 20468 4284
rect 20748 3892 20804 4284
rect 20748 3836 21140 3892
rect 20748 3442 20804 3454
rect 20748 3390 20750 3442
rect 20802 3390 20804 3442
rect 20748 3388 20804 3390
rect 20300 3332 20804 3388
rect 21084 3442 21140 3836
rect 21084 3390 21086 3442
rect 21138 3390 21140 3442
rect 21084 3378 21140 3390
rect 21532 3554 21588 4846
rect 21532 3502 21534 3554
rect 21586 3502 21588 3554
rect 21532 3388 21588 3502
rect 21308 3332 21588 3388
rect 21868 3442 21924 5068
rect 22204 5058 22260 5068
rect 22876 5010 22932 5022
rect 22876 4958 22878 5010
rect 22930 4958 22932 5010
rect 21980 4900 22036 4910
rect 21980 4898 22260 4900
rect 21980 4846 21982 4898
rect 22034 4846 22260 4898
rect 21980 4844 22260 4846
rect 21980 4834 22036 4844
rect 21868 3390 21870 3442
rect 21922 3390 21924 3442
rect 21868 3378 21924 3390
rect 22204 3556 22260 4844
rect 22764 4116 22820 4126
rect 22764 4022 22820 4060
rect 22428 3556 22484 3566
rect 22204 3554 22484 3556
rect 22204 3502 22430 3554
rect 22482 3502 22484 3554
rect 22204 3500 22484 3502
rect 20412 800 20468 3332
rect 21308 800 21364 3332
rect 22204 800 22260 3500
rect 22428 3490 22484 3500
rect 22764 3444 22820 3454
rect 22876 3444 22932 4958
rect 23660 5012 23716 5022
rect 22764 3442 22932 3444
rect 22764 3390 22766 3442
rect 22818 3390 22932 3442
rect 22764 3388 22932 3390
rect 23436 4116 23492 4126
rect 23436 3554 23492 4060
rect 23436 3502 23438 3554
rect 23490 3502 23492 3554
rect 23436 3388 23492 3502
rect 22764 3378 22820 3388
rect 23100 3332 23492 3388
rect 23660 3442 23716 4956
rect 23772 4898 23828 4910
rect 23772 4846 23774 4898
rect 23826 4846 23828 4898
rect 23772 4450 23828 4846
rect 23772 4398 23774 4450
rect 23826 4398 23828 4450
rect 23772 4386 23828 4398
rect 23660 3390 23662 3442
rect 23714 3390 23716 3442
rect 23660 3378 23716 3390
rect 23100 800 23156 3332
rect 23884 3220 23940 5740
rect 24332 5730 24388 5740
rect 24008 5516 25208 5526
rect 24064 5514 24112 5516
rect 24168 5514 24216 5516
rect 24076 5462 24112 5514
rect 24200 5462 24216 5514
rect 24064 5460 24112 5462
rect 24168 5460 24216 5462
rect 24272 5514 24320 5516
rect 24376 5514 24424 5516
rect 24480 5514 24528 5516
rect 24376 5462 24396 5514
rect 24480 5462 24520 5514
rect 24272 5460 24320 5462
rect 24376 5460 24424 5462
rect 24480 5460 24528 5462
rect 24584 5460 24632 5516
rect 24688 5514 24736 5516
rect 24792 5514 24840 5516
rect 24896 5514 24944 5516
rect 24696 5462 24736 5514
rect 24820 5462 24840 5514
rect 24688 5460 24736 5462
rect 24792 5460 24840 5462
rect 24896 5460 24944 5462
rect 25000 5514 25048 5516
rect 25104 5514 25152 5516
rect 25000 5462 25016 5514
rect 25104 5462 25140 5514
rect 25000 5460 25048 5462
rect 25104 5460 25152 5462
rect 24008 5450 25208 5460
rect 26012 5124 26068 5134
rect 25788 5122 26068 5124
rect 25788 5070 26014 5122
rect 26066 5070 26068 5122
rect 25788 5068 26068 5070
rect 24892 5012 24948 5022
rect 24892 4918 24948 4956
rect 24108 4564 24164 4574
rect 24108 4338 24164 4508
rect 25340 4564 25396 4602
rect 25340 4498 25396 4508
rect 24108 4286 24110 4338
rect 24162 4286 24164 4338
rect 24108 4274 24164 4286
rect 25340 4338 25396 4350
rect 25340 4286 25342 4338
rect 25394 4286 25396 4338
rect 24556 4226 24612 4238
rect 24556 4174 24558 4226
rect 24610 4174 24612 4226
rect 24556 4116 24612 4174
rect 24556 4050 24612 4060
rect 24008 3948 25208 3958
rect 24064 3946 24112 3948
rect 24168 3946 24216 3948
rect 24076 3894 24112 3946
rect 24200 3894 24216 3946
rect 24064 3892 24112 3894
rect 24168 3892 24216 3894
rect 24272 3946 24320 3948
rect 24376 3946 24424 3948
rect 24480 3946 24528 3948
rect 24376 3894 24396 3946
rect 24480 3894 24520 3946
rect 24272 3892 24320 3894
rect 24376 3892 24424 3894
rect 24480 3892 24528 3894
rect 24584 3892 24632 3948
rect 24688 3946 24736 3948
rect 24792 3946 24840 3948
rect 24896 3946 24944 3948
rect 24696 3894 24736 3946
rect 24820 3894 24840 3946
rect 24688 3892 24736 3894
rect 24792 3892 24840 3894
rect 24896 3892 24944 3894
rect 25000 3946 25048 3948
rect 25104 3946 25152 3948
rect 25000 3894 25016 3946
rect 25104 3894 25140 3946
rect 25000 3892 25048 3894
rect 25104 3892 25152 3894
rect 24008 3882 25208 3892
rect 25116 3668 25172 3678
rect 24556 3444 24612 3454
rect 24892 3442 24948 3454
rect 24892 3390 24894 3442
rect 24946 3390 24948 3442
rect 24892 3388 24948 3390
rect 24556 3350 24612 3388
rect 24668 3332 24948 3388
rect 25116 3444 25172 3612
rect 25228 3444 25284 3454
rect 25116 3442 25284 3444
rect 25116 3390 25230 3442
rect 25282 3390 25284 3442
rect 25116 3388 25284 3390
rect 25340 3444 25396 4286
rect 25564 3444 25620 3454
rect 25340 3442 25620 3444
rect 25340 3390 25566 3442
rect 25618 3390 25620 3442
rect 25340 3388 25620 3390
rect 24668 3220 24724 3332
rect 23884 3164 24724 3220
rect 23996 924 24388 980
rect 23996 800 24052 924
rect 2464 0 2576 800
rect 3360 0 3472 800
rect 4256 0 4368 800
rect 5152 0 5264 800
rect 6048 0 6160 800
rect 6944 0 7056 800
rect 7840 0 7952 800
rect 8736 0 8848 800
rect 9632 0 9744 800
rect 10528 0 10640 800
rect 11424 0 11536 800
rect 12320 0 12432 800
rect 13216 0 13328 800
rect 14112 0 14224 800
rect 15008 0 15120 800
rect 15904 0 16016 800
rect 16800 0 16912 800
rect 17696 0 17808 800
rect 18592 0 18704 800
rect 19488 0 19600 800
rect 20384 0 20496 800
rect 21280 0 21392 800
rect 22176 0 22288 800
rect 23072 0 23184 800
rect 23968 0 24080 800
rect 24332 756 24388 924
rect 24668 756 24724 3164
rect 25116 2212 25172 3388
rect 25228 3378 25284 3388
rect 25564 3378 25620 3388
rect 25788 3444 25844 5068
rect 26012 5058 26068 5068
rect 28140 5122 28196 5134
rect 28140 5070 28142 5122
rect 28194 5070 28196 5122
rect 26460 4898 26516 4910
rect 26908 4900 26964 4910
rect 26460 4846 26462 4898
rect 26514 4846 26516 4898
rect 25900 4452 25956 4462
rect 25900 4450 26068 4452
rect 25900 4398 25902 4450
rect 25954 4398 26068 4450
rect 25900 4396 26068 4398
rect 25900 4386 25956 4396
rect 25788 3378 25844 3388
rect 26012 3442 26068 4396
rect 26012 3390 26014 3442
rect 26066 3390 26068 3442
rect 26012 3378 26068 3390
rect 26348 3556 26404 3566
rect 26460 3556 26516 4846
rect 26348 3554 26516 3556
rect 26348 3502 26350 3554
rect 26402 3502 26516 3554
rect 26348 3500 26516 3502
rect 26684 4898 26964 4900
rect 26684 4846 26910 4898
rect 26962 4846 26964 4898
rect 26684 4844 26964 4846
rect 26348 3388 26404 3500
rect 26236 3332 26404 3388
rect 26684 3444 26740 4844
rect 26908 4834 26964 4844
rect 26236 2772 26292 3332
rect 24892 2156 25172 2212
rect 25788 2716 26292 2772
rect 24892 800 24948 2156
rect 25788 800 25844 2716
rect 26684 800 26740 3388
rect 26908 4508 27636 4564
rect 26908 3442 26964 4508
rect 27580 4452 27636 4508
rect 27916 4452 27972 4462
rect 27580 4450 27972 4452
rect 27580 4398 27918 4450
rect 27970 4398 27972 4450
rect 27580 4396 27972 4398
rect 27916 4386 27972 4396
rect 27468 4340 27524 4350
rect 27468 4338 27860 4340
rect 27468 4286 27470 4338
rect 27522 4286 27860 4338
rect 27468 4284 27860 4286
rect 27468 4274 27524 4284
rect 27804 3892 27860 4284
rect 28140 4004 28196 5070
rect 30156 5122 30212 5134
rect 32284 5124 32340 5134
rect 30156 5070 30158 5122
rect 30210 5070 30212 5122
rect 29484 4226 29540 4238
rect 29484 4174 29486 4226
rect 29538 4174 29540 4226
rect 29372 4114 29428 4126
rect 29372 4062 29374 4114
rect 29426 4062 29428 4114
rect 28140 3948 28644 4004
rect 27804 3836 28420 3892
rect 27692 3668 27748 3678
rect 27692 3574 27748 3612
rect 26908 3390 26910 3442
rect 26962 3390 26964 3442
rect 26908 3378 26964 3390
rect 27132 3554 27188 3566
rect 27132 3502 27134 3554
rect 27186 3502 27188 3554
rect 27132 3444 27188 3502
rect 27132 3378 27188 3388
rect 27580 3556 27636 3566
rect 27580 800 27636 3500
rect 28364 3442 28420 3836
rect 28588 3556 28644 3948
rect 28588 3462 28644 3500
rect 28364 3390 28366 3442
rect 28418 3390 28420 3442
rect 28364 3378 28420 3390
rect 28476 3444 28532 3454
rect 28476 800 28532 3388
rect 29036 3444 29092 3454
rect 29036 3350 29092 3388
rect 29372 3442 29428 4062
rect 29372 3390 29374 3442
rect 29426 3390 29428 3442
rect 29372 3378 29428 3390
rect 29484 3444 29540 4174
rect 29932 4226 29988 4238
rect 29932 4174 29934 4226
rect 29986 4174 29988 4226
rect 29484 3378 29540 3388
rect 29708 3444 29764 3454
rect 29932 3444 29988 4174
rect 30156 4226 30212 5070
rect 31724 5122 32340 5124
rect 31724 5070 32286 5122
rect 32338 5070 32340 5122
rect 31724 5068 32340 5070
rect 30156 4174 30158 4226
rect 30210 4174 30212 4226
rect 30156 4162 30212 4174
rect 30268 5010 30324 5022
rect 30268 4958 30270 5010
rect 30322 4958 30324 5010
rect 29708 3442 29988 3444
rect 29708 3390 29710 3442
rect 29762 3390 29988 3442
rect 29708 3388 29988 3390
rect 30044 3444 30100 3454
rect 30268 3444 30324 4958
rect 30828 5012 30884 5022
rect 30044 3442 30324 3444
rect 30044 3390 30046 3442
rect 30098 3390 30324 3442
rect 30044 3388 30324 3390
rect 30492 4226 30548 4238
rect 30492 4174 30494 4226
rect 30546 4174 30548 4226
rect 30492 3442 30548 4174
rect 30492 3390 30494 3442
rect 30546 3390 30548 3442
rect 29708 2548 29764 3388
rect 30044 3378 30100 3388
rect 30492 2548 30548 3390
rect 30828 3442 30884 4956
rect 31500 4114 31556 4126
rect 31500 4062 31502 4114
rect 31554 4062 31556 4114
rect 31276 3444 31332 3454
rect 31500 3444 31556 4062
rect 31724 3444 31780 5068
rect 32284 5058 32340 5068
rect 34972 5122 35028 5134
rect 34972 5070 34974 5122
rect 35026 5070 35028 5122
rect 32844 5012 32900 5022
rect 32844 4918 32900 4956
rect 33852 4898 33908 4910
rect 33852 4846 33854 4898
rect 33906 4846 33908 4898
rect 32508 4620 33348 4676
rect 32060 4340 32116 4350
rect 31836 4226 31892 4238
rect 31836 4174 31838 4226
rect 31890 4174 31892 4226
rect 31836 4114 31892 4174
rect 31836 4062 31838 4114
rect 31890 4062 31892 4114
rect 31836 4050 31892 4062
rect 32060 3666 32116 4284
rect 32508 4226 32564 4620
rect 32508 4174 32510 4226
rect 32562 4174 32564 4226
rect 32508 3780 32564 4174
rect 32060 3614 32062 3666
rect 32114 3614 32116 3666
rect 32060 3602 32116 3614
rect 32172 3724 32564 3780
rect 33068 4450 33124 4462
rect 33068 4398 33070 4450
rect 33122 4398 33124 4450
rect 30828 3390 30830 3442
rect 30882 3390 30884 3442
rect 30828 3378 30884 3390
rect 31164 3442 31556 3444
rect 31164 3390 31278 3442
rect 31330 3390 31556 3442
rect 31164 3388 31556 3390
rect 31612 3388 31780 3444
rect 29372 2492 29764 2548
rect 30268 2492 30548 2548
rect 29372 800 29428 2492
rect 30268 800 30324 2492
rect 31164 800 31220 3388
rect 31276 3378 31332 3388
rect 31612 3330 31668 3388
rect 31612 3278 31614 3330
rect 31666 3278 31668 3330
rect 31612 3266 31668 3278
rect 32172 2884 32228 3724
rect 32284 3556 32340 3566
rect 33068 3556 33124 4398
rect 32284 3554 33124 3556
rect 32284 3502 32286 3554
rect 32338 3502 33124 3554
rect 32284 3500 33124 3502
rect 33180 4340 33236 4350
rect 32284 3490 32340 3500
rect 33180 3444 33236 4284
rect 33292 4338 33348 4620
rect 33292 4286 33294 4338
rect 33346 4286 33348 4338
rect 33292 4274 33348 4286
rect 33740 4450 33796 4462
rect 33740 4398 33742 4450
rect 33794 4398 33796 4450
rect 32060 2828 32228 2884
rect 32956 3388 33236 3444
rect 33628 3668 33684 3678
rect 32060 800 32116 2828
rect 32956 800 33012 3388
rect 33628 3220 33684 3612
rect 33740 3442 33796 4398
rect 33740 3390 33742 3442
rect 33794 3390 33796 3442
rect 33740 3378 33796 3390
rect 33852 3444 33908 4846
rect 34412 4900 34468 4938
rect 34972 4900 35028 5070
rect 34972 4844 35364 4900
rect 34412 4834 34468 4844
rect 34008 4732 35208 4742
rect 34064 4730 34112 4732
rect 34168 4730 34216 4732
rect 34076 4678 34112 4730
rect 34200 4678 34216 4730
rect 34064 4676 34112 4678
rect 34168 4676 34216 4678
rect 34272 4730 34320 4732
rect 34376 4730 34424 4732
rect 34480 4730 34528 4732
rect 34376 4678 34396 4730
rect 34480 4678 34520 4730
rect 34272 4676 34320 4678
rect 34376 4676 34424 4678
rect 34480 4676 34528 4678
rect 34584 4676 34632 4732
rect 34688 4730 34736 4732
rect 34792 4730 34840 4732
rect 34896 4730 34944 4732
rect 34696 4678 34736 4730
rect 34820 4678 34840 4730
rect 34688 4676 34736 4678
rect 34792 4676 34840 4678
rect 34896 4676 34944 4678
rect 35000 4730 35048 4732
rect 35104 4730 35152 4732
rect 35000 4678 35016 4730
rect 35104 4678 35140 4730
rect 35000 4676 35048 4678
rect 35104 4676 35152 4678
rect 34008 4666 35208 4676
rect 34748 4452 34804 4462
rect 35084 4452 35140 4462
rect 34748 4450 35140 4452
rect 34748 4398 34750 4450
rect 34802 4398 35086 4450
rect 35138 4398 35140 4450
rect 34748 4396 35140 4398
rect 34748 4386 34804 4396
rect 35084 4386 35140 4396
rect 33964 4340 34020 4350
rect 33964 4246 34020 4284
rect 34412 4340 34468 4350
rect 34412 4246 34468 4284
rect 35308 4338 35364 4844
rect 35308 4286 35310 4338
rect 35362 4286 35364 4338
rect 34412 4114 34468 4126
rect 34412 4062 34414 4114
rect 34466 4062 34468 4114
rect 34412 3554 34468 4062
rect 35308 3668 35364 4286
rect 35756 4340 35812 4350
rect 35812 4284 35924 4340
rect 35756 4274 35812 4284
rect 35308 3602 35364 3612
rect 35644 4228 35700 4238
rect 34412 3502 34414 3554
rect 34466 3502 34468 3554
rect 34412 3490 34468 3502
rect 33852 3378 33908 3388
rect 34524 3444 34580 3454
rect 34524 3350 34580 3388
rect 35308 3444 35364 3454
rect 33628 3164 33908 3220
rect 33852 800 33908 3164
rect 34008 3164 35208 3174
rect 34064 3162 34112 3164
rect 34168 3162 34216 3164
rect 34076 3110 34112 3162
rect 34200 3110 34216 3162
rect 34064 3108 34112 3110
rect 34168 3108 34216 3110
rect 34272 3162 34320 3164
rect 34376 3162 34424 3164
rect 34480 3162 34528 3164
rect 34376 3110 34396 3162
rect 34480 3110 34520 3162
rect 34272 3108 34320 3110
rect 34376 3108 34424 3110
rect 34480 3108 34528 3110
rect 34584 3108 34632 3164
rect 34688 3162 34736 3164
rect 34792 3162 34840 3164
rect 34896 3162 34944 3164
rect 34696 3110 34736 3162
rect 34820 3110 34840 3162
rect 34688 3108 34736 3110
rect 34792 3108 34840 3110
rect 34896 3108 34944 3110
rect 35000 3162 35048 3164
rect 35104 3162 35152 3164
rect 35000 3110 35016 3162
rect 35104 3110 35140 3162
rect 35000 3108 35048 3110
rect 35104 3108 35152 3110
rect 34008 3098 35208 3108
rect 35308 2996 35364 3388
rect 35196 2940 35364 2996
rect 35196 2548 35252 2940
rect 34748 2492 35252 2548
rect 34748 800 34804 2492
rect 35644 800 35700 4172
rect 35868 3444 35924 4284
rect 35980 4226 36036 4238
rect 35980 4174 35982 4226
rect 36034 4174 36036 4226
rect 35980 3556 36036 4174
rect 36204 3556 36260 3566
rect 35980 3554 36260 3556
rect 35980 3502 36206 3554
rect 36258 3502 36260 3554
rect 35980 3500 36260 3502
rect 36204 3444 36260 3500
rect 35868 3388 36036 3444
rect 35980 3330 36036 3388
rect 36428 3444 36484 6636
rect 37884 6578 37940 8316
rect 37884 6526 37886 6578
rect 37938 6526 37940 6578
rect 37884 6514 37940 6526
rect 38220 6578 38276 6590
rect 38220 6526 38222 6578
rect 38274 6526 38276 6578
rect 37660 6466 37716 6478
rect 37660 6414 37662 6466
rect 37714 6414 37716 6466
rect 37660 6356 37716 6414
rect 37660 6290 37716 6300
rect 38220 6356 38276 6526
rect 38220 6290 38276 6300
rect 36540 4226 36596 4238
rect 36540 4174 36542 4226
rect 36594 4174 36596 4226
rect 36540 3556 36596 4174
rect 37436 4226 37492 4238
rect 37436 4174 37438 4226
rect 37490 4174 37492 4226
rect 37212 4116 37268 4126
rect 37268 4060 37380 4116
rect 37212 4050 37268 4060
rect 36988 3556 37044 3566
rect 36540 3554 37044 3556
rect 36540 3502 36990 3554
rect 37042 3502 37044 3554
rect 36540 3500 37044 3502
rect 36428 3388 36820 3444
rect 36204 3378 36260 3388
rect 35980 3278 35982 3330
rect 36034 3278 36036 3330
rect 35980 3266 36036 3278
rect 36764 3330 36820 3388
rect 36764 3278 36766 3330
rect 36818 3278 36820 3330
rect 36764 3266 36820 3278
rect 36876 2548 36932 3500
rect 36988 3490 37044 3500
rect 37324 3444 37380 4060
rect 37436 3556 37492 4174
rect 37884 3556 37940 3566
rect 37436 3554 37940 3556
rect 37436 3502 37886 3554
rect 37938 3502 37940 3554
rect 37436 3500 37940 3502
rect 37324 3388 37716 3444
rect 37660 3330 37716 3388
rect 37660 3278 37662 3330
rect 37714 3278 37716 3330
rect 37660 3266 37716 3278
rect 37884 2548 37940 3500
rect 36540 2492 36932 2548
rect 37436 2492 37940 2548
rect 36540 800 36596 2492
rect 37436 800 37492 2492
rect 24332 700 24724 756
rect 24864 0 24976 800
rect 25760 0 25872 800
rect 26656 0 26768 800
rect 27552 0 27664 800
rect 28448 0 28560 800
rect 29344 0 29456 800
rect 30240 0 30352 800
rect 31136 0 31248 800
rect 32032 0 32144 800
rect 32928 0 33040 800
rect 33824 0 33936 800
rect 34720 0 34832 800
rect 35616 0 35728 800
rect 36512 0 36624 800
rect 37408 0 37520 800
<< via2 >>
rect 2044 46956 2100 47012
rect 4008 46282 4064 46284
rect 4112 46282 4168 46284
rect 4008 46230 4024 46282
rect 4024 46230 4064 46282
rect 4112 46230 4148 46282
rect 4148 46230 4168 46282
rect 4008 46228 4064 46230
rect 4112 46228 4168 46230
rect 4216 46228 4272 46284
rect 4320 46282 4376 46284
rect 4424 46282 4480 46284
rect 4528 46282 4584 46284
rect 4320 46230 4324 46282
rect 4324 46230 4376 46282
rect 4424 46230 4448 46282
rect 4448 46230 4480 46282
rect 4528 46230 4572 46282
rect 4572 46230 4584 46282
rect 4320 46228 4376 46230
rect 4424 46228 4480 46230
rect 4528 46228 4584 46230
rect 4632 46282 4688 46284
rect 4736 46282 4792 46284
rect 4840 46282 4896 46284
rect 4632 46230 4644 46282
rect 4644 46230 4688 46282
rect 4736 46230 4768 46282
rect 4768 46230 4792 46282
rect 4840 46230 4892 46282
rect 4892 46230 4896 46282
rect 4632 46228 4688 46230
rect 4736 46228 4792 46230
rect 4840 46228 4896 46230
rect 4944 46228 5000 46284
rect 5048 46282 5104 46284
rect 5152 46282 5208 46284
rect 5048 46230 5068 46282
rect 5068 46230 5104 46282
rect 5152 46230 5192 46282
rect 5192 46230 5208 46282
rect 5048 46228 5104 46230
rect 5152 46228 5208 46230
rect 2156 45724 2212 45780
rect 1708 44380 1764 44436
rect 1820 44940 1876 44996
rect 1708 43036 1764 43092
rect 1708 41692 1764 41748
rect 1708 40348 1764 40404
rect 1708 39004 1764 39060
rect 1708 37826 1764 37828
rect 1708 37774 1710 37826
rect 1710 37774 1762 37826
rect 1762 37774 1764 37826
rect 1708 37772 1764 37774
rect 1708 36370 1764 36372
rect 1708 36318 1710 36370
rect 1710 36318 1762 36370
rect 1762 36318 1764 36370
rect 1708 36316 1764 36318
rect 1708 34972 1764 35028
rect 1708 33628 1764 33684
rect 1708 32284 1764 32340
rect 1708 30940 1764 30996
rect 1708 29596 1764 29652
rect 1708 28418 1764 28420
rect 1708 28366 1710 28418
rect 1710 28366 1762 28418
rect 1762 28366 1764 28418
rect 1708 28364 1764 28366
rect 1708 26908 1764 26964
rect 1708 25564 1764 25620
rect 1708 24220 1764 24276
rect 1708 22876 1764 22932
rect 1708 21532 1764 21588
rect 1708 20188 1764 20244
rect 1708 19010 1764 19012
rect 1708 18958 1710 19010
rect 1710 18958 1762 19010
rect 1762 18958 1764 19010
rect 1708 18956 1764 18958
rect 1708 17554 1764 17556
rect 1708 17502 1710 17554
rect 1710 17502 1762 17554
rect 1762 17502 1764 17554
rect 1708 17500 1764 17502
rect 1708 16156 1764 16212
rect 1708 14812 1764 14868
rect 1708 13468 1764 13524
rect 1708 12124 1764 12180
rect 1708 10780 1764 10836
rect 1708 9602 1764 9604
rect 1708 9550 1710 9602
rect 1710 9550 1762 9602
rect 1762 9550 1764 9602
rect 1708 9548 1764 9550
rect 1708 8146 1764 8148
rect 1708 8094 1710 8146
rect 1710 8094 1762 8146
rect 1762 8094 1764 8146
rect 1708 8092 1764 8094
rect 2716 44994 2772 44996
rect 2716 44942 2718 44994
rect 2718 44942 2770 44994
rect 2770 44942 2772 44994
rect 2716 44940 2772 44942
rect 12572 45948 12628 46004
rect 13580 46002 13636 46004
rect 13580 45950 13582 46002
rect 13582 45950 13634 46002
rect 13634 45950 13636 46002
rect 13580 45948 13636 45950
rect 3500 44940 3556 44996
rect 4008 44714 4064 44716
rect 4112 44714 4168 44716
rect 4008 44662 4024 44714
rect 4024 44662 4064 44714
rect 4112 44662 4148 44714
rect 4148 44662 4168 44714
rect 4008 44660 4064 44662
rect 4112 44660 4168 44662
rect 4216 44660 4272 44716
rect 4320 44714 4376 44716
rect 4424 44714 4480 44716
rect 4528 44714 4584 44716
rect 4320 44662 4324 44714
rect 4324 44662 4376 44714
rect 4424 44662 4448 44714
rect 4448 44662 4480 44714
rect 4528 44662 4572 44714
rect 4572 44662 4584 44714
rect 4320 44660 4376 44662
rect 4424 44660 4480 44662
rect 4528 44660 4584 44662
rect 4632 44714 4688 44716
rect 4736 44714 4792 44716
rect 4840 44714 4896 44716
rect 4632 44662 4644 44714
rect 4644 44662 4688 44714
rect 4736 44662 4768 44714
rect 4768 44662 4792 44714
rect 4840 44662 4892 44714
rect 4892 44662 4896 44714
rect 4632 44660 4688 44662
rect 4736 44660 4792 44662
rect 4840 44660 4896 44662
rect 4944 44660 5000 44716
rect 5048 44714 5104 44716
rect 5152 44714 5208 44716
rect 5048 44662 5068 44714
rect 5068 44662 5104 44714
rect 5152 44662 5192 44714
rect 5192 44662 5208 44714
rect 5048 44660 5104 44662
rect 5152 44660 5208 44662
rect 4008 43146 4064 43148
rect 4112 43146 4168 43148
rect 4008 43094 4024 43146
rect 4024 43094 4064 43146
rect 4112 43094 4148 43146
rect 4148 43094 4168 43146
rect 4008 43092 4064 43094
rect 4112 43092 4168 43094
rect 4216 43092 4272 43148
rect 4320 43146 4376 43148
rect 4424 43146 4480 43148
rect 4528 43146 4584 43148
rect 4320 43094 4324 43146
rect 4324 43094 4376 43146
rect 4424 43094 4448 43146
rect 4448 43094 4480 43146
rect 4528 43094 4572 43146
rect 4572 43094 4584 43146
rect 4320 43092 4376 43094
rect 4424 43092 4480 43094
rect 4528 43092 4584 43094
rect 4632 43146 4688 43148
rect 4736 43146 4792 43148
rect 4840 43146 4896 43148
rect 4632 43094 4644 43146
rect 4644 43094 4688 43146
rect 4736 43094 4768 43146
rect 4768 43094 4792 43146
rect 4840 43094 4892 43146
rect 4892 43094 4896 43146
rect 4632 43092 4688 43094
rect 4736 43092 4792 43094
rect 4840 43092 4896 43094
rect 4944 43092 5000 43148
rect 5048 43146 5104 43148
rect 5152 43146 5208 43148
rect 5048 43094 5068 43146
rect 5068 43094 5104 43146
rect 5152 43094 5192 43146
rect 5192 43094 5208 43146
rect 5048 43092 5104 43094
rect 5152 43092 5208 43094
rect 4008 41578 4064 41580
rect 4112 41578 4168 41580
rect 4008 41526 4024 41578
rect 4024 41526 4064 41578
rect 4112 41526 4148 41578
rect 4148 41526 4168 41578
rect 4008 41524 4064 41526
rect 4112 41524 4168 41526
rect 4216 41524 4272 41580
rect 4320 41578 4376 41580
rect 4424 41578 4480 41580
rect 4528 41578 4584 41580
rect 4320 41526 4324 41578
rect 4324 41526 4376 41578
rect 4424 41526 4448 41578
rect 4448 41526 4480 41578
rect 4528 41526 4572 41578
rect 4572 41526 4584 41578
rect 4320 41524 4376 41526
rect 4424 41524 4480 41526
rect 4528 41524 4584 41526
rect 4632 41578 4688 41580
rect 4736 41578 4792 41580
rect 4840 41578 4896 41580
rect 4632 41526 4644 41578
rect 4644 41526 4688 41578
rect 4736 41526 4768 41578
rect 4768 41526 4792 41578
rect 4840 41526 4892 41578
rect 4892 41526 4896 41578
rect 4632 41524 4688 41526
rect 4736 41524 4792 41526
rect 4840 41524 4896 41526
rect 4944 41524 5000 41580
rect 5048 41578 5104 41580
rect 5152 41578 5208 41580
rect 5048 41526 5068 41578
rect 5068 41526 5104 41578
rect 5152 41526 5192 41578
rect 5192 41526 5208 41578
rect 5048 41524 5104 41526
rect 5152 41524 5208 41526
rect 4008 40010 4064 40012
rect 4112 40010 4168 40012
rect 4008 39958 4024 40010
rect 4024 39958 4064 40010
rect 4112 39958 4148 40010
rect 4148 39958 4168 40010
rect 4008 39956 4064 39958
rect 4112 39956 4168 39958
rect 4216 39956 4272 40012
rect 4320 40010 4376 40012
rect 4424 40010 4480 40012
rect 4528 40010 4584 40012
rect 4320 39958 4324 40010
rect 4324 39958 4376 40010
rect 4424 39958 4448 40010
rect 4448 39958 4480 40010
rect 4528 39958 4572 40010
rect 4572 39958 4584 40010
rect 4320 39956 4376 39958
rect 4424 39956 4480 39958
rect 4528 39956 4584 39958
rect 4632 40010 4688 40012
rect 4736 40010 4792 40012
rect 4840 40010 4896 40012
rect 4632 39958 4644 40010
rect 4644 39958 4688 40010
rect 4736 39958 4768 40010
rect 4768 39958 4792 40010
rect 4840 39958 4892 40010
rect 4892 39958 4896 40010
rect 4632 39956 4688 39958
rect 4736 39956 4792 39958
rect 4840 39956 4896 39958
rect 4944 39956 5000 40012
rect 5048 40010 5104 40012
rect 5152 40010 5208 40012
rect 5048 39958 5068 40010
rect 5068 39958 5104 40010
rect 5152 39958 5192 40010
rect 5192 39958 5208 40010
rect 5048 39956 5104 39958
rect 5152 39956 5208 39958
rect 4008 38442 4064 38444
rect 4112 38442 4168 38444
rect 4008 38390 4024 38442
rect 4024 38390 4064 38442
rect 4112 38390 4148 38442
rect 4148 38390 4168 38442
rect 4008 38388 4064 38390
rect 4112 38388 4168 38390
rect 4216 38388 4272 38444
rect 4320 38442 4376 38444
rect 4424 38442 4480 38444
rect 4528 38442 4584 38444
rect 4320 38390 4324 38442
rect 4324 38390 4376 38442
rect 4424 38390 4448 38442
rect 4448 38390 4480 38442
rect 4528 38390 4572 38442
rect 4572 38390 4584 38442
rect 4320 38388 4376 38390
rect 4424 38388 4480 38390
rect 4528 38388 4584 38390
rect 4632 38442 4688 38444
rect 4736 38442 4792 38444
rect 4840 38442 4896 38444
rect 4632 38390 4644 38442
rect 4644 38390 4688 38442
rect 4736 38390 4768 38442
rect 4768 38390 4792 38442
rect 4840 38390 4892 38442
rect 4892 38390 4896 38442
rect 4632 38388 4688 38390
rect 4736 38388 4792 38390
rect 4840 38388 4896 38390
rect 4944 38388 5000 38444
rect 5048 38442 5104 38444
rect 5152 38442 5208 38444
rect 5048 38390 5068 38442
rect 5068 38390 5104 38442
rect 5152 38390 5192 38442
rect 5192 38390 5208 38442
rect 5048 38388 5104 38390
rect 5152 38388 5208 38390
rect 4008 36874 4064 36876
rect 4112 36874 4168 36876
rect 4008 36822 4024 36874
rect 4024 36822 4064 36874
rect 4112 36822 4148 36874
rect 4148 36822 4168 36874
rect 4008 36820 4064 36822
rect 4112 36820 4168 36822
rect 4216 36820 4272 36876
rect 4320 36874 4376 36876
rect 4424 36874 4480 36876
rect 4528 36874 4584 36876
rect 4320 36822 4324 36874
rect 4324 36822 4376 36874
rect 4424 36822 4448 36874
rect 4448 36822 4480 36874
rect 4528 36822 4572 36874
rect 4572 36822 4584 36874
rect 4320 36820 4376 36822
rect 4424 36820 4480 36822
rect 4528 36820 4584 36822
rect 4632 36874 4688 36876
rect 4736 36874 4792 36876
rect 4840 36874 4896 36876
rect 4632 36822 4644 36874
rect 4644 36822 4688 36874
rect 4736 36822 4768 36874
rect 4768 36822 4792 36874
rect 4840 36822 4892 36874
rect 4892 36822 4896 36874
rect 4632 36820 4688 36822
rect 4736 36820 4792 36822
rect 4840 36820 4896 36822
rect 4944 36820 5000 36876
rect 5048 36874 5104 36876
rect 5152 36874 5208 36876
rect 5048 36822 5068 36874
rect 5068 36822 5104 36874
rect 5152 36822 5192 36874
rect 5192 36822 5208 36874
rect 5048 36820 5104 36822
rect 5152 36820 5208 36822
rect 4008 35306 4064 35308
rect 4112 35306 4168 35308
rect 4008 35254 4024 35306
rect 4024 35254 4064 35306
rect 4112 35254 4148 35306
rect 4148 35254 4168 35306
rect 4008 35252 4064 35254
rect 4112 35252 4168 35254
rect 4216 35252 4272 35308
rect 4320 35306 4376 35308
rect 4424 35306 4480 35308
rect 4528 35306 4584 35308
rect 4320 35254 4324 35306
rect 4324 35254 4376 35306
rect 4424 35254 4448 35306
rect 4448 35254 4480 35306
rect 4528 35254 4572 35306
rect 4572 35254 4584 35306
rect 4320 35252 4376 35254
rect 4424 35252 4480 35254
rect 4528 35252 4584 35254
rect 4632 35306 4688 35308
rect 4736 35306 4792 35308
rect 4840 35306 4896 35308
rect 4632 35254 4644 35306
rect 4644 35254 4688 35306
rect 4736 35254 4768 35306
rect 4768 35254 4792 35306
rect 4840 35254 4892 35306
rect 4892 35254 4896 35306
rect 4632 35252 4688 35254
rect 4736 35252 4792 35254
rect 4840 35252 4896 35254
rect 4944 35252 5000 35308
rect 5048 35306 5104 35308
rect 5152 35306 5208 35308
rect 5048 35254 5068 35306
rect 5068 35254 5104 35306
rect 5152 35254 5192 35306
rect 5192 35254 5208 35306
rect 5048 35252 5104 35254
rect 5152 35252 5208 35254
rect 4008 33738 4064 33740
rect 4112 33738 4168 33740
rect 4008 33686 4024 33738
rect 4024 33686 4064 33738
rect 4112 33686 4148 33738
rect 4148 33686 4168 33738
rect 4008 33684 4064 33686
rect 4112 33684 4168 33686
rect 4216 33684 4272 33740
rect 4320 33738 4376 33740
rect 4424 33738 4480 33740
rect 4528 33738 4584 33740
rect 4320 33686 4324 33738
rect 4324 33686 4376 33738
rect 4424 33686 4448 33738
rect 4448 33686 4480 33738
rect 4528 33686 4572 33738
rect 4572 33686 4584 33738
rect 4320 33684 4376 33686
rect 4424 33684 4480 33686
rect 4528 33684 4584 33686
rect 4632 33738 4688 33740
rect 4736 33738 4792 33740
rect 4840 33738 4896 33740
rect 4632 33686 4644 33738
rect 4644 33686 4688 33738
rect 4736 33686 4768 33738
rect 4768 33686 4792 33738
rect 4840 33686 4892 33738
rect 4892 33686 4896 33738
rect 4632 33684 4688 33686
rect 4736 33684 4792 33686
rect 4840 33684 4896 33686
rect 4944 33684 5000 33740
rect 5048 33738 5104 33740
rect 5152 33738 5208 33740
rect 5048 33686 5068 33738
rect 5068 33686 5104 33738
rect 5152 33686 5192 33738
rect 5192 33686 5208 33738
rect 5048 33684 5104 33686
rect 5152 33684 5208 33686
rect 4008 32170 4064 32172
rect 4112 32170 4168 32172
rect 4008 32118 4024 32170
rect 4024 32118 4064 32170
rect 4112 32118 4148 32170
rect 4148 32118 4168 32170
rect 4008 32116 4064 32118
rect 4112 32116 4168 32118
rect 4216 32116 4272 32172
rect 4320 32170 4376 32172
rect 4424 32170 4480 32172
rect 4528 32170 4584 32172
rect 4320 32118 4324 32170
rect 4324 32118 4376 32170
rect 4424 32118 4448 32170
rect 4448 32118 4480 32170
rect 4528 32118 4572 32170
rect 4572 32118 4584 32170
rect 4320 32116 4376 32118
rect 4424 32116 4480 32118
rect 4528 32116 4584 32118
rect 4632 32170 4688 32172
rect 4736 32170 4792 32172
rect 4840 32170 4896 32172
rect 4632 32118 4644 32170
rect 4644 32118 4688 32170
rect 4736 32118 4768 32170
rect 4768 32118 4792 32170
rect 4840 32118 4892 32170
rect 4892 32118 4896 32170
rect 4632 32116 4688 32118
rect 4736 32116 4792 32118
rect 4840 32116 4896 32118
rect 4944 32116 5000 32172
rect 5048 32170 5104 32172
rect 5152 32170 5208 32172
rect 5048 32118 5068 32170
rect 5068 32118 5104 32170
rect 5152 32118 5192 32170
rect 5192 32118 5208 32170
rect 5048 32116 5104 32118
rect 5152 32116 5208 32118
rect 4008 30602 4064 30604
rect 4112 30602 4168 30604
rect 4008 30550 4024 30602
rect 4024 30550 4064 30602
rect 4112 30550 4148 30602
rect 4148 30550 4168 30602
rect 4008 30548 4064 30550
rect 4112 30548 4168 30550
rect 4216 30548 4272 30604
rect 4320 30602 4376 30604
rect 4424 30602 4480 30604
rect 4528 30602 4584 30604
rect 4320 30550 4324 30602
rect 4324 30550 4376 30602
rect 4424 30550 4448 30602
rect 4448 30550 4480 30602
rect 4528 30550 4572 30602
rect 4572 30550 4584 30602
rect 4320 30548 4376 30550
rect 4424 30548 4480 30550
rect 4528 30548 4584 30550
rect 4632 30602 4688 30604
rect 4736 30602 4792 30604
rect 4840 30602 4896 30604
rect 4632 30550 4644 30602
rect 4644 30550 4688 30602
rect 4736 30550 4768 30602
rect 4768 30550 4792 30602
rect 4840 30550 4892 30602
rect 4892 30550 4896 30602
rect 4632 30548 4688 30550
rect 4736 30548 4792 30550
rect 4840 30548 4896 30550
rect 4944 30548 5000 30604
rect 5048 30602 5104 30604
rect 5152 30602 5208 30604
rect 5048 30550 5068 30602
rect 5068 30550 5104 30602
rect 5152 30550 5192 30602
rect 5192 30550 5208 30602
rect 5048 30548 5104 30550
rect 5152 30548 5208 30550
rect 4008 29034 4064 29036
rect 4112 29034 4168 29036
rect 4008 28982 4024 29034
rect 4024 28982 4064 29034
rect 4112 28982 4148 29034
rect 4148 28982 4168 29034
rect 4008 28980 4064 28982
rect 4112 28980 4168 28982
rect 4216 28980 4272 29036
rect 4320 29034 4376 29036
rect 4424 29034 4480 29036
rect 4528 29034 4584 29036
rect 4320 28982 4324 29034
rect 4324 28982 4376 29034
rect 4424 28982 4448 29034
rect 4448 28982 4480 29034
rect 4528 28982 4572 29034
rect 4572 28982 4584 29034
rect 4320 28980 4376 28982
rect 4424 28980 4480 28982
rect 4528 28980 4584 28982
rect 4632 29034 4688 29036
rect 4736 29034 4792 29036
rect 4840 29034 4896 29036
rect 4632 28982 4644 29034
rect 4644 28982 4688 29034
rect 4736 28982 4768 29034
rect 4768 28982 4792 29034
rect 4840 28982 4892 29034
rect 4892 28982 4896 29034
rect 4632 28980 4688 28982
rect 4736 28980 4792 28982
rect 4840 28980 4896 28982
rect 4944 28980 5000 29036
rect 5048 29034 5104 29036
rect 5152 29034 5208 29036
rect 5048 28982 5068 29034
rect 5068 28982 5104 29034
rect 5152 28982 5192 29034
rect 5192 28982 5208 29034
rect 5048 28980 5104 28982
rect 5152 28980 5208 28982
rect 4008 27466 4064 27468
rect 4112 27466 4168 27468
rect 4008 27414 4024 27466
rect 4024 27414 4064 27466
rect 4112 27414 4148 27466
rect 4148 27414 4168 27466
rect 4008 27412 4064 27414
rect 4112 27412 4168 27414
rect 4216 27412 4272 27468
rect 4320 27466 4376 27468
rect 4424 27466 4480 27468
rect 4528 27466 4584 27468
rect 4320 27414 4324 27466
rect 4324 27414 4376 27466
rect 4424 27414 4448 27466
rect 4448 27414 4480 27466
rect 4528 27414 4572 27466
rect 4572 27414 4584 27466
rect 4320 27412 4376 27414
rect 4424 27412 4480 27414
rect 4528 27412 4584 27414
rect 4632 27466 4688 27468
rect 4736 27466 4792 27468
rect 4840 27466 4896 27468
rect 4632 27414 4644 27466
rect 4644 27414 4688 27466
rect 4736 27414 4768 27466
rect 4768 27414 4792 27466
rect 4840 27414 4892 27466
rect 4892 27414 4896 27466
rect 4632 27412 4688 27414
rect 4736 27412 4792 27414
rect 4840 27412 4896 27414
rect 4944 27412 5000 27468
rect 5048 27466 5104 27468
rect 5152 27466 5208 27468
rect 5048 27414 5068 27466
rect 5068 27414 5104 27466
rect 5152 27414 5192 27466
rect 5192 27414 5208 27466
rect 5048 27412 5104 27414
rect 5152 27412 5208 27414
rect 4008 25898 4064 25900
rect 4112 25898 4168 25900
rect 4008 25846 4024 25898
rect 4024 25846 4064 25898
rect 4112 25846 4148 25898
rect 4148 25846 4168 25898
rect 4008 25844 4064 25846
rect 4112 25844 4168 25846
rect 4216 25844 4272 25900
rect 4320 25898 4376 25900
rect 4424 25898 4480 25900
rect 4528 25898 4584 25900
rect 4320 25846 4324 25898
rect 4324 25846 4376 25898
rect 4424 25846 4448 25898
rect 4448 25846 4480 25898
rect 4528 25846 4572 25898
rect 4572 25846 4584 25898
rect 4320 25844 4376 25846
rect 4424 25844 4480 25846
rect 4528 25844 4584 25846
rect 4632 25898 4688 25900
rect 4736 25898 4792 25900
rect 4840 25898 4896 25900
rect 4632 25846 4644 25898
rect 4644 25846 4688 25898
rect 4736 25846 4768 25898
rect 4768 25846 4792 25898
rect 4840 25846 4892 25898
rect 4892 25846 4896 25898
rect 4632 25844 4688 25846
rect 4736 25844 4792 25846
rect 4840 25844 4896 25846
rect 4944 25844 5000 25900
rect 5048 25898 5104 25900
rect 5152 25898 5208 25900
rect 5048 25846 5068 25898
rect 5068 25846 5104 25898
rect 5152 25846 5192 25898
rect 5192 25846 5208 25898
rect 5048 25844 5104 25846
rect 5152 25844 5208 25846
rect 4008 24330 4064 24332
rect 4112 24330 4168 24332
rect 4008 24278 4024 24330
rect 4024 24278 4064 24330
rect 4112 24278 4148 24330
rect 4148 24278 4168 24330
rect 4008 24276 4064 24278
rect 4112 24276 4168 24278
rect 4216 24276 4272 24332
rect 4320 24330 4376 24332
rect 4424 24330 4480 24332
rect 4528 24330 4584 24332
rect 4320 24278 4324 24330
rect 4324 24278 4376 24330
rect 4424 24278 4448 24330
rect 4448 24278 4480 24330
rect 4528 24278 4572 24330
rect 4572 24278 4584 24330
rect 4320 24276 4376 24278
rect 4424 24276 4480 24278
rect 4528 24276 4584 24278
rect 4632 24330 4688 24332
rect 4736 24330 4792 24332
rect 4840 24330 4896 24332
rect 4632 24278 4644 24330
rect 4644 24278 4688 24330
rect 4736 24278 4768 24330
rect 4768 24278 4792 24330
rect 4840 24278 4892 24330
rect 4892 24278 4896 24330
rect 4632 24276 4688 24278
rect 4736 24276 4792 24278
rect 4840 24276 4896 24278
rect 4944 24276 5000 24332
rect 5048 24330 5104 24332
rect 5152 24330 5208 24332
rect 5048 24278 5068 24330
rect 5068 24278 5104 24330
rect 5152 24278 5192 24330
rect 5192 24278 5208 24330
rect 5048 24276 5104 24278
rect 5152 24276 5208 24278
rect 4008 22762 4064 22764
rect 4112 22762 4168 22764
rect 4008 22710 4024 22762
rect 4024 22710 4064 22762
rect 4112 22710 4148 22762
rect 4148 22710 4168 22762
rect 4008 22708 4064 22710
rect 4112 22708 4168 22710
rect 4216 22708 4272 22764
rect 4320 22762 4376 22764
rect 4424 22762 4480 22764
rect 4528 22762 4584 22764
rect 4320 22710 4324 22762
rect 4324 22710 4376 22762
rect 4424 22710 4448 22762
rect 4448 22710 4480 22762
rect 4528 22710 4572 22762
rect 4572 22710 4584 22762
rect 4320 22708 4376 22710
rect 4424 22708 4480 22710
rect 4528 22708 4584 22710
rect 4632 22762 4688 22764
rect 4736 22762 4792 22764
rect 4840 22762 4896 22764
rect 4632 22710 4644 22762
rect 4644 22710 4688 22762
rect 4736 22710 4768 22762
rect 4768 22710 4792 22762
rect 4840 22710 4892 22762
rect 4892 22710 4896 22762
rect 4632 22708 4688 22710
rect 4736 22708 4792 22710
rect 4840 22708 4896 22710
rect 4944 22708 5000 22764
rect 5048 22762 5104 22764
rect 5152 22762 5208 22764
rect 5048 22710 5068 22762
rect 5068 22710 5104 22762
rect 5152 22710 5192 22762
rect 5192 22710 5208 22762
rect 5048 22708 5104 22710
rect 5152 22708 5208 22710
rect 4008 21194 4064 21196
rect 4112 21194 4168 21196
rect 4008 21142 4024 21194
rect 4024 21142 4064 21194
rect 4112 21142 4148 21194
rect 4148 21142 4168 21194
rect 4008 21140 4064 21142
rect 4112 21140 4168 21142
rect 4216 21140 4272 21196
rect 4320 21194 4376 21196
rect 4424 21194 4480 21196
rect 4528 21194 4584 21196
rect 4320 21142 4324 21194
rect 4324 21142 4376 21194
rect 4424 21142 4448 21194
rect 4448 21142 4480 21194
rect 4528 21142 4572 21194
rect 4572 21142 4584 21194
rect 4320 21140 4376 21142
rect 4424 21140 4480 21142
rect 4528 21140 4584 21142
rect 4632 21194 4688 21196
rect 4736 21194 4792 21196
rect 4840 21194 4896 21196
rect 4632 21142 4644 21194
rect 4644 21142 4688 21194
rect 4736 21142 4768 21194
rect 4768 21142 4792 21194
rect 4840 21142 4892 21194
rect 4892 21142 4896 21194
rect 4632 21140 4688 21142
rect 4736 21140 4792 21142
rect 4840 21140 4896 21142
rect 4944 21140 5000 21196
rect 5048 21194 5104 21196
rect 5152 21194 5208 21196
rect 5048 21142 5068 21194
rect 5068 21142 5104 21194
rect 5152 21142 5192 21194
rect 5192 21142 5208 21194
rect 5048 21140 5104 21142
rect 5152 21140 5208 21142
rect 4008 19626 4064 19628
rect 4112 19626 4168 19628
rect 4008 19574 4024 19626
rect 4024 19574 4064 19626
rect 4112 19574 4148 19626
rect 4148 19574 4168 19626
rect 4008 19572 4064 19574
rect 4112 19572 4168 19574
rect 4216 19572 4272 19628
rect 4320 19626 4376 19628
rect 4424 19626 4480 19628
rect 4528 19626 4584 19628
rect 4320 19574 4324 19626
rect 4324 19574 4376 19626
rect 4424 19574 4448 19626
rect 4448 19574 4480 19626
rect 4528 19574 4572 19626
rect 4572 19574 4584 19626
rect 4320 19572 4376 19574
rect 4424 19572 4480 19574
rect 4528 19572 4584 19574
rect 4632 19626 4688 19628
rect 4736 19626 4792 19628
rect 4840 19626 4896 19628
rect 4632 19574 4644 19626
rect 4644 19574 4688 19626
rect 4736 19574 4768 19626
rect 4768 19574 4792 19626
rect 4840 19574 4892 19626
rect 4892 19574 4896 19626
rect 4632 19572 4688 19574
rect 4736 19572 4792 19574
rect 4840 19572 4896 19574
rect 4944 19572 5000 19628
rect 5048 19626 5104 19628
rect 5152 19626 5208 19628
rect 5048 19574 5068 19626
rect 5068 19574 5104 19626
rect 5152 19574 5192 19626
rect 5192 19574 5208 19626
rect 5048 19572 5104 19574
rect 5152 19572 5208 19574
rect 4008 18058 4064 18060
rect 4112 18058 4168 18060
rect 4008 18006 4024 18058
rect 4024 18006 4064 18058
rect 4112 18006 4148 18058
rect 4148 18006 4168 18058
rect 4008 18004 4064 18006
rect 4112 18004 4168 18006
rect 4216 18004 4272 18060
rect 4320 18058 4376 18060
rect 4424 18058 4480 18060
rect 4528 18058 4584 18060
rect 4320 18006 4324 18058
rect 4324 18006 4376 18058
rect 4424 18006 4448 18058
rect 4448 18006 4480 18058
rect 4528 18006 4572 18058
rect 4572 18006 4584 18058
rect 4320 18004 4376 18006
rect 4424 18004 4480 18006
rect 4528 18004 4584 18006
rect 4632 18058 4688 18060
rect 4736 18058 4792 18060
rect 4840 18058 4896 18060
rect 4632 18006 4644 18058
rect 4644 18006 4688 18058
rect 4736 18006 4768 18058
rect 4768 18006 4792 18058
rect 4840 18006 4892 18058
rect 4892 18006 4896 18058
rect 4632 18004 4688 18006
rect 4736 18004 4792 18006
rect 4840 18004 4896 18006
rect 4944 18004 5000 18060
rect 5048 18058 5104 18060
rect 5152 18058 5208 18060
rect 5048 18006 5068 18058
rect 5068 18006 5104 18058
rect 5152 18006 5192 18058
rect 5192 18006 5208 18058
rect 5048 18004 5104 18006
rect 5152 18004 5208 18006
rect 4008 16490 4064 16492
rect 4112 16490 4168 16492
rect 4008 16438 4024 16490
rect 4024 16438 4064 16490
rect 4112 16438 4148 16490
rect 4148 16438 4168 16490
rect 4008 16436 4064 16438
rect 4112 16436 4168 16438
rect 4216 16436 4272 16492
rect 4320 16490 4376 16492
rect 4424 16490 4480 16492
rect 4528 16490 4584 16492
rect 4320 16438 4324 16490
rect 4324 16438 4376 16490
rect 4424 16438 4448 16490
rect 4448 16438 4480 16490
rect 4528 16438 4572 16490
rect 4572 16438 4584 16490
rect 4320 16436 4376 16438
rect 4424 16436 4480 16438
rect 4528 16436 4584 16438
rect 4632 16490 4688 16492
rect 4736 16490 4792 16492
rect 4840 16490 4896 16492
rect 4632 16438 4644 16490
rect 4644 16438 4688 16490
rect 4736 16438 4768 16490
rect 4768 16438 4792 16490
rect 4840 16438 4892 16490
rect 4892 16438 4896 16490
rect 4632 16436 4688 16438
rect 4736 16436 4792 16438
rect 4840 16436 4896 16438
rect 4944 16436 5000 16492
rect 5048 16490 5104 16492
rect 5152 16490 5208 16492
rect 5048 16438 5068 16490
rect 5068 16438 5104 16490
rect 5152 16438 5192 16490
rect 5192 16438 5208 16490
rect 5048 16436 5104 16438
rect 5152 16436 5208 16438
rect 4008 14922 4064 14924
rect 4112 14922 4168 14924
rect 4008 14870 4024 14922
rect 4024 14870 4064 14922
rect 4112 14870 4148 14922
rect 4148 14870 4168 14922
rect 4008 14868 4064 14870
rect 4112 14868 4168 14870
rect 4216 14868 4272 14924
rect 4320 14922 4376 14924
rect 4424 14922 4480 14924
rect 4528 14922 4584 14924
rect 4320 14870 4324 14922
rect 4324 14870 4376 14922
rect 4424 14870 4448 14922
rect 4448 14870 4480 14922
rect 4528 14870 4572 14922
rect 4572 14870 4584 14922
rect 4320 14868 4376 14870
rect 4424 14868 4480 14870
rect 4528 14868 4584 14870
rect 4632 14922 4688 14924
rect 4736 14922 4792 14924
rect 4840 14922 4896 14924
rect 4632 14870 4644 14922
rect 4644 14870 4688 14922
rect 4736 14870 4768 14922
rect 4768 14870 4792 14922
rect 4840 14870 4892 14922
rect 4892 14870 4896 14922
rect 4632 14868 4688 14870
rect 4736 14868 4792 14870
rect 4840 14868 4896 14870
rect 4944 14868 5000 14924
rect 5048 14922 5104 14924
rect 5152 14922 5208 14924
rect 5048 14870 5068 14922
rect 5068 14870 5104 14922
rect 5152 14870 5192 14922
rect 5192 14870 5208 14922
rect 5048 14868 5104 14870
rect 5152 14868 5208 14870
rect 4008 13354 4064 13356
rect 4112 13354 4168 13356
rect 4008 13302 4024 13354
rect 4024 13302 4064 13354
rect 4112 13302 4148 13354
rect 4148 13302 4168 13354
rect 4008 13300 4064 13302
rect 4112 13300 4168 13302
rect 4216 13300 4272 13356
rect 4320 13354 4376 13356
rect 4424 13354 4480 13356
rect 4528 13354 4584 13356
rect 4320 13302 4324 13354
rect 4324 13302 4376 13354
rect 4424 13302 4448 13354
rect 4448 13302 4480 13354
rect 4528 13302 4572 13354
rect 4572 13302 4584 13354
rect 4320 13300 4376 13302
rect 4424 13300 4480 13302
rect 4528 13300 4584 13302
rect 4632 13354 4688 13356
rect 4736 13354 4792 13356
rect 4840 13354 4896 13356
rect 4632 13302 4644 13354
rect 4644 13302 4688 13354
rect 4736 13302 4768 13354
rect 4768 13302 4792 13354
rect 4840 13302 4892 13354
rect 4892 13302 4896 13354
rect 4632 13300 4688 13302
rect 4736 13300 4792 13302
rect 4840 13300 4896 13302
rect 4944 13300 5000 13356
rect 5048 13354 5104 13356
rect 5152 13354 5208 13356
rect 5048 13302 5068 13354
rect 5068 13302 5104 13354
rect 5152 13302 5192 13354
rect 5192 13302 5208 13354
rect 5048 13300 5104 13302
rect 5152 13300 5208 13302
rect 4008 11786 4064 11788
rect 4112 11786 4168 11788
rect 4008 11734 4024 11786
rect 4024 11734 4064 11786
rect 4112 11734 4148 11786
rect 4148 11734 4168 11786
rect 4008 11732 4064 11734
rect 4112 11732 4168 11734
rect 4216 11732 4272 11788
rect 4320 11786 4376 11788
rect 4424 11786 4480 11788
rect 4528 11786 4584 11788
rect 4320 11734 4324 11786
rect 4324 11734 4376 11786
rect 4424 11734 4448 11786
rect 4448 11734 4480 11786
rect 4528 11734 4572 11786
rect 4572 11734 4584 11786
rect 4320 11732 4376 11734
rect 4424 11732 4480 11734
rect 4528 11732 4584 11734
rect 4632 11786 4688 11788
rect 4736 11786 4792 11788
rect 4840 11786 4896 11788
rect 4632 11734 4644 11786
rect 4644 11734 4688 11786
rect 4736 11734 4768 11786
rect 4768 11734 4792 11786
rect 4840 11734 4892 11786
rect 4892 11734 4896 11786
rect 4632 11732 4688 11734
rect 4736 11732 4792 11734
rect 4840 11732 4896 11734
rect 4944 11732 5000 11788
rect 5048 11786 5104 11788
rect 5152 11786 5208 11788
rect 5048 11734 5068 11786
rect 5068 11734 5104 11786
rect 5152 11734 5192 11786
rect 5192 11734 5208 11786
rect 5048 11732 5104 11734
rect 5152 11732 5208 11734
rect 10332 10556 10388 10612
rect 4008 10218 4064 10220
rect 4112 10218 4168 10220
rect 4008 10166 4024 10218
rect 4024 10166 4064 10218
rect 4112 10166 4148 10218
rect 4148 10166 4168 10218
rect 4008 10164 4064 10166
rect 4112 10164 4168 10166
rect 4216 10164 4272 10220
rect 4320 10218 4376 10220
rect 4424 10218 4480 10220
rect 4528 10218 4584 10220
rect 4320 10166 4324 10218
rect 4324 10166 4376 10218
rect 4424 10166 4448 10218
rect 4448 10166 4480 10218
rect 4528 10166 4572 10218
rect 4572 10166 4584 10218
rect 4320 10164 4376 10166
rect 4424 10164 4480 10166
rect 4528 10164 4584 10166
rect 4632 10218 4688 10220
rect 4736 10218 4792 10220
rect 4840 10218 4896 10220
rect 4632 10166 4644 10218
rect 4644 10166 4688 10218
rect 4736 10166 4768 10218
rect 4768 10166 4792 10218
rect 4840 10166 4892 10218
rect 4892 10166 4896 10218
rect 4632 10164 4688 10166
rect 4736 10164 4792 10166
rect 4840 10164 4896 10166
rect 4944 10164 5000 10220
rect 5048 10218 5104 10220
rect 5152 10218 5208 10220
rect 5048 10166 5068 10218
rect 5068 10166 5104 10218
rect 5152 10166 5192 10218
rect 5192 10166 5208 10218
rect 5048 10164 5104 10166
rect 5152 10164 5208 10166
rect 7756 9714 7812 9716
rect 7756 9662 7758 9714
rect 7758 9662 7810 9714
rect 7810 9662 7812 9714
rect 7756 9660 7812 9662
rect 8316 9714 8372 9716
rect 8316 9662 8318 9714
rect 8318 9662 8370 9714
rect 8370 9662 8372 9714
rect 8316 9660 8372 9662
rect 4008 8650 4064 8652
rect 4112 8650 4168 8652
rect 4008 8598 4024 8650
rect 4024 8598 4064 8650
rect 4112 8598 4148 8650
rect 4148 8598 4168 8650
rect 4008 8596 4064 8598
rect 4112 8596 4168 8598
rect 4216 8596 4272 8652
rect 4320 8650 4376 8652
rect 4424 8650 4480 8652
rect 4528 8650 4584 8652
rect 4320 8598 4324 8650
rect 4324 8598 4376 8650
rect 4424 8598 4448 8650
rect 4448 8598 4480 8650
rect 4528 8598 4572 8650
rect 4572 8598 4584 8650
rect 4320 8596 4376 8598
rect 4424 8596 4480 8598
rect 4528 8596 4584 8598
rect 4632 8650 4688 8652
rect 4736 8650 4792 8652
rect 4840 8650 4896 8652
rect 4632 8598 4644 8650
rect 4644 8598 4688 8650
rect 4736 8598 4768 8650
rect 4768 8598 4792 8650
rect 4840 8598 4892 8650
rect 4892 8598 4896 8650
rect 4632 8596 4688 8598
rect 4736 8596 4792 8598
rect 4840 8596 4896 8598
rect 4944 8596 5000 8652
rect 5048 8650 5104 8652
rect 5152 8650 5208 8652
rect 5048 8598 5068 8650
rect 5068 8598 5104 8650
rect 5152 8598 5192 8650
rect 5192 8598 5208 8650
rect 5048 8596 5104 8598
rect 5152 8596 5208 8598
rect 5964 8258 6020 8260
rect 5964 8206 5966 8258
rect 5966 8206 6018 8258
rect 6018 8206 6020 8258
rect 5964 8204 6020 8206
rect 2940 7196 2996 7252
rect 1932 6748 1988 6804
rect 2268 6412 2324 6468
rect 2604 6076 2660 6132
rect 1932 5906 1988 5908
rect 1932 5854 1934 5906
rect 1934 5854 1986 5906
rect 1986 5854 1988 5906
rect 1932 5852 1988 5854
rect 1708 4396 1764 4452
rect 2156 5346 2212 5348
rect 2156 5294 2158 5346
rect 2158 5294 2210 5346
rect 2210 5294 2212 5346
rect 2156 5292 2212 5294
rect 2044 4396 2100 4452
rect 2492 5068 2548 5124
rect 2156 2716 2212 2772
rect 3052 5068 3108 5124
rect 3500 6300 3556 6356
rect 3052 4060 3108 4116
rect 3724 5292 3780 5348
rect 4284 7196 4340 7252
rect 4008 7082 4064 7084
rect 4112 7082 4168 7084
rect 4008 7030 4024 7082
rect 4024 7030 4064 7082
rect 4112 7030 4148 7082
rect 4148 7030 4168 7082
rect 4008 7028 4064 7030
rect 4112 7028 4168 7030
rect 4216 7028 4272 7084
rect 4320 7082 4376 7084
rect 4424 7082 4480 7084
rect 4528 7082 4584 7084
rect 4320 7030 4324 7082
rect 4324 7030 4376 7082
rect 4424 7030 4448 7082
rect 4448 7030 4480 7082
rect 4528 7030 4572 7082
rect 4572 7030 4584 7082
rect 4320 7028 4376 7030
rect 4424 7028 4480 7030
rect 4528 7028 4584 7030
rect 4632 7082 4688 7084
rect 4736 7082 4792 7084
rect 4840 7082 4896 7084
rect 4632 7030 4644 7082
rect 4644 7030 4688 7082
rect 4736 7030 4768 7082
rect 4768 7030 4792 7082
rect 4840 7030 4892 7082
rect 4892 7030 4896 7082
rect 4632 7028 4688 7030
rect 4736 7028 4792 7030
rect 4840 7028 4896 7030
rect 4944 7028 5000 7084
rect 5048 7082 5104 7084
rect 5152 7082 5208 7084
rect 5048 7030 5068 7082
rect 5068 7030 5104 7082
rect 5152 7030 5192 7082
rect 5192 7030 5208 7082
rect 5048 7028 5104 7030
rect 5152 7028 5208 7030
rect 3948 6300 4004 6356
rect 4732 5964 4788 6020
rect 4732 5794 4788 5796
rect 4732 5742 4734 5794
rect 4734 5742 4786 5794
rect 4786 5742 4788 5794
rect 4732 5740 4788 5742
rect 4008 5514 4064 5516
rect 4112 5514 4168 5516
rect 4008 5462 4024 5514
rect 4024 5462 4064 5514
rect 4112 5462 4148 5514
rect 4148 5462 4168 5514
rect 4008 5460 4064 5462
rect 4112 5460 4168 5462
rect 4216 5460 4272 5516
rect 4320 5514 4376 5516
rect 4424 5514 4480 5516
rect 4528 5514 4584 5516
rect 4320 5462 4324 5514
rect 4324 5462 4376 5514
rect 4424 5462 4448 5514
rect 4448 5462 4480 5514
rect 4528 5462 4572 5514
rect 4572 5462 4584 5514
rect 4320 5460 4376 5462
rect 4424 5460 4480 5462
rect 4528 5460 4584 5462
rect 4632 5514 4688 5516
rect 4736 5514 4792 5516
rect 4840 5514 4896 5516
rect 4632 5462 4644 5514
rect 4644 5462 4688 5514
rect 4736 5462 4768 5514
rect 4768 5462 4792 5514
rect 4840 5462 4892 5514
rect 4892 5462 4896 5514
rect 4632 5460 4688 5462
rect 4736 5460 4792 5462
rect 4840 5460 4896 5462
rect 4944 5460 5000 5516
rect 5048 5514 5104 5516
rect 5152 5514 5208 5516
rect 5048 5462 5068 5514
rect 5068 5462 5104 5514
rect 5152 5462 5192 5514
rect 5192 5462 5208 5514
rect 5048 5460 5104 5462
rect 5152 5460 5208 5462
rect 4620 5180 4676 5236
rect 4060 5122 4116 5124
rect 4060 5070 4062 5122
rect 4062 5070 4114 5122
rect 4114 5070 4116 5122
rect 4060 5068 4116 5070
rect 4396 5068 4452 5124
rect 3500 3612 3556 3668
rect 3612 4060 3668 4116
rect 3836 4450 3892 4452
rect 3836 4398 3838 4450
rect 3838 4398 3890 4450
rect 3890 4398 3892 4450
rect 3836 4396 3892 4398
rect 5068 4844 5124 4900
rect 4956 4620 5012 4676
rect 5964 7644 6020 7700
rect 5516 6466 5572 6468
rect 5516 6414 5518 6466
rect 5518 6414 5570 6466
rect 5570 6414 5572 6466
rect 5516 6412 5572 6414
rect 5852 6300 5908 6356
rect 4844 4060 4900 4116
rect 5404 5292 5460 5348
rect 5516 5964 5572 6020
rect 7420 8652 7476 8708
rect 7196 8540 7252 8596
rect 6524 8034 6580 8036
rect 6524 7982 6526 8034
rect 6526 7982 6578 8034
rect 6578 7982 6580 8034
rect 6524 7980 6580 7982
rect 6972 8034 7028 8036
rect 6972 7982 6974 8034
rect 6974 7982 7026 8034
rect 7026 7982 7028 8034
rect 6972 7980 7028 7982
rect 6524 7532 6580 7588
rect 6412 7362 6468 7364
rect 6412 7310 6414 7362
rect 6414 7310 6466 7362
rect 6466 7310 6468 7362
rect 6412 7308 6468 7310
rect 6300 6466 6356 6468
rect 6300 6414 6302 6466
rect 6302 6414 6354 6466
rect 6354 6414 6356 6466
rect 6300 6412 6356 6414
rect 6188 6188 6244 6244
rect 6076 5794 6132 5796
rect 6076 5742 6078 5794
rect 6078 5742 6130 5794
rect 6130 5742 6132 5794
rect 6076 5740 6132 5742
rect 5516 5180 5572 5236
rect 6188 5068 6244 5124
rect 5852 4956 5908 5012
rect 4008 3946 4064 3948
rect 4112 3946 4168 3948
rect 4008 3894 4024 3946
rect 4024 3894 4064 3946
rect 4112 3894 4148 3946
rect 4148 3894 4168 3946
rect 4008 3892 4064 3894
rect 4112 3892 4168 3894
rect 4216 3892 4272 3948
rect 4320 3946 4376 3948
rect 4424 3946 4480 3948
rect 4528 3946 4584 3948
rect 4320 3894 4324 3946
rect 4324 3894 4376 3946
rect 4424 3894 4448 3946
rect 4448 3894 4480 3946
rect 4528 3894 4572 3946
rect 4572 3894 4584 3946
rect 4320 3892 4376 3894
rect 4424 3892 4480 3894
rect 4528 3892 4584 3894
rect 4632 3946 4688 3948
rect 4736 3946 4792 3948
rect 4840 3946 4896 3948
rect 4632 3894 4644 3946
rect 4644 3894 4688 3946
rect 4736 3894 4768 3946
rect 4768 3894 4792 3946
rect 4840 3894 4892 3946
rect 4892 3894 4896 3946
rect 4632 3892 4688 3894
rect 4736 3892 4792 3894
rect 4840 3892 4896 3894
rect 4944 3892 5000 3948
rect 5048 3946 5104 3948
rect 5152 3946 5208 3948
rect 5048 3894 5068 3946
rect 5068 3894 5104 3946
rect 5152 3894 5192 3946
rect 5192 3894 5208 3946
rect 5048 3892 5104 3894
rect 5152 3892 5208 3894
rect 5404 4060 5460 4116
rect 4284 3724 4340 3780
rect 4060 3612 4116 3668
rect 3948 3554 4004 3556
rect 3948 3502 3950 3554
rect 3950 3502 4002 3554
rect 4002 3502 4004 3554
rect 3948 3500 4004 3502
rect 5180 3500 5236 3556
rect 4956 3442 5012 3444
rect 4956 3390 4958 3442
rect 4958 3390 5010 3442
rect 5010 3390 5012 3442
rect 4956 3388 5012 3390
rect 7420 8370 7476 8372
rect 7420 8318 7422 8370
rect 7422 8318 7474 8370
rect 7474 8318 7476 8370
rect 7420 8316 7476 8318
rect 7868 8652 7924 8708
rect 7756 8370 7812 8372
rect 7756 8318 7758 8370
rect 7758 8318 7810 8370
rect 7810 8318 7812 8370
rect 7756 8316 7812 8318
rect 8204 8204 8260 8260
rect 6748 6860 6804 6916
rect 7756 7474 7812 7476
rect 7756 7422 7758 7474
rect 7758 7422 7810 7474
rect 7810 7422 7812 7474
rect 7756 7420 7812 7422
rect 8316 7980 8372 8036
rect 7980 7644 8036 7700
rect 7980 7362 8036 7364
rect 7980 7310 7982 7362
rect 7982 7310 8034 7362
rect 8034 7310 8036 7362
rect 7980 7308 8036 7310
rect 6636 6412 6692 6468
rect 6860 6188 6916 6244
rect 7084 5964 7140 6020
rect 7308 6188 7364 6244
rect 6412 4956 6468 5012
rect 6300 4508 6356 4564
rect 6860 4844 6916 4900
rect 6412 4338 6468 4340
rect 6412 4286 6414 4338
rect 6414 4286 6466 4338
rect 6466 4286 6468 4338
rect 6412 4284 6468 4286
rect 5740 3554 5796 3556
rect 5740 3502 5742 3554
rect 5742 3502 5794 3554
rect 5794 3502 5796 3554
rect 5740 3500 5796 3502
rect 6076 3836 6132 3892
rect 6524 3724 6580 3780
rect 6860 4562 6916 4564
rect 6860 4510 6862 4562
rect 6862 4510 6914 4562
rect 6914 4510 6916 4562
rect 6860 4508 6916 4510
rect 7084 5682 7140 5684
rect 7084 5630 7086 5682
rect 7086 5630 7138 5682
rect 7138 5630 7140 5682
rect 7084 5628 7140 5630
rect 6860 4060 6916 4116
rect 7980 6636 8036 6692
rect 7868 6466 7924 6468
rect 7868 6414 7870 6466
rect 7870 6414 7922 6466
rect 7922 6414 7924 6466
rect 7868 6412 7924 6414
rect 8204 7474 8260 7476
rect 8204 7422 8206 7474
rect 8206 7422 8258 7474
rect 8258 7422 8260 7474
rect 8204 7420 8260 7422
rect 8316 7308 8372 7364
rect 8204 6466 8260 6468
rect 8204 6414 8206 6466
rect 8206 6414 8258 6466
rect 8258 6414 8260 6466
rect 8204 6412 8260 6414
rect 7756 6188 7812 6244
rect 7308 4620 7364 4676
rect 7644 6018 7700 6020
rect 7644 5966 7646 6018
rect 7646 5966 7698 6018
rect 7698 5966 7700 6018
rect 7644 5964 7700 5966
rect 7756 5852 7812 5908
rect 7980 4844 8036 4900
rect 8764 8204 8820 8260
rect 8876 8876 8932 8932
rect 8652 7474 8708 7476
rect 8652 7422 8654 7474
rect 8654 7422 8706 7474
rect 8706 7422 8708 7474
rect 8652 7420 8708 7422
rect 9660 8930 9716 8932
rect 9660 8878 9662 8930
rect 9662 8878 9714 8930
rect 9714 8878 9716 8930
rect 9660 8876 9716 8878
rect 11900 10610 11956 10612
rect 11900 10558 11902 10610
rect 11902 10558 11954 10610
rect 11954 10558 11956 10610
rect 11900 10556 11956 10558
rect 12124 10610 12180 10612
rect 12124 10558 12126 10610
rect 12126 10558 12178 10610
rect 12178 10558 12180 10610
rect 12124 10556 12180 10558
rect 10780 10444 10836 10500
rect 12012 10498 12068 10500
rect 12012 10446 12014 10498
rect 12014 10446 12066 10498
rect 12066 10446 12068 10498
rect 12012 10444 12068 10446
rect 12908 10610 12964 10612
rect 12908 10558 12910 10610
rect 12910 10558 12962 10610
rect 12962 10558 12964 10610
rect 12908 10556 12964 10558
rect 9772 8540 9828 8596
rect 9324 8092 9380 8148
rect 8988 7980 9044 8036
rect 8652 6578 8708 6580
rect 8652 6526 8654 6578
rect 8654 6526 8706 6578
rect 8706 6526 8708 6578
rect 8652 6524 8708 6526
rect 8988 6076 9044 6132
rect 8540 5906 8596 5908
rect 8540 5854 8542 5906
rect 8542 5854 8594 5906
rect 8594 5854 8596 5906
rect 8540 5852 8596 5854
rect 8652 5068 8708 5124
rect 8092 3948 8148 4004
rect 7868 3724 7924 3780
rect 6972 3500 7028 3556
rect 6524 924 6580 980
rect 7420 3500 7476 3556
rect 9436 6524 9492 6580
rect 8316 3724 8372 3780
rect 8428 4172 8484 4228
rect 7084 3330 7140 3332
rect 7084 3278 7086 3330
rect 7086 3278 7138 3330
rect 7138 3278 7140 3330
rect 7084 3276 7140 3278
rect 10108 7586 10164 7588
rect 10108 7534 10110 7586
rect 10110 7534 10162 7586
rect 10162 7534 10164 7586
rect 10108 7532 10164 7534
rect 9660 5292 9716 5348
rect 8876 5180 8932 5236
rect 9436 4844 9492 4900
rect 9884 4732 9940 4788
rect 9884 4060 9940 4116
rect 10444 7308 10500 7364
rect 10780 7084 10836 7140
rect 10220 6076 10276 6132
rect 9772 3554 9828 3556
rect 9772 3502 9774 3554
rect 9774 3502 9826 3554
rect 9826 3502 9828 3554
rect 9772 3500 9828 3502
rect 9884 3724 9940 3780
rect 10220 4956 10276 5012
rect 10108 3836 10164 3892
rect 10220 4620 10276 4676
rect 9996 3612 10052 3668
rect 10668 4060 10724 4116
rect 10780 6636 10836 6692
rect 10556 3612 10612 3668
rect 10892 4956 10948 5012
rect 12684 8876 12740 8932
rect 11564 8204 11620 8260
rect 11564 7420 11620 7476
rect 11676 7084 11732 7140
rect 11452 6076 11508 6132
rect 11228 5068 11284 5124
rect 11564 5852 11620 5908
rect 12908 7308 12964 7364
rect 11788 5964 11844 6020
rect 12124 6524 12180 6580
rect 12236 5292 12292 5348
rect 12460 4898 12516 4900
rect 12460 4846 12462 4898
rect 12462 4846 12514 4898
rect 12514 4846 12516 4898
rect 12460 4844 12516 4846
rect 12572 4732 12628 4788
rect 12012 4284 12068 4340
rect 12348 4172 12404 4228
rect 11228 3388 11284 3444
rect 11452 3500 11508 3556
rect 7868 924 7924 980
rect 11676 3554 11732 3556
rect 11676 3502 11678 3554
rect 11678 3502 11730 3554
rect 11730 3502 11732 3554
rect 11676 3500 11732 3502
rect 12572 3724 12628 3780
rect 13468 8540 13524 8596
rect 24008 46282 24064 46284
rect 24112 46282 24168 46284
rect 24008 46230 24024 46282
rect 24024 46230 24064 46282
rect 24112 46230 24148 46282
rect 24148 46230 24168 46282
rect 24008 46228 24064 46230
rect 24112 46228 24168 46230
rect 24216 46228 24272 46284
rect 24320 46282 24376 46284
rect 24424 46282 24480 46284
rect 24528 46282 24584 46284
rect 24320 46230 24324 46282
rect 24324 46230 24376 46282
rect 24424 46230 24448 46282
rect 24448 46230 24480 46282
rect 24528 46230 24572 46282
rect 24572 46230 24584 46282
rect 24320 46228 24376 46230
rect 24424 46228 24480 46230
rect 24528 46228 24584 46230
rect 24632 46282 24688 46284
rect 24736 46282 24792 46284
rect 24840 46282 24896 46284
rect 24632 46230 24644 46282
rect 24644 46230 24688 46282
rect 24736 46230 24768 46282
rect 24768 46230 24792 46282
rect 24840 46230 24892 46282
rect 24892 46230 24896 46282
rect 24632 46228 24688 46230
rect 24736 46228 24792 46230
rect 24840 46228 24896 46230
rect 24944 46228 25000 46284
rect 25048 46282 25104 46284
rect 25152 46282 25208 46284
rect 25048 46230 25068 46282
rect 25068 46230 25104 46282
rect 25152 46230 25192 46282
rect 25192 46230 25208 46282
rect 25048 46228 25104 46230
rect 25152 46228 25208 46230
rect 27356 46060 27412 46116
rect 28812 46060 28868 46116
rect 14008 45498 14064 45500
rect 14112 45498 14168 45500
rect 14008 45446 14024 45498
rect 14024 45446 14064 45498
rect 14112 45446 14148 45498
rect 14148 45446 14168 45498
rect 14008 45444 14064 45446
rect 14112 45444 14168 45446
rect 14216 45444 14272 45500
rect 14320 45498 14376 45500
rect 14424 45498 14480 45500
rect 14528 45498 14584 45500
rect 14320 45446 14324 45498
rect 14324 45446 14376 45498
rect 14424 45446 14448 45498
rect 14448 45446 14480 45498
rect 14528 45446 14572 45498
rect 14572 45446 14584 45498
rect 14320 45444 14376 45446
rect 14424 45444 14480 45446
rect 14528 45444 14584 45446
rect 14632 45498 14688 45500
rect 14736 45498 14792 45500
rect 14840 45498 14896 45500
rect 14632 45446 14644 45498
rect 14644 45446 14688 45498
rect 14736 45446 14768 45498
rect 14768 45446 14792 45498
rect 14840 45446 14892 45498
rect 14892 45446 14896 45498
rect 14632 45444 14688 45446
rect 14736 45444 14792 45446
rect 14840 45444 14896 45446
rect 14944 45444 15000 45500
rect 15048 45498 15104 45500
rect 15152 45498 15208 45500
rect 15048 45446 15068 45498
rect 15068 45446 15104 45498
rect 15152 45446 15192 45498
rect 15192 45446 15208 45498
rect 15048 45444 15104 45446
rect 15152 45444 15208 45446
rect 24008 44714 24064 44716
rect 24112 44714 24168 44716
rect 24008 44662 24024 44714
rect 24024 44662 24064 44714
rect 24112 44662 24148 44714
rect 24148 44662 24168 44714
rect 24008 44660 24064 44662
rect 24112 44660 24168 44662
rect 24216 44660 24272 44716
rect 24320 44714 24376 44716
rect 24424 44714 24480 44716
rect 24528 44714 24584 44716
rect 24320 44662 24324 44714
rect 24324 44662 24376 44714
rect 24424 44662 24448 44714
rect 24448 44662 24480 44714
rect 24528 44662 24572 44714
rect 24572 44662 24584 44714
rect 24320 44660 24376 44662
rect 24424 44660 24480 44662
rect 24528 44660 24584 44662
rect 24632 44714 24688 44716
rect 24736 44714 24792 44716
rect 24840 44714 24896 44716
rect 24632 44662 24644 44714
rect 24644 44662 24688 44714
rect 24736 44662 24768 44714
rect 24768 44662 24792 44714
rect 24840 44662 24892 44714
rect 24892 44662 24896 44714
rect 24632 44660 24688 44662
rect 24736 44660 24792 44662
rect 24840 44660 24896 44662
rect 24944 44660 25000 44716
rect 25048 44714 25104 44716
rect 25152 44714 25208 44716
rect 25048 44662 25068 44714
rect 25068 44662 25104 44714
rect 25152 44662 25192 44714
rect 25192 44662 25208 44714
rect 25048 44660 25104 44662
rect 25152 44660 25208 44662
rect 14008 43930 14064 43932
rect 14112 43930 14168 43932
rect 14008 43878 14024 43930
rect 14024 43878 14064 43930
rect 14112 43878 14148 43930
rect 14148 43878 14168 43930
rect 14008 43876 14064 43878
rect 14112 43876 14168 43878
rect 14216 43876 14272 43932
rect 14320 43930 14376 43932
rect 14424 43930 14480 43932
rect 14528 43930 14584 43932
rect 14320 43878 14324 43930
rect 14324 43878 14376 43930
rect 14424 43878 14448 43930
rect 14448 43878 14480 43930
rect 14528 43878 14572 43930
rect 14572 43878 14584 43930
rect 14320 43876 14376 43878
rect 14424 43876 14480 43878
rect 14528 43876 14584 43878
rect 14632 43930 14688 43932
rect 14736 43930 14792 43932
rect 14840 43930 14896 43932
rect 14632 43878 14644 43930
rect 14644 43878 14688 43930
rect 14736 43878 14768 43930
rect 14768 43878 14792 43930
rect 14840 43878 14892 43930
rect 14892 43878 14896 43930
rect 14632 43876 14688 43878
rect 14736 43876 14792 43878
rect 14840 43876 14896 43878
rect 14944 43876 15000 43932
rect 15048 43930 15104 43932
rect 15152 43930 15208 43932
rect 15048 43878 15068 43930
rect 15068 43878 15104 43930
rect 15152 43878 15192 43930
rect 15192 43878 15208 43930
rect 15048 43876 15104 43878
rect 15152 43876 15208 43878
rect 24008 43146 24064 43148
rect 24112 43146 24168 43148
rect 24008 43094 24024 43146
rect 24024 43094 24064 43146
rect 24112 43094 24148 43146
rect 24148 43094 24168 43146
rect 24008 43092 24064 43094
rect 24112 43092 24168 43094
rect 24216 43092 24272 43148
rect 24320 43146 24376 43148
rect 24424 43146 24480 43148
rect 24528 43146 24584 43148
rect 24320 43094 24324 43146
rect 24324 43094 24376 43146
rect 24424 43094 24448 43146
rect 24448 43094 24480 43146
rect 24528 43094 24572 43146
rect 24572 43094 24584 43146
rect 24320 43092 24376 43094
rect 24424 43092 24480 43094
rect 24528 43092 24584 43094
rect 24632 43146 24688 43148
rect 24736 43146 24792 43148
rect 24840 43146 24896 43148
rect 24632 43094 24644 43146
rect 24644 43094 24688 43146
rect 24736 43094 24768 43146
rect 24768 43094 24792 43146
rect 24840 43094 24892 43146
rect 24892 43094 24896 43146
rect 24632 43092 24688 43094
rect 24736 43092 24792 43094
rect 24840 43092 24896 43094
rect 24944 43092 25000 43148
rect 25048 43146 25104 43148
rect 25152 43146 25208 43148
rect 25048 43094 25068 43146
rect 25068 43094 25104 43146
rect 25152 43094 25192 43146
rect 25192 43094 25208 43146
rect 25048 43092 25104 43094
rect 25152 43092 25208 43094
rect 14008 42362 14064 42364
rect 14112 42362 14168 42364
rect 14008 42310 14024 42362
rect 14024 42310 14064 42362
rect 14112 42310 14148 42362
rect 14148 42310 14168 42362
rect 14008 42308 14064 42310
rect 14112 42308 14168 42310
rect 14216 42308 14272 42364
rect 14320 42362 14376 42364
rect 14424 42362 14480 42364
rect 14528 42362 14584 42364
rect 14320 42310 14324 42362
rect 14324 42310 14376 42362
rect 14424 42310 14448 42362
rect 14448 42310 14480 42362
rect 14528 42310 14572 42362
rect 14572 42310 14584 42362
rect 14320 42308 14376 42310
rect 14424 42308 14480 42310
rect 14528 42308 14584 42310
rect 14632 42362 14688 42364
rect 14736 42362 14792 42364
rect 14840 42362 14896 42364
rect 14632 42310 14644 42362
rect 14644 42310 14688 42362
rect 14736 42310 14768 42362
rect 14768 42310 14792 42362
rect 14840 42310 14892 42362
rect 14892 42310 14896 42362
rect 14632 42308 14688 42310
rect 14736 42308 14792 42310
rect 14840 42308 14896 42310
rect 14944 42308 15000 42364
rect 15048 42362 15104 42364
rect 15152 42362 15208 42364
rect 15048 42310 15068 42362
rect 15068 42310 15104 42362
rect 15152 42310 15192 42362
rect 15192 42310 15208 42362
rect 15048 42308 15104 42310
rect 15152 42308 15208 42310
rect 24008 41578 24064 41580
rect 24112 41578 24168 41580
rect 24008 41526 24024 41578
rect 24024 41526 24064 41578
rect 24112 41526 24148 41578
rect 24148 41526 24168 41578
rect 24008 41524 24064 41526
rect 24112 41524 24168 41526
rect 24216 41524 24272 41580
rect 24320 41578 24376 41580
rect 24424 41578 24480 41580
rect 24528 41578 24584 41580
rect 24320 41526 24324 41578
rect 24324 41526 24376 41578
rect 24424 41526 24448 41578
rect 24448 41526 24480 41578
rect 24528 41526 24572 41578
rect 24572 41526 24584 41578
rect 24320 41524 24376 41526
rect 24424 41524 24480 41526
rect 24528 41524 24584 41526
rect 24632 41578 24688 41580
rect 24736 41578 24792 41580
rect 24840 41578 24896 41580
rect 24632 41526 24644 41578
rect 24644 41526 24688 41578
rect 24736 41526 24768 41578
rect 24768 41526 24792 41578
rect 24840 41526 24892 41578
rect 24892 41526 24896 41578
rect 24632 41524 24688 41526
rect 24736 41524 24792 41526
rect 24840 41524 24896 41526
rect 24944 41524 25000 41580
rect 25048 41578 25104 41580
rect 25152 41578 25208 41580
rect 25048 41526 25068 41578
rect 25068 41526 25104 41578
rect 25152 41526 25192 41578
rect 25192 41526 25208 41578
rect 25048 41524 25104 41526
rect 25152 41524 25208 41526
rect 14008 40794 14064 40796
rect 14112 40794 14168 40796
rect 14008 40742 14024 40794
rect 14024 40742 14064 40794
rect 14112 40742 14148 40794
rect 14148 40742 14168 40794
rect 14008 40740 14064 40742
rect 14112 40740 14168 40742
rect 14216 40740 14272 40796
rect 14320 40794 14376 40796
rect 14424 40794 14480 40796
rect 14528 40794 14584 40796
rect 14320 40742 14324 40794
rect 14324 40742 14376 40794
rect 14424 40742 14448 40794
rect 14448 40742 14480 40794
rect 14528 40742 14572 40794
rect 14572 40742 14584 40794
rect 14320 40740 14376 40742
rect 14424 40740 14480 40742
rect 14528 40740 14584 40742
rect 14632 40794 14688 40796
rect 14736 40794 14792 40796
rect 14840 40794 14896 40796
rect 14632 40742 14644 40794
rect 14644 40742 14688 40794
rect 14736 40742 14768 40794
rect 14768 40742 14792 40794
rect 14840 40742 14892 40794
rect 14892 40742 14896 40794
rect 14632 40740 14688 40742
rect 14736 40740 14792 40742
rect 14840 40740 14896 40742
rect 14944 40740 15000 40796
rect 15048 40794 15104 40796
rect 15152 40794 15208 40796
rect 15048 40742 15068 40794
rect 15068 40742 15104 40794
rect 15152 40742 15192 40794
rect 15192 40742 15208 40794
rect 15048 40740 15104 40742
rect 15152 40740 15208 40742
rect 24008 40010 24064 40012
rect 24112 40010 24168 40012
rect 24008 39958 24024 40010
rect 24024 39958 24064 40010
rect 24112 39958 24148 40010
rect 24148 39958 24168 40010
rect 24008 39956 24064 39958
rect 24112 39956 24168 39958
rect 24216 39956 24272 40012
rect 24320 40010 24376 40012
rect 24424 40010 24480 40012
rect 24528 40010 24584 40012
rect 24320 39958 24324 40010
rect 24324 39958 24376 40010
rect 24424 39958 24448 40010
rect 24448 39958 24480 40010
rect 24528 39958 24572 40010
rect 24572 39958 24584 40010
rect 24320 39956 24376 39958
rect 24424 39956 24480 39958
rect 24528 39956 24584 39958
rect 24632 40010 24688 40012
rect 24736 40010 24792 40012
rect 24840 40010 24896 40012
rect 24632 39958 24644 40010
rect 24644 39958 24688 40010
rect 24736 39958 24768 40010
rect 24768 39958 24792 40010
rect 24840 39958 24892 40010
rect 24892 39958 24896 40010
rect 24632 39956 24688 39958
rect 24736 39956 24792 39958
rect 24840 39956 24896 39958
rect 24944 39956 25000 40012
rect 25048 40010 25104 40012
rect 25152 40010 25208 40012
rect 25048 39958 25068 40010
rect 25068 39958 25104 40010
rect 25152 39958 25192 40010
rect 25192 39958 25208 40010
rect 25048 39956 25104 39958
rect 25152 39956 25208 39958
rect 14008 39226 14064 39228
rect 14112 39226 14168 39228
rect 14008 39174 14024 39226
rect 14024 39174 14064 39226
rect 14112 39174 14148 39226
rect 14148 39174 14168 39226
rect 14008 39172 14064 39174
rect 14112 39172 14168 39174
rect 14216 39172 14272 39228
rect 14320 39226 14376 39228
rect 14424 39226 14480 39228
rect 14528 39226 14584 39228
rect 14320 39174 14324 39226
rect 14324 39174 14376 39226
rect 14424 39174 14448 39226
rect 14448 39174 14480 39226
rect 14528 39174 14572 39226
rect 14572 39174 14584 39226
rect 14320 39172 14376 39174
rect 14424 39172 14480 39174
rect 14528 39172 14584 39174
rect 14632 39226 14688 39228
rect 14736 39226 14792 39228
rect 14840 39226 14896 39228
rect 14632 39174 14644 39226
rect 14644 39174 14688 39226
rect 14736 39174 14768 39226
rect 14768 39174 14792 39226
rect 14840 39174 14892 39226
rect 14892 39174 14896 39226
rect 14632 39172 14688 39174
rect 14736 39172 14792 39174
rect 14840 39172 14896 39174
rect 14944 39172 15000 39228
rect 15048 39226 15104 39228
rect 15152 39226 15208 39228
rect 15048 39174 15068 39226
rect 15068 39174 15104 39226
rect 15152 39174 15192 39226
rect 15192 39174 15208 39226
rect 15048 39172 15104 39174
rect 15152 39172 15208 39174
rect 24008 38442 24064 38444
rect 24112 38442 24168 38444
rect 24008 38390 24024 38442
rect 24024 38390 24064 38442
rect 24112 38390 24148 38442
rect 24148 38390 24168 38442
rect 24008 38388 24064 38390
rect 24112 38388 24168 38390
rect 24216 38388 24272 38444
rect 24320 38442 24376 38444
rect 24424 38442 24480 38444
rect 24528 38442 24584 38444
rect 24320 38390 24324 38442
rect 24324 38390 24376 38442
rect 24424 38390 24448 38442
rect 24448 38390 24480 38442
rect 24528 38390 24572 38442
rect 24572 38390 24584 38442
rect 24320 38388 24376 38390
rect 24424 38388 24480 38390
rect 24528 38388 24584 38390
rect 24632 38442 24688 38444
rect 24736 38442 24792 38444
rect 24840 38442 24896 38444
rect 24632 38390 24644 38442
rect 24644 38390 24688 38442
rect 24736 38390 24768 38442
rect 24768 38390 24792 38442
rect 24840 38390 24892 38442
rect 24892 38390 24896 38442
rect 24632 38388 24688 38390
rect 24736 38388 24792 38390
rect 24840 38388 24896 38390
rect 24944 38388 25000 38444
rect 25048 38442 25104 38444
rect 25152 38442 25208 38444
rect 25048 38390 25068 38442
rect 25068 38390 25104 38442
rect 25152 38390 25192 38442
rect 25192 38390 25208 38442
rect 25048 38388 25104 38390
rect 25152 38388 25208 38390
rect 14008 37658 14064 37660
rect 14112 37658 14168 37660
rect 14008 37606 14024 37658
rect 14024 37606 14064 37658
rect 14112 37606 14148 37658
rect 14148 37606 14168 37658
rect 14008 37604 14064 37606
rect 14112 37604 14168 37606
rect 14216 37604 14272 37660
rect 14320 37658 14376 37660
rect 14424 37658 14480 37660
rect 14528 37658 14584 37660
rect 14320 37606 14324 37658
rect 14324 37606 14376 37658
rect 14424 37606 14448 37658
rect 14448 37606 14480 37658
rect 14528 37606 14572 37658
rect 14572 37606 14584 37658
rect 14320 37604 14376 37606
rect 14424 37604 14480 37606
rect 14528 37604 14584 37606
rect 14632 37658 14688 37660
rect 14736 37658 14792 37660
rect 14840 37658 14896 37660
rect 14632 37606 14644 37658
rect 14644 37606 14688 37658
rect 14736 37606 14768 37658
rect 14768 37606 14792 37658
rect 14840 37606 14892 37658
rect 14892 37606 14896 37658
rect 14632 37604 14688 37606
rect 14736 37604 14792 37606
rect 14840 37604 14896 37606
rect 14944 37604 15000 37660
rect 15048 37658 15104 37660
rect 15152 37658 15208 37660
rect 15048 37606 15068 37658
rect 15068 37606 15104 37658
rect 15152 37606 15192 37658
rect 15192 37606 15208 37658
rect 15048 37604 15104 37606
rect 15152 37604 15208 37606
rect 24008 36874 24064 36876
rect 24112 36874 24168 36876
rect 24008 36822 24024 36874
rect 24024 36822 24064 36874
rect 24112 36822 24148 36874
rect 24148 36822 24168 36874
rect 24008 36820 24064 36822
rect 24112 36820 24168 36822
rect 24216 36820 24272 36876
rect 24320 36874 24376 36876
rect 24424 36874 24480 36876
rect 24528 36874 24584 36876
rect 24320 36822 24324 36874
rect 24324 36822 24376 36874
rect 24424 36822 24448 36874
rect 24448 36822 24480 36874
rect 24528 36822 24572 36874
rect 24572 36822 24584 36874
rect 24320 36820 24376 36822
rect 24424 36820 24480 36822
rect 24528 36820 24584 36822
rect 24632 36874 24688 36876
rect 24736 36874 24792 36876
rect 24840 36874 24896 36876
rect 24632 36822 24644 36874
rect 24644 36822 24688 36874
rect 24736 36822 24768 36874
rect 24768 36822 24792 36874
rect 24840 36822 24892 36874
rect 24892 36822 24896 36874
rect 24632 36820 24688 36822
rect 24736 36820 24792 36822
rect 24840 36820 24896 36822
rect 24944 36820 25000 36876
rect 25048 36874 25104 36876
rect 25152 36874 25208 36876
rect 25048 36822 25068 36874
rect 25068 36822 25104 36874
rect 25152 36822 25192 36874
rect 25192 36822 25208 36874
rect 25048 36820 25104 36822
rect 25152 36820 25208 36822
rect 14008 36090 14064 36092
rect 14112 36090 14168 36092
rect 14008 36038 14024 36090
rect 14024 36038 14064 36090
rect 14112 36038 14148 36090
rect 14148 36038 14168 36090
rect 14008 36036 14064 36038
rect 14112 36036 14168 36038
rect 14216 36036 14272 36092
rect 14320 36090 14376 36092
rect 14424 36090 14480 36092
rect 14528 36090 14584 36092
rect 14320 36038 14324 36090
rect 14324 36038 14376 36090
rect 14424 36038 14448 36090
rect 14448 36038 14480 36090
rect 14528 36038 14572 36090
rect 14572 36038 14584 36090
rect 14320 36036 14376 36038
rect 14424 36036 14480 36038
rect 14528 36036 14584 36038
rect 14632 36090 14688 36092
rect 14736 36090 14792 36092
rect 14840 36090 14896 36092
rect 14632 36038 14644 36090
rect 14644 36038 14688 36090
rect 14736 36038 14768 36090
rect 14768 36038 14792 36090
rect 14840 36038 14892 36090
rect 14892 36038 14896 36090
rect 14632 36036 14688 36038
rect 14736 36036 14792 36038
rect 14840 36036 14896 36038
rect 14944 36036 15000 36092
rect 15048 36090 15104 36092
rect 15152 36090 15208 36092
rect 15048 36038 15068 36090
rect 15068 36038 15104 36090
rect 15152 36038 15192 36090
rect 15192 36038 15208 36090
rect 15048 36036 15104 36038
rect 15152 36036 15208 36038
rect 24008 35306 24064 35308
rect 24112 35306 24168 35308
rect 24008 35254 24024 35306
rect 24024 35254 24064 35306
rect 24112 35254 24148 35306
rect 24148 35254 24168 35306
rect 24008 35252 24064 35254
rect 24112 35252 24168 35254
rect 24216 35252 24272 35308
rect 24320 35306 24376 35308
rect 24424 35306 24480 35308
rect 24528 35306 24584 35308
rect 24320 35254 24324 35306
rect 24324 35254 24376 35306
rect 24424 35254 24448 35306
rect 24448 35254 24480 35306
rect 24528 35254 24572 35306
rect 24572 35254 24584 35306
rect 24320 35252 24376 35254
rect 24424 35252 24480 35254
rect 24528 35252 24584 35254
rect 24632 35306 24688 35308
rect 24736 35306 24792 35308
rect 24840 35306 24896 35308
rect 24632 35254 24644 35306
rect 24644 35254 24688 35306
rect 24736 35254 24768 35306
rect 24768 35254 24792 35306
rect 24840 35254 24892 35306
rect 24892 35254 24896 35306
rect 24632 35252 24688 35254
rect 24736 35252 24792 35254
rect 24840 35252 24896 35254
rect 24944 35252 25000 35308
rect 25048 35306 25104 35308
rect 25152 35306 25208 35308
rect 25048 35254 25068 35306
rect 25068 35254 25104 35306
rect 25152 35254 25192 35306
rect 25192 35254 25208 35306
rect 25048 35252 25104 35254
rect 25152 35252 25208 35254
rect 14008 34522 14064 34524
rect 14112 34522 14168 34524
rect 14008 34470 14024 34522
rect 14024 34470 14064 34522
rect 14112 34470 14148 34522
rect 14148 34470 14168 34522
rect 14008 34468 14064 34470
rect 14112 34468 14168 34470
rect 14216 34468 14272 34524
rect 14320 34522 14376 34524
rect 14424 34522 14480 34524
rect 14528 34522 14584 34524
rect 14320 34470 14324 34522
rect 14324 34470 14376 34522
rect 14424 34470 14448 34522
rect 14448 34470 14480 34522
rect 14528 34470 14572 34522
rect 14572 34470 14584 34522
rect 14320 34468 14376 34470
rect 14424 34468 14480 34470
rect 14528 34468 14584 34470
rect 14632 34522 14688 34524
rect 14736 34522 14792 34524
rect 14840 34522 14896 34524
rect 14632 34470 14644 34522
rect 14644 34470 14688 34522
rect 14736 34470 14768 34522
rect 14768 34470 14792 34522
rect 14840 34470 14892 34522
rect 14892 34470 14896 34522
rect 14632 34468 14688 34470
rect 14736 34468 14792 34470
rect 14840 34468 14896 34470
rect 14944 34468 15000 34524
rect 15048 34522 15104 34524
rect 15152 34522 15208 34524
rect 15048 34470 15068 34522
rect 15068 34470 15104 34522
rect 15152 34470 15192 34522
rect 15192 34470 15208 34522
rect 15048 34468 15104 34470
rect 15152 34468 15208 34470
rect 24008 33738 24064 33740
rect 24112 33738 24168 33740
rect 24008 33686 24024 33738
rect 24024 33686 24064 33738
rect 24112 33686 24148 33738
rect 24148 33686 24168 33738
rect 24008 33684 24064 33686
rect 24112 33684 24168 33686
rect 24216 33684 24272 33740
rect 24320 33738 24376 33740
rect 24424 33738 24480 33740
rect 24528 33738 24584 33740
rect 24320 33686 24324 33738
rect 24324 33686 24376 33738
rect 24424 33686 24448 33738
rect 24448 33686 24480 33738
rect 24528 33686 24572 33738
rect 24572 33686 24584 33738
rect 24320 33684 24376 33686
rect 24424 33684 24480 33686
rect 24528 33684 24584 33686
rect 24632 33738 24688 33740
rect 24736 33738 24792 33740
rect 24840 33738 24896 33740
rect 24632 33686 24644 33738
rect 24644 33686 24688 33738
rect 24736 33686 24768 33738
rect 24768 33686 24792 33738
rect 24840 33686 24892 33738
rect 24892 33686 24896 33738
rect 24632 33684 24688 33686
rect 24736 33684 24792 33686
rect 24840 33684 24896 33686
rect 24944 33684 25000 33740
rect 25048 33738 25104 33740
rect 25152 33738 25208 33740
rect 25048 33686 25068 33738
rect 25068 33686 25104 33738
rect 25152 33686 25192 33738
rect 25192 33686 25208 33738
rect 25048 33684 25104 33686
rect 25152 33684 25208 33686
rect 14008 32954 14064 32956
rect 14112 32954 14168 32956
rect 14008 32902 14024 32954
rect 14024 32902 14064 32954
rect 14112 32902 14148 32954
rect 14148 32902 14168 32954
rect 14008 32900 14064 32902
rect 14112 32900 14168 32902
rect 14216 32900 14272 32956
rect 14320 32954 14376 32956
rect 14424 32954 14480 32956
rect 14528 32954 14584 32956
rect 14320 32902 14324 32954
rect 14324 32902 14376 32954
rect 14424 32902 14448 32954
rect 14448 32902 14480 32954
rect 14528 32902 14572 32954
rect 14572 32902 14584 32954
rect 14320 32900 14376 32902
rect 14424 32900 14480 32902
rect 14528 32900 14584 32902
rect 14632 32954 14688 32956
rect 14736 32954 14792 32956
rect 14840 32954 14896 32956
rect 14632 32902 14644 32954
rect 14644 32902 14688 32954
rect 14736 32902 14768 32954
rect 14768 32902 14792 32954
rect 14840 32902 14892 32954
rect 14892 32902 14896 32954
rect 14632 32900 14688 32902
rect 14736 32900 14792 32902
rect 14840 32900 14896 32902
rect 14944 32900 15000 32956
rect 15048 32954 15104 32956
rect 15152 32954 15208 32956
rect 15048 32902 15068 32954
rect 15068 32902 15104 32954
rect 15152 32902 15192 32954
rect 15192 32902 15208 32954
rect 15048 32900 15104 32902
rect 15152 32900 15208 32902
rect 24008 32170 24064 32172
rect 24112 32170 24168 32172
rect 24008 32118 24024 32170
rect 24024 32118 24064 32170
rect 24112 32118 24148 32170
rect 24148 32118 24168 32170
rect 24008 32116 24064 32118
rect 24112 32116 24168 32118
rect 24216 32116 24272 32172
rect 24320 32170 24376 32172
rect 24424 32170 24480 32172
rect 24528 32170 24584 32172
rect 24320 32118 24324 32170
rect 24324 32118 24376 32170
rect 24424 32118 24448 32170
rect 24448 32118 24480 32170
rect 24528 32118 24572 32170
rect 24572 32118 24584 32170
rect 24320 32116 24376 32118
rect 24424 32116 24480 32118
rect 24528 32116 24584 32118
rect 24632 32170 24688 32172
rect 24736 32170 24792 32172
rect 24840 32170 24896 32172
rect 24632 32118 24644 32170
rect 24644 32118 24688 32170
rect 24736 32118 24768 32170
rect 24768 32118 24792 32170
rect 24840 32118 24892 32170
rect 24892 32118 24896 32170
rect 24632 32116 24688 32118
rect 24736 32116 24792 32118
rect 24840 32116 24896 32118
rect 24944 32116 25000 32172
rect 25048 32170 25104 32172
rect 25152 32170 25208 32172
rect 25048 32118 25068 32170
rect 25068 32118 25104 32170
rect 25152 32118 25192 32170
rect 25192 32118 25208 32170
rect 25048 32116 25104 32118
rect 25152 32116 25208 32118
rect 14008 31386 14064 31388
rect 14112 31386 14168 31388
rect 14008 31334 14024 31386
rect 14024 31334 14064 31386
rect 14112 31334 14148 31386
rect 14148 31334 14168 31386
rect 14008 31332 14064 31334
rect 14112 31332 14168 31334
rect 14216 31332 14272 31388
rect 14320 31386 14376 31388
rect 14424 31386 14480 31388
rect 14528 31386 14584 31388
rect 14320 31334 14324 31386
rect 14324 31334 14376 31386
rect 14424 31334 14448 31386
rect 14448 31334 14480 31386
rect 14528 31334 14572 31386
rect 14572 31334 14584 31386
rect 14320 31332 14376 31334
rect 14424 31332 14480 31334
rect 14528 31332 14584 31334
rect 14632 31386 14688 31388
rect 14736 31386 14792 31388
rect 14840 31386 14896 31388
rect 14632 31334 14644 31386
rect 14644 31334 14688 31386
rect 14736 31334 14768 31386
rect 14768 31334 14792 31386
rect 14840 31334 14892 31386
rect 14892 31334 14896 31386
rect 14632 31332 14688 31334
rect 14736 31332 14792 31334
rect 14840 31332 14896 31334
rect 14944 31332 15000 31388
rect 15048 31386 15104 31388
rect 15152 31386 15208 31388
rect 15048 31334 15068 31386
rect 15068 31334 15104 31386
rect 15152 31334 15192 31386
rect 15192 31334 15208 31386
rect 15048 31332 15104 31334
rect 15152 31332 15208 31334
rect 24008 30602 24064 30604
rect 24112 30602 24168 30604
rect 24008 30550 24024 30602
rect 24024 30550 24064 30602
rect 24112 30550 24148 30602
rect 24148 30550 24168 30602
rect 24008 30548 24064 30550
rect 24112 30548 24168 30550
rect 24216 30548 24272 30604
rect 24320 30602 24376 30604
rect 24424 30602 24480 30604
rect 24528 30602 24584 30604
rect 24320 30550 24324 30602
rect 24324 30550 24376 30602
rect 24424 30550 24448 30602
rect 24448 30550 24480 30602
rect 24528 30550 24572 30602
rect 24572 30550 24584 30602
rect 24320 30548 24376 30550
rect 24424 30548 24480 30550
rect 24528 30548 24584 30550
rect 24632 30602 24688 30604
rect 24736 30602 24792 30604
rect 24840 30602 24896 30604
rect 24632 30550 24644 30602
rect 24644 30550 24688 30602
rect 24736 30550 24768 30602
rect 24768 30550 24792 30602
rect 24840 30550 24892 30602
rect 24892 30550 24896 30602
rect 24632 30548 24688 30550
rect 24736 30548 24792 30550
rect 24840 30548 24896 30550
rect 24944 30548 25000 30604
rect 25048 30602 25104 30604
rect 25152 30602 25208 30604
rect 25048 30550 25068 30602
rect 25068 30550 25104 30602
rect 25152 30550 25192 30602
rect 25192 30550 25208 30602
rect 25048 30548 25104 30550
rect 25152 30548 25208 30550
rect 14008 29818 14064 29820
rect 14112 29818 14168 29820
rect 14008 29766 14024 29818
rect 14024 29766 14064 29818
rect 14112 29766 14148 29818
rect 14148 29766 14168 29818
rect 14008 29764 14064 29766
rect 14112 29764 14168 29766
rect 14216 29764 14272 29820
rect 14320 29818 14376 29820
rect 14424 29818 14480 29820
rect 14528 29818 14584 29820
rect 14320 29766 14324 29818
rect 14324 29766 14376 29818
rect 14424 29766 14448 29818
rect 14448 29766 14480 29818
rect 14528 29766 14572 29818
rect 14572 29766 14584 29818
rect 14320 29764 14376 29766
rect 14424 29764 14480 29766
rect 14528 29764 14584 29766
rect 14632 29818 14688 29820
rect 14736 29818 14792 29820
rect 14840 29818 14896 29820
rect 14632 29766 14644 29818
rect 14644 29766 14688 29818
rect 14736 29766 14768 29818
rect 14768 29766 14792 29818
rect 14840 29766 14892 29818
rect 14892 29766 14896 29818
rect 14632 29764 14688 29766
rect 14736 29764 14792 29766
rect 14840 29764 14896 29766
rect 14944 29764 15000 29820
rect 15048 29818 15104 29820
rect 15152 29818 15208 29820
rect 15048 29766 15068 29818
rect 15068 29766 15104 29818
rect 15152 29766 15192 29818
rect 15192 29766 15208 29818
rect 15048 29764 15104 29766
rect 15152 29764 15208 29766
rect 24008 29034 24064 29036
rect 24112 29034 24168 29036
rect 24008 28982 24024 29034
rect 24024 28982 24064 29034
rect 24112 28982 24148 29034
rect 24148 28982 24168 29034
rect 24008 28980 24064 28982
rect 24112 28980 24168 28982
rect 24216 28980 24272 29036
rect 24320 29034 24376 29036
rect 24424 29034 24480 29036
rect 24528 29034 24584 29036
rect 24320 28982 24324 29034
rect 24324 28982 24376 29034
rect 24424 28982 24448 29034
rect 24448 28982 24480 29034
rect 24528 28982 24572 29034
rect 24572 28982 24584 29034
rect 24320 28980 24376 28982
rect 24424 28980 24480 28982
rect 24528 28980 24584 28982
rect 24632 29034 24688 29036
rect 24736 29034 24792 29036
rect 24840 29034 24896 29036
rect 24632 28982 24644 29034
rect 24644 28982 24688 29034
rect 24736 28982 24768 29034
rect 24768 28982 24792 29034
rect 24840 28982 24892 29034
rect 24892 28982 24896 29034
rect 24632 28980 24688 28982
rect 24736 28980 24792 28982
rect 24840 28980 24896 28982
rect 24944 28980 25000 29036
rect 25048 29034 25104 29036
rect 25152 29034 25208 29036
rect 25048 28982 25068 29034
rect 25068 28982 25104 29034
rect 25152 28982 25192 29034
rect 25192 28982 25208 29034
rect 25048 28980 25104 28982
rect 25152 28980 25208 28982
rect 14008 28250 14064 28252
rect 14112 28250 14168 28252
rect 14008 28198 14024 28250
rect 14024 28198 14064 28250
rect 14112 28198 14148 28250
rect 14148 28198 14168 28250
rect 14008 28196 14064 28198
rect 14112 28196 14168 28198
rect 14216 28196 14272 28252
rect 14320 28250 14376 28252
rect 14424 28250 14480 28252
rect 14528 28250 14584 28252
rect 14320 28198 14324 28250
rect 14324 28198 14376 28250
rect 14424 28198 14448 28250
rect 14448 28198 14480 28250
rect 14528 28198 14572 28250
rect 14572 28198 14584 28250
rect 14320 28196 14376 28198
rect 14424 28196 14480 28198
rect 14528 28196 14584 28198
rect 14632 28250 14688 28252
rect 14736 28250 14792 28252
rect 14840 28250 14896 28252
rect 14632 28198 14644 28250
rect 14644 28198 14688 28250
rect 14736 28198 14768 28250
rect 14768 28198 14792 28250
rect 14840 28198 14892 28250
rect 14892 28198 14896 28250
rect 14632 28196 14688 28198
rect 14736 28196 14792 28198
rect 14840 28196 14896 28198
rect 14944 28196 15000 28252
rect 15048 28250 15104 28252
rect 15152 28250 15208 28252
rect 15048 28198 15068 28250
rect 15068 28198 15104 28250
rect 15152 28198 15192 28250
rect 15192 28198 15208 28250
rect 15048 28196 15104 28198
rect 15152 28196 15208 28198
rect 24008 27466 24064 27468
rect 24112 27466 24168 27468
rect 24008 27414 24024 27466
rect 24024 27414 24064 27466
rect 24112 27414 24148 27466
rect 24148 27414 24168 27466
rect 24008 27412 24064 27414
rect 24112 27412 24168 27414
rect 24216 27412 24272 27468
rect 24320 27466 24376 27468
rect 24424 27466 24480 27468
rect 24528 27466 24584 27468
rect 24320 27414 24324 27466
rect 24324 27414 24376 27466
rect 24424 27414 24448 27466
rect 24448 27414 24480 27466
rect 24528 27414 24572 27466
rect 24572 27414 24584 27466
rect 24320 27412 24376 27414
rect 24424 27412 24480 27414
rect 24528 27412 24584 27414
rect 24632 27466 24688 27468
rect 24736 27466 24792 27468
rect 24840 27466 24896 27468
rect 24632 27414 24644 27466
rect 24644 27414 24688 27466
rect 24736 27414 24768 27466
rect 24768 27414 24792 27466
rect 24840 27414 24892 27466
rect 24892 27414 24896 27466
rect 24632 27412 24688 27414
rect 24736 27412 24792 27414
rect 24840 27412 24896 27414
rect 24944 27412 25000 27468
rect 25048 27466 25104 27468
rect 25152 27466 25208 27468
rect 25048 27414 25068 27466
rect 25068 27414 25104 27466
rect 25152 27414 25192 27466
rect 25192 27414 25208 27466
rect 25048 27412 25104 27414
rect 25152 27412 25208 27414
rect 14008 26682 14064 26684
rect 14112 26682 14168 26684
rect 14008 26630 14024 26682
rect 14024 26630 14064 26682
rect 14112 26630 14148 26682
rect 14148 26630 14168 26682
rect 14008 26628 14064 26630
rect 14112 26628 14168 26630
rect 14216 26628 14272 26684
rect 14320 26682 14376 26684
rect 14424 26682 14480 26684
rect 14528 26682 14584 26684
rect 14320 26630 14324 26682
rect 14324 26630 14376 26682
rect 14424 26630 14448 26682
rect 14448 26630 14480 26682
rect 14528 26630 14572 26682
rect 14572 26630 14584 26682
rect 14320 26628 14376 26630
rect 14424 26628 14480 26630
rect 14528 26628 14584 26630
rect 14632 26682 14688 26684
rect 14736 26682 14792 26684
rect 14840 26682 14896 26684
rect 14632 26630 14644 26682
rect 14644 26630 14688 26682
rect 14736 26630 14768 26682
rect 14768 26630 14792 26682
rect 14840 26630 14892 26682
rect 14892 26630 14896 26682
rect 14632 26628 14688 26630
rect 14736 26628 14792 26630
rect 14840 26628 14896 26630
rect 14944 26628 15000 26684
rect 15048 26682 15104 26684
rect 15152 26682 15208 26684
rect 15048 26630 15068 26682
rect 15068 26630 15104 26682
rect 15152 26630 15192 26682
rect 15192 26630 15208 26682
rect 15048 26628 15104 26630
rect 15152 26628 15208 26630
rect 24008 25898 24064 25900
rect 24112 25898 24168 25900
rect 24008 25846 24024 25898
rect 24024 25846 24064 25898
rect 24112 25846 24148 25898
rect 24148 25846 24168 25898
rect 24008 25844 24064 25846
rect 24112 25844 24168 25846
rect 24216 25844 24272 25900
rect 24320 25898 24376 25900
rect 24424 25898 24480 25900
rect 24528 25898 24584 25900
rect 24320 25846 24324 25898
rect 24324 25846 24376 25898
rect 24424 25846 24448 25898
rect 24448 25846 24480 25898
rect 24528 25846 24572 25898
rect 24572 25846 24584 25898
rect 24320 25844 24376 25846
rect 24424 25844 24480 25846
rect 24528 25844 24584 25846
rect 24632 25898 24688 25900
rect 24736 25898 24792 25900
rect 24840 25898 24896 25900
rect 24632 25846 24644 25898
rect 24644 25846 24688 25898
rect 24736 25846 24768 25898
rect 24768 25846 24792 25898
rect 24840 25846 24892 25898
rect 24892 25846 24896 25898
rect 24632 25844 24688 25846
rect 24736 25844 24792 25846
rect 24840 25844 24896 25846
rect 24944 25844 25000 25900
rect 25048 25898 25104 25900
rect 25152 25898 25208 25900
rect 25048 25846 25068 25898
rect 25068 25846 25104 25898
rect 25152 25846 25192 25898
rect 25192 25846 25208 25898
rect 25048 25844 25104 25846
rect 25152 25844 25208 25846
rect 14008 25114 14064 25116
rect 14112 25114 14168 25116
rect 14008 25062 14024 25114
rect 14024 25062 14064 25114
rect 14112 25062 14148 25114
rect 14148 25062 14168 25114
rect 14008 25060 14064 25062
rect 14112 25060 14168 25062
rect 14216 25060 14272 25116
rect 14320 25114 14376 25116
rect 14424 25114 14480 25116
rect 14528 25114 14584 25116
rect 14320 25062 14324 25114
rect 14324 25062 14376 25114
rect 14424 25062 14448 25114
rect 14448 25062 14480 25114
rect 14528 25062 14572 25114
rect 14572 25062 14584 25114
rect 14320 25060 14376 25062
rect 14424 25060 14480 25062
rect 14528 25060 14584 25062
rect 14632 25114 14688 25116
rect 14736 25114 14792 25116
rect 14840 25114 14896 25116
rect 14632 25062 14644 25114
rect 14644 25062 14688 25114
rect 14736 25062 14768 25114
rect 14768 25062 14792 25114
rect 14840 25062 14892 25114
rect 14892 25062 14896 25114
rect 14632 25060 14688 25062
rect 14736 25060 14792 25062
rect 14840 25060 14896 25062
rect 14944 25060 15000 25116
rect 15048 25114 15104 25116
rect 15152 25114 15208 25116
rect 15048 25062 15068 25114
rect 15068 25062 15104 25114
rect 15152 25062 15192 25114
rect 15192 25062 15208 25114
rect 15048 25060 15104 25062
rect 15152 25060 15208 25062
rect 24008 24330 24064 24332
rect 24112 24330 24168 24332
rect 24008 24278 24024 24330
rect 24024 24278 24064 24330
rect 24112 24278 24148 24330
rect 24148 24278 24168 24330
rect 24008 24276 24064 24278
rect 24112 24276 24168 24278
rect 24216 24276 24272 24332
rect 24320 24330 24376 24332
rect 24424 24330 24480 24332
rect 24528 24330 24584 24332
rect 24320 24278 24324 24330
rect 24324 24278 24376 24330
rect 24424 24278 24448 24330
rect 24448 24278 24480 24330
rect 24528 24278 24572 24330
rect 24572 24278 24584 24330
rect 24320 24276 24376 24278
rect 24424 24276 24480 24278
rect 24528 24276 24584 24278
rect 24632 24330 24688 24332
rect 24736 24330 24792 24332
rect 24840 24330 24896 24332
rect 24632 24278 24644 24330
rect 24644 24278 24688 24330
rect 24736 24278 24768 24330
rect 24768 24278 24792 24330
rect 24840 24278 24892 24330
rect 24892 24278 24896 24330
rect 24632 24276 24688 24278
rect 24736 24276 24792 24278
rect 24840 24276 24896 24278
rect 24944 24276 25000 24332
rect 25048 24330 25104 24332
rect 25152 24330 25208 24332
rect 25048 24278 25068 24330
rect 25068 24278 25104 24330
rect 25152 24278 25192 24330
rect 25192 24278 25208 24330
rect 25048 24276 25104 24278
rect 25152 24276 25208 24278
rect 14008 23546 14064 23548
rect 14112 23546 14168 23548
rect 14008 23494 14024 23546
rect 14024 23494 14064 23546
rect 14112 23494 14148 23546
rect 14148 23494 14168 23546
rect 14008 23492 14064 23494
rect 14112 23492 14168 23494
rect 14216 23492 14272 23548
rect 14320 23546 14376 23548
rect 14424 23546 14480 23548
rect 14528 23546 14584 23548
rect 14320 23494 14324 23546
rect 14324 23494 14376 23546
rect 14424 23494 14448 23546
rect 14448 23494 14480 23546
rect 14528 23494 14572 23546
rect 14572 23494 14584 23546
rect 14320 23492 14376 23494
rect 14424 23492 14480 23494
rect 14528 23492 14584 23494
rect 14632 23546 14688 23548
rect 14736 23546 14792 23548
rect 14840 23546 14896 23548
rect 14632 23494 14644 23546
rect 14644 23494 14688 23546
rect 14736 23494 14768 23546
rect 14768 23494 14792 23546
rect 14840 23494 14892 23546
rect 14892 23494 14896 23546
rect 14632 23492 14688 23494
rect 14736 23492 14792 23494
rect 14840 23492 14896 23494
rect 14944 23492 15000 23548
rect 15048 23546 15104 23548
rect 15152 23546 15208 23548
rect 15048 23494 15068 23546
rect 15068 23494 15104 23546
rect 15152 23494 15192 23546
rect 15192 23494 15208 23546
rect 15048 23492 15104 23494
rect 15152 23492 15208 23494
rect 24008 22762 24064 22764
rect 24112 22762 24168 22764
rect 24008 22710 24024 22762
rect 24024 22710 24064 22762
rect 24112 22710 24148 22762
rect 24148 22710 24168 22762
rect 24008 22708 24064 22710
rect 24112 22708 24168 22710
rect 24216 22708 24272 22764
rect 24320 22762 24376 22764
rect 24424 22762 24480 22764
rect 24528 22762 24584 22764
rect 24320 22710 24324 22762
rect 24324 22710 24376 22762
rect 24424 22710 24448 22762
rect 24448 22710 24480 22762
rect 24528 22710 24572 22762
rect 24572 22710 24584 22762
rect 24320 22708 24376 22710
rect 24424 22708 24480 22710
rect 24528 22708 24584 22710
rect 24632 22762 24688 22764
rect 24736 22762 24792 22764
rect 24840 22762 24896 22764
rect 24632 22710 24644 22762
rect 24644 22710 24688 22762
rect 24736 22710 24768 22762
rect 24768 22710 24792 22762
rect 24840 22710 24892 22762
rect 24892 22710 24896 22762
rect 24632 22708 24688 22710
rect 24736 22708 24792 22710
rect 24840 22708 24896 22710
rect 24944 22708 25000 22764
rect 25048 22762 25104 22764
rect 25152 22762 25208 22764
rect 25048 22710 25068 22762
rect 25068 22710 25104 22762
rect 25152 22710 25192 22762
rect 25192 22710 25208 22762
rect 25048 22708 25104 22710
rect 25152 22708 25208 22710
rect 14008 21978 14064 21980
rect 14112 21978 14168 21980
rect 14008 21926 14024 21978
rect 14024 21926 14064 21978
rect 14112 21926 14148 21978
rect 14148 21926 14168 21978
rect 14008 21924 14064 21926
rect 14112 21924 14168 21926
rect 14216 21924 14272 21980
rect 14320 21978 14376 21980
rect 14424 21978 14480 21980
rect 14528 21978 14584 21980
rect 14320 21926 14324 21978
rect 14324 21926 14376 21978
rect 14424 21926 14448 21978
rect 14448 21926 14480 21978
rect 14528 21926 14572 21978
rect 14572 21926 14584 21978
rect 14320 21924 14376 21926
rect 14424 21924 14480 21926
rect 14528 21924 14584 21926
rect 14632 21978 14688 21980
rect 14736 21978 14792 21980
rect 14840 21978 14896 21980
rect 14632 21926 14644 21978
rect 14644 21926 14688 21978
rect 14736 21926 14768 21978
rect 14768 21926 14792 21978
rect 14840 21926 14892 21978
rect 14892 21926 14896 21978
rect 14632 21924 14688 21926
rect 14736 21924 14792 21926
rect 14840 21924 14896 21926
rect 14944 21924 15000 21980
rect 15048 21978 15104 21980
rect 15152 21978 15208 21980
rect 15048 21926 15068 21978
rect 15068 21926 15104 21978
rect 15152 21926 15192 21978
rect 15192 21926 15208 21978
rect 15048 21924 15104 21926
rect 15152 21924 15208 21926
rect 24008 21194 24064 21196
rect 24112 21194 24168 21196
rect 24008 21142 24024 21194
rect 24024 21142 24064 21194
rect 24112 21142 24148 21194
rect 24148 21142 24168 21194
rect 24008 21140 24064 21142
rect 24112 21140 24168 21142
rect 24216 21140 24272 21196
rect 24320 21194 24376 21196
rect 24424 21194 24480 21196
rect 24528 21194 24584 21196
rect 24320 21142 24324 21194
rect 24324 21142 24376 21194
rect 24424 21142 24448 21194
rect 24448 21142 24480 21194
rect 24528 21142 24572 21194
rect 24572 21142 24584 21194
rect 24320 21140 24376 21142
rect 24424 21140 24480 21142
rect 24528 21140 24584 21142
rect 24632 21194 24688 21196
rect 24736 21194 24792 21196
rect 24840 21194 24896 21196
rect 24632 21142 24644 21194
rect 24644 21142 24688 21194
rect 24736 21142 24768 21194
rect 24768 21142 24792 21194
rect 24840 21142 24892 21194
rect 24892 21142 24896 21194
rect 24632 21140 24688 21142
rect 24736 21140 24792 21142
rect 24840 21140 24896 21142
rect 24944 21140 25000 21196
rect 25048 21194 25104 21196
rect 25152 21194 25208 21196
rect 25048 21142 25068 21194
rect 25068 21142 25104 21194
rect 25152 21142 25192 21194
rect 25192 21142 25208 21194
rect 25048 21140 25104 21142
rect 25152 21140 25208 21142
rect 14008 20410 14064 20412
rect 14112 20410 14168 20412
rect 14008 20358 14024 20410
rect 14024 20358 14064 20410
rect 14112 20358 14148 20410
rect 14148 20358 14168 20410
rect 14008 20356 14064 20358
rect 14112 20356 14168 20358
rect 14216 20356 14272 20412
rect 14320 20410 14376 20412
rect 14424 20410 14480 20412
rect 14528 20410 14584 20412
rect 14320 20358 14324 20410
rect 14324 20358 14376 20410
rect 14424 20358 14448 20410
rect 14448 20358 14480 20410
rect 14528 20358 14572 20410
rect 14572 20358 14584 20410
rect 14320 20356 14376 20358
rect 14424 20356 14480 20358
rect 14528 20356 14584 20358
rect 14632 20410 14688 20412
rect 14736 20410 14792 20412
rect 14840 20410 14896 20412
rect 14632 20358 14644 20410
rect 14644 20358 14688 20410
rect 14736 20358 14768 20410
rect 14768 20358 14792 20410
rect 14840 20358 14892 20410
rect 14892 20358 14896 20410
rect 14632 20356 14688 20358
rect 14736 20356 14792 20358
rect 14840 20356 14896 20358
rect 14944 20356 15000 20412
rect 15048 20410 15104 20412
rect 15152 20410 15208 20412
rect 15048 20358 15068 20410
rect 15068 20358 15104 20410
rect 15152 20358 15192 20410
rect 15192 20358 15208 20410
rect 15048 20356 15104 20358
rect 15152 20356 15208 20358
rect 24008 19626 24064 19628
rect 24112 19626 24168 19628
rect 24008 19574 24024 19626
rect 24024 19574 24064 19626
rect 24112 19574 24148 19626
rect 24148 19574 24168 19626
rect 24008 19572 24064 19574
rect 24112 19572 24168 19574
rect 24216 19572 24272 19628
rect 24320 19626 24376 19628
rect 24424 19626 24480 19628
rect 24528 19626 24584 19628
rect 24320 19574 24324 19626
rect 24324 19574 24376 19626
rect 24424 19574 24448 19626
rect 24448 19574 24480 19626
rect 24528 19574 24572 19626
rect 24572 19574 24584 19626
rect 24320 19572 24376 19574
rect 24424 19572 24480 19574
rect 24528 19572 24584 19574
rect 24632 19626 24688 19628
rect 24736 19626 24792 19628
rect 24840 19626 24896 19628
rect 24632 19574 24644 19626
rect 24644 19574 24688 19626
rect 24736 19574 24768 19626
rect 24768 19574 24792 19626
rect 24840 19574 24892 19626
rect 24892 19574 24896 19626
rect 24632 19572 24688 19574
rect 24736 19572 24792 19574
rect 24840 19572 24896 19574
rect 24944 19572 25000 19628
rect 25048 19626 25104 19628
rect 25152 19626 25208 19628
rect 25048 19574 25068 19626
rect 25068 19574 25104 19626
rect 25152 19574 25192 19626
rect 25192 19574 25208 19626
rect 25048 19572 25104 19574
rect 25152 19572 25208 19574
rect 14008 18842 14064 18844
rect 14112 18842 14168 18844
rect 14008 18790 14024 18842
rect 14024 18790 14064 18842
rect 14112 18790 14148 18842
rect 14148 18790 14168 18842
rect 14008 18788 14064 18790
rect 14112 18788 14168 18790
rect 14216 18788 14272 18844
rect 14320 18842 14376 18844
rect 14424 18842 14480 18844
rect 14528 18842 14584 18844
rect 14320 18790 14324 18842
rect 14324 18790 14376 18842
rect 14424 18790 14448 18842
rect 14448 18790 14480 18842
rect 14528 18790 14572 18842
rect 14572 18790 14584 18842
rect 14320 18788 14376 18790
rect 14424 18788 14480 18790
rect 14528 18788 14584 18790
rect 14632 18842 14688 18844
rect 14736 18842 14792 18844
rect 14840 18842 14896 18844
rect 14632 18790 14644 18842
rect 14644 18790 14688 18842
rect 14736 18790 14768 18842
rect 14768 18790 14792 18842
rect 14840 18790 14892 18842
rect 14892 18790 14896 18842
rect 14632 18788 14688 18790
rect 14736 18788 14792 18790
rect 14840 18788 14896 18790
rect 14944 18788 15000 18844
rect 15048 18842 15104 18844
rect 15152 18842 15208 18844
rect 15048 18790 15068 18842
rect 15068 18790 15104 18842
rect 15152 18790 15192 18842
rect 15192 18790 15208 18842
rect 15048 18788 15104 18790
rect 15152 18788 15208 18790
rect 24008 18058 24064 18060
rect 24112 18058 24168 18060
rect 24008 18006 24024 18058
rect 24024 18006 24064 18058
rect 24112 18006 24148 18058
rect 24148 18006 24168 18058
rect 24008 18004 24064 18006
rect 24112 18004 24168 18006
rect 24216 18004 24272 18060
rect 24320 18058 24376 18060
rect 24424 18058 24480 18060
rect 24528 18058 24584 18060
rect 24320 18006 24324 18058
rect 24324 18006 24376 18058
rect 24424 18006 24448 18058
rect 24448 18006 24480 18058
rect 24528 18006 24572 18058
rect 24572 18006 24584 18058
rect 24320 18004 24376 18006
rect 24424 18004 24480 18006
rect 24528 18004 24584 18006
rect 24632 18058 24688 18060
rect 24736 18058 24792 18060
rect 24840 18058 24896 18060
rect 24632 18006 24644 18058
rect 24644 18006 24688 18058
rect 24736 18006 24768 18058
rect 24768 18006 24792 18058
rect 24840 18006 24892 18058
rect 24892 18006 24896 18058
rect 24632 18004 24688 18006
rect 24736 18004 24792 18006
rect 24840 18004 24896 18006
rect 24944 18004 25000 18060
rect 25048 18058 25104 18060
rect 25152 18058 25208 18060
rect 25048 18006 25068 18058
rect 25068 18006 25104 18058
rect 25152 18006 25192 18058
rect 25192 18006 25208 18058
rect 25048 18004 25104 18006
rect 25152 18004 25208 18006
rect 14008 17274 14064 17276
rect 14112 17274 14168 17276
rect 14008 17222 14024 17274
rect 14024 17222 14064 17274
rect 14112 17222 14148 17274
rect 14148 17222 14168 17274
rect 14008 17220 14064 17222
rect 14112 17220 14168 17222
rect 14216 17220 14272 17276
rect 14320 17274 14376 17276
rect 14424 17274 14480 17276
rect 14528 17274 14584 17276
rect 14320 17222 14324 17274
rect 14324 17222 14376 17274
rect 14424 17222 14448 17274
rect 14448 17222 14480 17274
rect 14528 17222 14572 17274
rect 14572 17222 14584 17274
rect 14320 17220 14376 17222
rect 14424 17220 14480 17222
rect 14528 17220 14584 17222
rect 14632 17274 14688 17276
rect 14736 17274 14792 17276
rect 14840 17274 14896 17276
rect 14632 17222 14644 17274
rect 14644 17222 14688 17274
rect 14736 17222 14768 17274
rect 14768 17222 14792 17274
rect 14840 17222 14892 17274
rect 14892 17222 14896 17274
rect 14632 17220 14688 17222
rect 14736 17220 14792 17222
rect 14840 17220 14896 17222
rect 14944 17220 15000 17276
rect 15048 17274 15104 17276
rect 15152 17274 15208 17276
rect 15048 17222 15068 17274
rect 15068 17222 15104 17274
rect 15152 17222 15192 17274
rect 15192 17222 15208 17274
rect 15048 17220 15104 17222
rect 15152 17220 15208 17222
rect 24008 16490 24064 16492
rect 24112 16490 24168 16492
rect 24008 16438 24024 16490
rect 24024 16438 24064 16490
rect 24112 16438 24148 16490
rect 24148 16438 24168 16490
rect 24008 16436 24064 16438
rect 24112 16436 24168 16438
rect 24216 16436 24272 16492
rect 24320 16490 24376 16492
rect 24424 16490 24480 16492
rect 24528 16490 24584 16492
rect 24320 16438 24324 16490
rect 24324 16438 24376 16490
rect 24424 16438 24448 16490
rect 24448 16438 24480 16490
rect 24528 16438 24572 16490
rect 24572 16438 24584 16490
rect 24320 16436 24376 16438
rect 24424 16436 24480 16438
rect 24528 16436 24584 16438
rect 24632 16490 24688 16492
rect 24736 16490 24792 16492
rect 24840 16490 24896 16492
rect 24632 16438 24644 16490
rect 24644 16438 24688 16490
rect 24736 16438 24768 16490
rect 24768 16438 24792 16490
rect 24840 16438 24892 16490
rect 24892 16438 24896 16490
rect 24632 16436 24688 16438
rect 24736 16436 24792 16438
rect 24840 16436 24896 16438
rect 24944 16436 25000 16492
rect 25048 16490 25104 16492
rect 25152 16490 25208 16492
rect 25048 16438 25068 16490
rect 25068 16438 25104 16490
rect 25152 16438 25192 16490
rect 25192 16438 25208 16490
rect 25048 16436 25104 16438
rect 25152 16436 25208 16438
rect 14008 15706 14064 15708
rect 14112 15706 14168 15708
rect 14008 15654 14024 15706
rect 14024 15654 14064 15706
rect 14112 15654 14148 15706
rect 14148 15654 14168 15706
rect 14008 15652 14064 15654
rect 14112 15652 14168 15654
rect 14216 15652 14272 15708
rect 14320 15706 14376 15708
rect 14424 15706 14480 15708
rect 14528 15706 14584 15708
rect 14320 15654 14324 15706
rect 14324 15654 14376 15706
rect 14424 15654 14448 15706
rect 14448 15654 14480 15706
rect 14528 15654 14572 15706
rect 14572 15654 14584 15706
rect 14320 15652 14376 15654
rect 14424 15652 14480 15654
rect 14528 15652 14584 15654
rect 14632 15706 14688 15708
rect 14736 15706 14792 15708
rect 14840 15706 14896 15708
rect 14632 15654 14644 15706
rect 14644 15654 14688 15706
rect 14736 15654 14768 15706
rect 14768 15654 14792 15706
rect 14840 15654 14892 15706
rect 14892 15654 14896 15706
rect 14632 15652 14688 15654
rect 14736 15652 14792 15654
rect 14840 15652 14896 15654
rect 14944 15652 15000 15708
rect 15048 15706 15104 15708
rect 15152 15706 15208 15708
rect 15048 15654 15068 15706
rect 15068 15654 15104 15706
rect 15152 15654 15192 15706
rect 15192 15654 15208 15706
rect 15048 15652 15104 15654
rect 15152 15652 15208 15654
rect 24008 14922 24064 14924
rect 24112 14922 24168 14924
rect 24008 14870 24024 14922
rect 24024 14870 24064 14922
rect 24112 14870 24148 14922
rect 24148 14870 24168 14922
rect 24008 14868 24064 14870
rect 24112 14868 24168 14870
rect 24216 14868 24272 14924
rect 24320 14922 24376 14924
rect 24424 14922 24480 14924
rect 24528 14922 24584 14924
rect 24320 14870 24324 14922
rect 24324 14870 24376 14922
rect 24424 14870 24448 14922
rect 24448 14870 24480 14922
rect 24528 14870 24572 14922
rect 24572 14870 24584 14922
rect 24320 14868 24376 14870
rect 24424 14868 24480 14870
rect 24528 14868 24584 14870
rect 24632 14922 24688 14924
rect 24736 14922 24792 14924
rect 24840 14922 24896 14924
rect 24632 14870 24644 14922
rect 24644 14870 24688 14922
rect 24736 14870 24768 14922
rect 24768 14870 24792 14922
rect 24840 14870 24892 14922
rect 24892 14870 24896 14922
rect 24632 14868 24688 14870
rect 24736 14868 24792 14870
rect 24840 14868 24896 14870
rect 24944 14868 25000 14924
rect 25048 14922 25104 14924
rect 25152 14922 25208 14924
rect 25048 14870 25068 14922
rect 25068 14870 25104 14922
rect 25152 14870 25192 14922
rect 25192 14870 25208 14922
rect 25048 14868 25104 14870
rect 25152 14868 25208 14870
rect 14008 14138 14064 14140
rect 14112 14138 14168 14140
rect 14008 14086 14024 14138
rect 14024 14086 14064 14138
rect 14112 14086 14148 14138
rect 14148 14086 14168 14138
rect 14008 14084 14064 14086
rect 14112 14084 14168 14086
rect 14216 14084 14272 14140
rect 14320 14138 14376 14140
rect 14424 14138 14480 14140
rect 14528 14138 14584 14140
rect 14320 14086 14324 14138
rect 14324 14086 14376 14138
rect 14424 14086 14448 14138
rect 14448 14086 14480 14138
rect 14528 14086 14572 14138
rect 14572 14086 14584 14138
rect 14320 14084 14376 14086
rect 14424 14084 14480 14086
rect 14528 14084 14584 14086
rect 14632 14138 14688 14140
rect 14736 14138 14792 14140
rect 14840 14138 14896 14140
rect 14632 14086 14644 14138
rect 14644 14086 14688 14138
rect 14736 14086 14768 14138
rect 14768 14086 14792 14138
rect 14840 14086 14892 14138
rect 14892 14086 14896 14138
rect 14632 14084 14688 14086
rect 14736 14084 14792 14086
rect 14840 14084 14896 14086
rect 14944 14084 15000 14140
rect 15048 14138 15104 14140
rect 15152 14138 15208 14140
rect 15048 14086 15068 14138
rect 15068 14086 15104 14138
rect 15152 14086 15192 14138
rect 15192 14086 15208 14138
rect 15048 14084 15104 14086
rect 15152 14084 15208 14086
rect 24008 13354 24064 13356
rect 24112 13354 24168 13356
rect 24008 13302 24024 13354
rect 24024 13302 24064 13354
rect 24112 13302 24148 13354
rect 24148 13302 24168 13354
rect 24008 13300 24064 13302
rect 24112 13300 24168 13302
rect 24216 13300 24272 13356
rect 24320 13354 24376 13356
rect 24424 13354 24480 13356
rect 24528 13354 24584 13356
rect 24320 13302 24324 13354
rect 24324 13302 24376 13354
rect 24424 13302 24448 13354
rect 24448 13302 24480 13354
rect 24528 13302 24572 13354
rect 24572 13302 24584 13354
rect 24320 13300 24376 13302
rect 24424 13300 24480 13302
rect 24528 13300 24584 13302
rect 24632 13354 24688 13356
rect 24736 13354 24792 13356
rect 24840 13354 24896 13356
rect 24632 13302 24644 13354
rect 24644 13302 24688 13354
rect 24736 13302 24768 13354
rect 24768 13302 24792 13354
rect 24840 13302 24892 13354
rect 24892 13302 24896 13354
rect 24632 13300 24688 13302
rect 24736 13300 24792 13302
rect 24840 13300 24896 13302
rect 24944 13300 25000 13356
rect 25048 13354 25104 13356
rect 25152 13354 25208 13356
rect 25048 13302 25068 13354
rect 25068 13302 25104 13354
rect 25152 13302 25192 13354
rect 25192 13302 25208 13354
rect 25048 13300 25104 13302
rect 25152 13300 25208 13302
rect 14008 12570 14064 12572
rect 14112 12570 14168 12572
rect 14008 12518 14024 12570
rect 14024 12518 14064 12570
rect 14112 12518 14148 12570
rect 14148 12518 14168 12570
rect 14008 12516 14064 12518
rect 14112 12516 14168 12518
rect 14216 12516 14272 12572
rect 14320 12570 14376 12572
rect 14424 12570 14480 12572
rect 14528 12570 14584 12572
rect 14320 12518 14324 12570
rect 14324 12518 14376 12570
rect 14424 12518 14448 12570
rect 14448 12518 14480 12570
rect 14528 12518 14572 12570
rect 14572 12518 14584 12570
rect 14320 12516 14376 12518
rect 14424 12516 14480 12518
rect 14528 12516 14584 12518
rect 14632 12570 14688 12572
rect 14736 12570 14792 12572
rect 14840 12570 14896 12572
rect 14632 12518 14644 12570
rect 14644 12518 14688 12570
rect 14736 12518 14768 12570
rect 14768 12518 14792 12570
rect 14840 12518 14892 12570
rect 14892 12518 14896 12570
rect 14632 12516 14688 12518
rect 14736 12516 14792 12518
rect 14840 12516 14896 12518
rect 14944 12516 15000 12572
rect 15048 12570 15104 12572
rect 15152 12570 15208 12572
rect 15048 12518 15068 12570
rect 15068 12518 15104 12570
rect 15152 12518 15192 12570
rect 15192 12518 15208 12570
rect 15048 12516 15104 12518
rect 15152 12516 15208 12518
rect 24008 11786 24064 11788
rect 24112 11786 24168 11788
rect 24008 11734 24024 11786
rect 24024 11734 24064 11786
rect 24112 11734 24148 11786
rect 24148 11734 24168 11786
rect 24008 11732 24064 11734
rect 24112 11732 24168 11734
rect 24216 11732 24272 11788
rect 24320 11786 24376 11788
rect 24424 11786 24480 11788
rect 24528 11786 24584 11788
rect 24320 11734 24324 11786
rect 24324 11734 24376 11786
rect 24424 11734 24448 11786
rect 24448 11734 24480 11786
rect 24528 11734 24572 11786
rect 24572 11734 24584 11786
rect 24320 11732 24376 11734
rect 24424 11732 24480 11734
rect 24528 11732 24584 11734
rect 24632 11786 24688 11788
rect 24736 11786 24792 11788
rect 24840 11786 24896 11788
rect 24632 11734 24644 11786
rect 24644 11734 24688 11786
rect 24736 11734 24768 11786
rect 24768 11734 24792 11786
rect 24840 11734 24892 11786
rect 24892 11734 24896 11786
rect 24632 11732 24688 11734
rect 24736 11732 24792 11734
rect 24840 11732 24896 11734
rect 24944 11732 25000 11788
rect 25048 11786 25104 11788
rect 25152 11786 25208 11788
rect 25048 11734 25068 11786
rect 25068 11734 25104 11786
rect 25152 11734 25192 11786
rect 25192 11734 25208 11786
rect 25048 11732 25104 11734
rect 25152 11732 25208 11734
rect 14008 11002 14064 11004
rect 14112 11002 14168 11004
rect 14008 10950 14024 11002
rect 14024 10950 14064 11002
rect 14112 10950 14148 11002
rect 14148 10950 14168 11002
rect 14008 10948 14064 10950
rect 14112 10948 14168 10950
rect 14216 10948 14272 11004
rect 14320 11002 14376 11004
rect 14424 11002 14480 11004
rect 14528 11002 14584 11004
rect 14320 10950 14324 11002
rect 14324 10950 14376 11002
rect 14424 10950 14448 11002
rect 14448 10950 14480 11002
rect 14528 10950 14572 11002
rect 14572 10950 14584 11002
rect 14320 10948 14376 10950
rect 14424 10948 14480 10950
rect 14528 10948 14584 10950
rect 14632 11002 14688 11004
rect 14736 11002 14792 11004
rect 14840 11002 14896 11004
rect 14632 10950 14644 11002
rect 14644 10950 14688 11002
rect 14736 10950 14768 11002
rect 14768 10950 14792 11002
rect 14840 10950 14892 11002
rect 14892 10950 14896 11002
rect 14632 10948 14688 10950
rect 14736 10948 14792 10950
rect 14840 10948 14896 10950
rect 14944 10948 15000 11004
rect 15048 11002 15104 11004
rect 15152 11002 15208 11004
rect 15048 10950 15068 11002
rect 15068 10950 15104 11002
rect 15152 10950 15192 11002
rect 15192 10950 15208 11002
rect 15048 10948 15104 10950
rect 15152 10948 15208 10950
rect 24008 10218 24064 10220
rect 24112 10218 24168 10220
rect 24008 10166 24024 10218
rect 24024 10166 24064 10218
rect 24112 10166 24148 10218
rect 24148 10166 24168 10218
rect 24008 10164 24064 10166
rect 24112 10164 24168 10166
rect 24216 10164 24272 10220
rect 24320 10218 24376 10220
rect 24424 10218 24480 10220
rect 24528 10218 24584 10220
rect 24320 10166 24324 10218
rect 24324 10166 24376 10218
rect 24424 10166 24448 10218
rect 24448 10166 24480 10218
rect 24528 10166 24572 10218
rect 24572 10166 24584 10218
rect 24320 10164 24376 10166
rect 24424 10164 24480 10166
rect 24528 10164 24584 10166
rect 24632 10218 24688 10220
rect 24736 10218 24792 10220
rect 24840 10218 24896 10220
rect 24632 10166 24644 10218
rect 24644 10166 24688 10218
rect 24736 10166 24768 10218
rect 24768 10166 24792 10218
rect 24840 10166 24892 10218
rect 24892 10166 24896 10218
rect 24632 10164 24688 10166
rect 24736 10164 24792 10166
rect 24840 10164 24896 10166
rect 24944 10164 25000 10220
rect 25048 10218 25104 10220
rect 25152 10218 25208 10220
rect 25048 10166 25068 10218
rect 25068 10166 25104 10218
rect 25152 10166 25192 10218
rect 25192 10166 25208 10218
rect 25048 10164 25104 10166
rect 25152 10164 25208 10166
rect 14008 9434 14064 9436
rect 14112 9434 14168 9436
rect 14008 9382 14024 9434
rect 14024 9382 14064 9434
rect 14112 9382 14148 9434
rect 14148 9382 14168 9434
rect 14008 9380 14064 9382
rect 14112 9380 14168 9382
rect 14216 9380 14272 9436
rect 14320 9434 14376 9436
rect 14424 9434 14480 9436
rect 14528 9434 14584 9436
rect 14320 9382 14324 9434
rect 14324 9382 14376 9434
rect 14424 9382 14448 9434
rect 14448 9382 14480 9434
rect 14528 9382 14572 9434
rect 14572 9382 14584 9434
rect 14320 9380 14376 9382
rect 14424 9380 14480 9382
rect 14528 9380 14584 9382
rect 14632 9434 14688 9436
rect 14736 9434 14792 9436
rect 14840 9434 14896 9436
rect 14632 9382 14644 9434
rect 14644 9382 14688 9434
rect 14736 9382 14768 9434
rect 14768 9382 14792 9434
rect 14840 9382 14892 9434
rect 14892 9382 14896 9434
rect 14632 9380 14688 9382
rect 14736 9380 14792 9382
rect 14840 9380 14896 9382
rect 14944 9380 15000 9436
rect 15048 9434 15104 9436
rect 15152 9434 15208 9436
rect 15048 9382 15068 9434
rect 15068 9382 15104 9434
rect 15152 9382 15192 9434
rect 15192 9382 15208 9434
rect 15048 9380 15104 9382
rect 15152 9380 15208 9382
rect 24008 8650 24064 8652
rect 24112 8650 24168 8652
rect 24008 8598 24024 8650
rect 24024 8598 24064 8650
rect 24112 8598 24148 8650
rect 24148 8598 24168 8650
rect 24008 8596 24064 8598
rect 24112 8596 24168 8598
rect 24216 8596 24272 8652
rect 24320 8650 24376 8652
rect 24424 8650 24480 8652
rect 24528 8650 24584 8652
rect 24320 8598 24324 8650
rect 24324 8598 24376 8650
rect 24424 8598 24448 8650
rect 24448 8598 24480 8650
rect 24528 8598 24572 8650
rect 24572 8598 24584 8650
rect 24320 8596 24376 8598
rect 24424 8596 24480 8598
rect 24528 8596 24584 8598
rect 24632 8650 24688 8652
rect 24736 8650 24792 8652
rect 24840 8650 24896 8652
rect 24632 8598 24644 8650
rect 24644 8598 24688 8650
rect 24736 8598 24768 8650
rect 24768 8598 24792 8650
rect 24840 8598 24892 8650
rect 24892 8598 24896 8650
rect 24632 8596 24688 8598
rect 24736 8596 24792 8598
rect 24840 8596 24896 8598
rect 24944 8596 25000 8652
rect 25048 8650 25104 8652
rect 25152 8650 25208 8652
rect 25048 8598 25068 8650
rect 25068 8598 25104 8650
rect 25152 8598 25192 8650
rect 25192 8598 25208 8650
rect 25048 8596 25104 8598
rect 25152 8596 25208 8598
rect 14252 8146 14308 8148
rect 14252 8094 14254 8146
rect 14254 8094 14306 8146
rect 14306 8094 14308 8146
rect 14252 8092 14308 8094
rect 16492 8034 16548 8036
rect 16492 7982 16494 8034
rect 16494 7982 16546 8034
rect 16546 7982 16548 8034
rect 16492 7980 16548 7982
rect 34008 45498 34064 45500
rect 34112 45498 34168 45500
rect 34008 45446 34024 45498
rect 34024 45446 34064 45498
rect 34112 45446 34148 45498
rect 34148 45446 34168 45498
rect 34008 45444 34064 45446
rect 34112 45444 34168 45446
rect 34216 45444 34272 45500
rect 34320 45498 34376 45500
rect 34424 45498 34480 45500
rect 34528 45498 34584 45500
rect 34320 45446 34324 45498
rect 34324 45446 34376 45498
rect 34424 45446 34448 45498
rect 34448 45446 34480 45498
rect 34528 45446 34572 45498
rect 34572 45446 34584 45498
rect 34320 45444 34376 45446
rect 34424 45444 34480 45446
rect 34528 45444 34584 45446
rect 34632 45498 34688 45500
rect 34736 45498 34792 45500
rect 34840 45498 34896 45500
rect 34632 45446 34644 45498
rect 34644 45446 34688 45498
rect 34736 45446 34768 45498
rect 34768 45446 34792 45498
rect 34840 45446 34892 45498
rect 34892 45446 34896 45498
rect 34632 45444 34688 45446
rect 34736 45444 34792 45446
rect 34840 45444 34896 45446
rect 34944 45444 35000 45500
rect 35048 45498 35104 45500
rect 35152 45498 35208 45500
rect 35048 45446 35068 45498
rect 35068 45446 35104 45498
rect 35152 45446 35192 45498
rect 35192 45446 35208 45498
rect 35048 45444 35104 45446
rect 35152 45444 35208 45446
rect 34008 43930 34064 43932
rect 34112 43930 34168 43932
rect 34008 43878 34024 43930
rect 34024 43878 34064 43930
rect 34112 43878 34148 43930
rect 34148 43878 34168 43930
rect 34008 43876 34064 43878
rect 34112 43876 34168 43878
rect 34216 43876 34272 43932
rect 34320 43930 34376 43932
rect 34424 43930 34480 43932
rect 34528 43930 34584 43932
rect 34320 43878 34324 43930
rect 34324 43878 34376 43930
rect 34424 43878 34448 43930
rect 34448 43878 34480 43930
rect 34528 43878 34572 43930
rect 34572 43878 34584 43930
rect 34320 43876 34376 43878
rect 34424 43876 34480 43878
rect 34528 43876 34584 43878
rect 34632 43930 34688 43932
rect 34736 43930 34792 43932
rect 34840 43930 34896 43932
rect 34632 43878 34644 43930
rect 34644 43878 34688 43930
rect 34736 43878 34768 43930
rect 34768 43878 34792 43930
rect 34840 43878 34892 43930
rect 34892 43878 34896 43930
rect 34632 43876 34688 43878
rect 34736 43876 34792 43878
rect 34840 43876 34896 43878
rect 34944 43876 35000 43932
rect 35048 43930 35104 43932
rect 35152 43930 35208 43932
rect 35048 43878 35068 43930
rect 35068 43878 35104 43930
rect 35152 43878 35192 43930
rect 35192 43878 35208 43930
rect 35048 43876 35104 43878
rect 35152 43876 35208 43878
rect 34008 42362 34064 42364
rect 34112 42362 34168 42364
rect 34008 42310 34024 42362
rect 34024 42310 34064 42362
rect 34112 42310 34148 42362
rect 34148 42310 34168 42362
rect 34008 42308 34064 42310
rect 34112 42308 34168 42310
rect 34216 42308 34272 42364
rect 34320 42362 34376 42364
rect 34424 42362 34480 42364
rect 34528 42362 34584 42364
rect 34320 42310 34324 42362
rect 34324 42310 34376 42362
rect 34424 42310 34448 42362
rect 34448 42310 34480 42362
rect 34528 42310 34572 42362
rect 34572 42310 34584 42362
rect 34320 42308 34376 42310
rect 34424 42308 34480 42310
rect 34528 42308 34584 42310
rect 34632 42362 34688 42364
rect 34736 42362 34792 42364
rect 34840 42362 34896 42364
rect 34632 42310 34644 42362
rect 34644 42310 34688 42362
rect 34736 42310 34768 42362
rect 34768 42310 34792 42362
rect 34840 42310 34892 42362
rect 34892 42310 34896 42362
rect 34632 42308 34688 42310
rect 34736 42308 34792 42310
rect 34840 42308 34896 42310
rect 34944 42308 35000 42364
rect 35048 42362 35104 42364
rect 35152 42362 35208 42364
rect 35048 42310 35068 42362
rect 35068 42310 35104 42362
rect 35152 42310 35192 42362
rect 35192 42310 35208 42362
rect 35048 42308 35104 42310
rect 35152 42308 35208 42310
rect 34008 40794 34064 40796
rect 34112 40794 34168 40796
rect 34008 40742 34024 40794
rect 34024 40742 34064 40794
rect 34112 40742 34148 40794
rect 34148 40742 34168 40794
rect 34008 40740 34064 40742
rect 34112 40740 34168 40742
rect 34216 40740 34272 40796
rect 34320 40794 34376 40796
rect 34424 40794 34480 40796
rect 34528 40794 34584 40796
rect 34320 40742 34324 40794
rect 34324 40742 34376 40794
rect 34424 40742 34448 40794
rect 34448 40742 34480 40794
rect 34528 40742 34572 40794
rect 34572 40742 34584 40794
rect 34320 40740 34376 40742
rect 34424 40740 34480 40742
rect 34528 40740 34584 40742
rect 34632 40794 34688 40796
rect 34736 40794 34792 40796
rect 34840 40794 34896 40796
rect 34632 40742 34644 40794
rect 34644 40742 34688 40794
rect 34736 40742 34768 40794
rect 34768 40742 34792 40794
rect 34840 40742 34892 40794
rect 34892 40742 34896 40794
rect 34632 40740 34688 40742
rect 34736 40740 34792 40742
rect 34840 40740 34896 40742
rect 34944 40740 35000 40796
rect 35048 40794 35104 40796
rect 35152 40794 35208 40796
rect 35048 40742 35068 40794
rect 35068 40742 35104 40794
rect 35152 40742 35192 40794
rect 35192 40742 35208 40794
rect 35048 40740 35104 40742
rect 35152 40740 35208 40742
rect 34008 39226 34064 39228
rect 34112 39226 34168 39228
rect 34008 39174 34024 39226
rect 34024 39174 34064 39226
rect 34112 39174 34148 39226
rect 34148 39174 34168 39226
rect 34008 39172 34064 39174
rect 34112 39172 34168 39174
rect 34216 39172 34272 39228
rect 34320 39226 34376 39228
rect 34424 39226 34480 39228
rect 34528 39226 34584 39228
rect 34320 39174 34324 39226
rect 34324 39174 34376 39226
rect 34424 39174 34448 39226
rect 34448 39174 34480 39226
rect 34528 39174 34572 39226
rect 34572 39174 34584 39226
rect 34320 39172 34376 39174
rect 34424 39172 34480 39174
rect 34528 39172 34584 39174
rect 34632 39226 34688 39228
rect 34736 39226 34792 39228
rect 34840 39226 34896 39228
rect 34632 39174 34644 39226
rect 34644 39174 34688 39226
rect 34736 39174 34768 39226
rect 34768 39174 34792 39226
rect 34840 39174 34892 39226
rect 34892 39174 34896 39226
rect 34632 39172 34688 39174
rect 34736 39172 34792 39174
rect 34840 39172 34896 39174
rect 34944 39172 35000 39228
rect 35048 39226 35104 39228
rect 35152 39226 35208 39228
rect 35048 39174 35068 39226
rect 35068 39174 35104 39226
rect 35152 39174 35192 39226
rect 35192 39174 35208 39226
rect 35048 39172 35104 39174
rect 35152 39172 35208 39174
rect 34008 37658 34064 37660
rect 34112 37658 34168 37660
rect 34008 37606 34024 37658
rect 34024 37606 34064 37658
rect 34112 37606 34148 37658
rect 34148 37606 34168 37658
rect 34008 37604 34064 37606
rect 34112 37604 34168 37606
rect 34216 37604 34272 37660
rect 34320 37658 34376 37660
rect 34424 37658 34480 37660
rect 34528 37658 34584 37660
rect 34320 37606 34324 37658
rect 34324 37606 34376 37658
rect 34424 37606 34448 37658
rect 34448 37606 34480 37658
rect 34528 37606 34572 37658
rect 34572 37606 34584 37658
rect 34320 37604 34376 37606
rect 34424 37604 34480 37606
rect 34528 37604 34584 37606
rect 34632 37658 34688 37660
rect 34736 37658 34792 37660
rect 34840 37658 34896 37660
rect 34632 37606 34644 37658
rect 34644 37606 34688 37658
rect 34736 37606 34768 37658
rect 34768 37606 34792 37658
rect 34840 37606 34892 37658
rect 34892 37606 34896 37658
rect 34632 37604 34688 37606
rect 34736 37604 34792 37606
rect 34840 37604 34896 37606
rect 34944 37604 35000 37660
rect 35048 37658 35104 37660
rect 35152 37658 35208 37660
rect 35048 37606 35068 37658
rect 35068 37606 35104 37658
rect 35152 37606 35192 37658
rect 35192 37606 35208 37658
rect 35048 37604 35104 37606
rect 35152 37604 35208 37606
rect 34008 36090 34064 36092
rect 34112 36090 34168 36092
rect 34008 36038 34024 36090
rect 34024 36038 34064 36090
rect 34112 36038 34148 36090
rect 34148 36038 34168 36090
rect 34008 36036 34064 36038
rect 34112 36036 34168 36038
rect 34216 36036 34272 36092
rect 34320 36090 34376 36092
rect 34424 36090 34480 36092
rect 34528 36090 34584 36092
rect 34320 36038 34324 36090
rect 34324 36038 34376 36090
rect 34424 36038 34448 36090
rect 34448 36038 34480 36090
rect 34528 36038 34572 36090
rect 34572 36038 34584 36090
rect 34320 36036 34376 36038
rect 34424 36036 34480 36038
rect 34528 36036 34584 36038
rect 34632 36090 34688 36092
rect 34736 36090 34792 36092
rect 34840 36090 34896 36092
rect 34632 36038 34644 36090
rect 34644 36038 34688 36090
rect 34736 36038 34768 36090
rect 34768 36038 34792 36090
rect 34840 36038 34892 36090
rect 34892 36038 34896 36090
rect 34632 36036 34688 36038
rect 34736 36036 34792 36038
rect 34840 36036 34896 36038
rect 34944 36036 35000 36092
rect 35048 36090 35104 36092
rect 35152 36090 35208 36092
rect 35048 36038 35068 36090
rect 35068 36038 35104 36090
rect 35152 36038 35192 36090
rect 35192 36038 35208 36090
rect 35048 36036 35104 36038
rect 35152 36036 35208 36038
rect 34008 34522 34064 34524
rect 34112 34522 34168 34524
rect 34008 34470 34024 34522
rect 34024 34470 34064 34522
rect 34112 34470 34148 34522
rect 34148 34470 34168 34522
rect 34008 34468 34064 34470
rect 34112 34468 34168 34470
rect 34216 34468 34272 34524
rect 34320 34522 34376 34524
rect 34424 34522 34480 34524
rect 34528 34522 34584 34524
rect 34320 34470 34324 34522
rect 34324 34470 34376 34522
rect 34424 34470 34448 34522
rect 34448 34470 34480 34522
rect 34528 34470 34572 34522
rect 34572 34470 34584 34522
rect 34320 34468 34376 34470
rect 34424 34468 34480 34470
rect 34528 34468 34584 34470
rect 34632 34522 34688 34524
rect 34736 34522 34792 34524
rect 34840 34522 34896 34524
rect 34632 34470 34644 34522
rect 34644 34470 34688 34522
rect 34736 34470 34768 34522
rect 34768 34470 34792 34522
rect 34840 34470 34892 34522
rect 34892 34470 34896 34522
rect 34632 34468 34688 34470
rect 34736 34468 34792 34470
rect 34840 34468 34896 34470
rect 34944 34468 35000 34524
rect 35048 34522 35104 34524
rect 35152 34522 35208 34524
rect 35048 34470 35068 34522
rect 35068 34470 35104 34522
rect 35152 34470 35192 34522
rect 35192 34470 35208 34522
rect 35048 34468 35104 34470
rect 35152 34468 35208 34470
rect 34008 32954 34064 32956
rect 34112 32954 34168 32956
rect 34008 32902 34024 32954
rect 34024 32902 34064 32954
rect 34112 32902 34148 32954
rect 34148 32902 34168 32954
rect 34008 32900 34064 32902
rect 34112 32900 34168 32902
rect 34216 32900 34272 32956
rect 34320 32954 34376 32956
rect 34424 32954 34480 32956
rect 34528 32954 34584 32956
rect 34320 32902 34324 32954
rect 34324 32902 34376 32954
rect 34424 32902 34448 32954
rect 34448 32902 34480 32954
rect 34528 32902 34572 32954
rect 34572 32902 34584 32954
rect 34320 32900 34376 32902
rect 34424 32900 34480 32902
rect 34528 32900 34584 32902
rect 34632 32954 34688 32956
rect 34736 32954 34792 32956
rect 34840 32954 34896 32956
rect 34632 32902 34644 32954
rect 34644 32902 34688 32954
rect 34736 32902 34768 32954
rect 34768 32902 34792 32954
rect 34840 32902 34892 32954
rect 34892 32902 34896 32954
rect 34632 32900 34688 32902
rect 34736 32900 34792 32902
rect 34840 32900 34896 32902
rect 34944 32900 35000 32956
rect 35048 32954 35104 32956
rect 35152 32954 35208 32956
rect 35048 32902 35068 32954
rect 35068 32902 35104 32954
rect 35152 32902 35192 32954
rect 35192 32902 35208 32954
rect 35048 32900 35104 32902
rect 35152 32900 35208 32902
rect 34008 31386 34064 31388
rect 34112 31386 34168 31388
rect 34008 31334 34024 31386
rect 34024 31334 34064 31386
rect 34112 31334 34148 31386
rect 34148 31334 34168 31386
rect 34008 31332 34064 31334
rect 34112 31332 34168 31334
rect 34216 31332 34272 31388
rect 34320 31386 34376 31388
rect 34424 31386 34480 31388
rect 34528 31386 34584 31388
rect 34320 31334 34324 31386
rect 34324 31334 34376 31386
rect 34424 31334 34448 31386
rect 34448 31334 34480 31386
rect 34528 31334 34572 31386
rect 34572 31334 34584 31386
rect 34320 31332 34376 31334
rect 34424 31332 34480 31334
rect 34528 31332 34584 31334
rect 34632 31386 34688 31388
rect 34736 31386 34792 31388
rect 34840 31386 34896 31388
rect 34632 31334 34644 31386
rect 34644 31334 34688 31386
rect 34736 31334 34768 31386
rect 34768 31334 34792 31386
rect 34840 31334 34892 31386
rect 34892 31334 34896 31386
rect 34632 31332 34688 31334
rect 34736 31332 34792 31334
rect 34840 31332 34896 31334
rect 34944 31332 35000 31388
rect 35048 31386 35104 31388
rect 35152 31386 35208 31388
rect 35048 31334 35068 31386
rect 35068 31334 35104 31386
rect 35152 31334 35192 31386
rect 35192 31334 35208 31386
rect 35048 31332 35104 31334
rect 35152 31332 35208 31334
rect 34008 29818 34064 29820
rect 34112 29818 34168 29820
rect 34008 29766 34024 29818
rect 34024 29766 34064 29818
rect 34112 29766 34148 29818
rect 34148 29766 34168 29818
rect 34008 29764 34064 29766
rect 34112 29764 34168 29766
rect 34216 29764 34272 29820
rect 34320 29818 34376 29820
rect 34424 29818 34480 29820
rect 34528 29818 34584 29820
rect 34320 29766 34324 29818
rect 34324 29766 34376 29818
rect 34424 29766 34448 29818
rect 34448 29766 34480 29818
rect 34528 29766 34572 29818
rect 34572 29766 34584 29818
rect 34320 29764 34376 29766
rect 34424 29764 34480 29766
rect 34528 29764 34584 29766
rect 34632 29818 34688 29820
rect 34736 29818 34792 29820
rect 34840 29818 34896 29820
rect 34632 29766 34644 29818
rect 34644 29766 34688 29818
rect 34736 29766 34768 29818
rect 34768 29766 34792 29818
rect 34840 29766 34892 29818
rect 34892 29766 34896 29818
rect 34632 29764 34688 29766
rect 34736 29764 34792 29766
rect 34840 29764 34896 29766
rect 34944 29764 35000 29820
rect 35048 29818 35104 29820
rect 35152 29818 35208 29820
rect 35048 29766 35068 29818
rect 35068 29766 35104 29818
rect 35152 29766 35192 29818
rect 35192 29766 35208 29818
rect 35048 29764 35104 29766
rect 35152 29764 35208 29766
rect 34008 28250 34064 28252
rect 34112 28250 34168 28252
rect 34008 28198 34024 28250
rect 34024 28198 34064 28250
rect 34112 28198 34148 28250
rect 34148 28198 34168 28250
rect 34008 28196 34064 28198
rect 34112 28196 34168 28198
rect 34216 28196 34272 28252
rect 34320 28250 34376 28252
rect 34424 28250 34480 28252
rect 34528 28250 34584 28252
rect 34320 28198 34324 28250
rect 34324 28198 34376 28250
rect 34424 28198 34448 28250
rect 34448 28198 34480 28250
rect 34528 28198 34572 28250
rect 34572 28198 34584 28250
rect 34320 28196 34376 28198
rect 34424 28196 34480 28198
rect 34528 28196 34584 28198
rect 34632 28250 34688 28252
rect 34736 28250 34792 28252
rect 34840 28250 34896 28252
rect 34632 28198 34644 28250
rect 34644 28198 34688 28250
rect 34736 28198 34768 28250
rect 34768 28198 34792 28250
rect 34840 28198 34892 28250
rect 34892 28198 34896 28250
rect 34632 28196 34688 28198
rect 34736 28196 34792 28198
rect 34840 28196 34896 28198
rect 34944 28196 35000 28252
rect 35048 28250 35104 28252
rect 35152 28250 35208 28252
rect 35048 28198 35068 28250
rect 35068 28198 35104 28250
rect 35152 28198 35192 28250
rect 35192 28198 35208 28250
rect 35048 28196 35104 28198
rect 35152 28196 35208 28198
rect 34008 26682 34064 26684
rect 34112 26682 34168 26684
rect 34008 26630 34024 26682
rect 34024 26630 34064 26682
rect 34112 26630 34148 26682
rect 34148 26630 34168 26682
rect 34008 26628 34064 26630
rect 34112 26628 34168 26630
rect 34216 26628 34272 26684
rect 34320 26682 34376 26684
rect 34424 26682 34480 26684
rect 34528 26682 34584 26684
rect 34320 26630 34324 26682
rect 34324 26630 34376 26682
rect 34424 26630 34448 26682
rect 34448 26630 34480 26682
rect 34528 26630 34572 26682
rect 34572 26630 34584 26682
rect 34320 26628 34376 26630
rect 34424 26628 34480 26630
rect 34528 26628 34584 26630
rect 34632 26682 34688 26684
rect 34736 26682 34792 26684
rect 34840 26682 34896 26684
rect 34632 26630 34644 26682
rect 34644 26630 34688 26682
rect 34736 26630 34768 26682
rect 34768 26630 34792 26682
rect 34840 26630 34892 26682
rect 34892 26630 34896 26682
rect 34632 26628 34688 26630
rect 34736 26628 34792 26630
rect 34840 26628 34896 26630
rect 34944 26628 35000 26684
rect 35048 26682 35104 26684
rect 35152 26682 35208 26684
rect 35048 26630 35068 26682
rect 35068 26630 35104 26682
rect 35152 26630 35192 26682
rect 35192 26630 35208 26682
rect 35048 26628 35104 26630
rect 35152 26628 35208 26630
rect 34008 25114 34064 25116
rect 34112 25114 34168 25116
rect 34008 25062 34024 25114
rect 34024 25062 34064 25114
rect 34112 25062 34148 25114
rect 34148 25062 34168 25114
rect 34008 25060 34064 25062
rect 34112 25060 34168 25062
rect 34216 25060 34272 25116
rect 34320 25114 34376 25116
rect 34424 25114 34480 25116
rect 34528 25114 34584 25116
rect 34320 25062 34324 25114
rect 34324 25062 34376 25114
rect 34424 25062 34448 25114
rect 34448 25062 34480 25114
rect 34528 25062 34572 25114
rect 34572 25062 34584 25114
rect 34320 25060 34376 25062
rect 34424 25060 34480 25062
rect 34528 25060 34584 25062
rect 34632 25114 34688 25116
rect 34736 25114 34792 25116
rect 34840 25114 34896 25116
rect 34632 25062 34644 25114
rect 34644 25062 34688 25114
rect 34736 25062 34768 25114
rect 34768 25062 34792 25114
rect 34840 25062 34892 25114
rect 34892 25062 34896 25114
rect 34632 25060 34688 25062
rect 34736 25060 34792 25062
rect 34840 25060 34896 25062
rect 34944 25060 35000 25116
rect 35048 25114 35104 25116
rect 35152 25114 35208 25116
rect 35048 25062 35068 25114
rect 35068 25062 35104 25114
rect 35152 25062 35192 25114
rect 35192 25062 35208 25114
rect 35048 25060 35104 25062
rect 35152 25060 35208 25062
rect 34008 23546 34064 23548
rect 34112 23546 34168 23548
rect 34008 23494 34024 23546
rect 34024 23494 34064 23546
rect 34112 23494 34148 23546
rect 34148 23494 34168 23546
rect 34008 23492 34064 23494
rect 34112 23492 34168 23494
rect 34216 23492 34272 23548
rect 34320 23546 34376 23548
rect 34424 23546 34480 23548
rect 34528 23546 34584 23548
rect 34320 23494 34324 23546
rect 34324 23494 34376 23546
rect 34424 23494 34448 23546
rect 34448 23494 34480 23546
rect 34528 23494 34572 23546
rect 34572 23494 34584 23546
rect 34320 23492 34376 23494
rect 34424 23492 34480 23494
rect 34528 23492 34584 23494
rect 34632 23546 34688 23548
rect 34736 23546 34792 23548
rect 34840 23546 34896 23548
rect 34632 23494 34644 23546
rect 34644 23494 34688 23546
rect 34736 23494 34768 23546
rect 34768 23494 34792 23546
rect 34840 23494 34892 23546
rect 34892 23494 34896 23546
rect 34632 23492 34688 23494
rect 34736 23492 34792 23494
rect 34840 23492 34896 23494
rect 34944 23492 35000 23548
rect 35048 23546 35104 23548
rect 35152 23546 35208 23548
rect 35048 23494 35068 23546
rect 35068 23494 35104 23546
rect 35152 23494 35192 23546
rect 35192 23494 35208 23546
rect 35048 23492 35104 23494
rect 35152 23492 35208 23494
rect 34008 21978 34064 21980
rect 34112 21978 34168 21980
rect 34008 21926 34024 21978
rect 34024 21926 34064 21978
rect 34112 21926 34148 21978
rect 34148 21926 34168 21978
rect 34008 21924 34064 21926
rect 34112 21924 34168 21926
rect 34216 21924 34272 21980
rect 34320 21978 34376 21980
rect 34424 21978 34480 21980
rect 34528 21978 34584 21980
rect 34320 21926 34324 21978
rect 34324 21926 34376 21978
rect 34424 21926 34448 21978
rect 34448 21926 34480 21978
rect 34528 21926 34572 21978
rect 34572 21926 34584 21978
rect 34320 21924 34376 21926
rect 34424 21924 34480 21926
rect 34528 21924 34584 21926
rect 34632 21978 34688 21980
rect 34736 21978 34792 21980
rect 34840 21978 34896 21980
rect 34632 21926 34644 21978
rect 34644 21926 34688 21978
rect 34736 21926 34768 21978
rect 34768 21926 34792 21978
rect 34840 21926 34892 21978
rect 34892 21926 34896 21978
rect 34632 21924 34688 21926
rect 34736 21924 34792 21926
rect 34840 21924 34896 21926
rect 34944 21924 35000 21980
rect 35048 21978 35104 21980
rect 35152 21978 35208 21980
rect 35048 21926 35068 21978
rect 35068 21926 35104 21978
rect 35152 21926 35192 21978
rect 35192 21926 35208 21978
rect 35048 21924 35104 21926
rect 35152 21924 35208 21926
rect 34008 20410 34064 20412
rect 34112 20410 34168 20412
rect 34008 20358 34024 20410
rect 34024 20358 34064 20410
rect 34112 20358 34148 20410
rect 34148 20358 34168 20410
rect 34008 20356 34064 20358
rect 34112 20356 34168 20358
rect 34216 20356 34272 20412
rect 34320 20410 34376 20412
rect 34424 20410 34480 20412
rect 34528 20410 34584 20412
rect 34320 20358 34324 20410
rect 34324 20358 34376 20410
rect 34424 20358 34448 20410
rect 34448 20358 34480 20410
rect 34528 20358 34572 20410
rect 34572 20358 34584 20410
rect 34320 20356 34376 20358
rect 34424 20356 34480 20358
rect 34528 20356 34584 20358
rect 34632 20410 34688 20412
rect 34736 20410 34792 20412
rect 34840 20410 34896 20412
rect 34632 20358 34644 20410
rect 34644 20358 34688 20410
rect 34736 20358 34768 20410
rect 34768 20358 34792 20410
rect 34840 20358 34892 20410
rect 34892 20358 34896 20410
rect 34632 20356 34688 20358
rect 34736 20356 34792 20358
rect 34840 20356 34896 20358
rect 34944 20356 35000 20412
rect 35048 20410 35104 20412
rect 35152 20410 35208 20412
rect 35048 20358 35068 20410
rect 35068 20358 35104 20410
rect 35152 20358 35192 20410
rect 35192 20358 35208 20410
rect 35048 20356 35104 20358
rect 35152 20356 35208 20358
rect 34008 18842 34064 18844
rect 34112 18842 34168 18844
rect 34008 18790 34024 18842
rect 34024 18790 34064 18842
rect 34112 18790 34148 18842
rect 34148 18790 34168 18842
rect 34008 18788 34064 18790
rect 34112 18788 34168 18790
rect 34216 18788 34272 18844
rect 34320 18842 34376 18844
rect 34424 18842 34480 18844
rect 34528 18842 34584 18844
rect 34320 18790 34324 18842
rect 34324 18790 34376 18842
rect 34424 18790 34448 18842
rect 34448 18790 34480 18842
rect 34528 18790 34572 18842
rect 34572 18790 34584 18842
rect 34320 18788 34376 18790
rect 34424 18788 34480 18790
rect 34528 18788 34584 18790
rect 34632 18842 34688 18844
rect 34736 18842 34792 18844
rect 34840 18842 34896 18844
rect 34632 18790 34644 18842
rect 34644 18790 34688 18842
rect 34736 18790 34768 18842
rect 34768 18790 34792 18842
rect 34840 18790 34892 18842
rect 34892 18790 34896 18842
rect 34632 18788 34688 18790
rect 34736 18788 34792 18790
rect 34840 18788 34896 18790
rect 34944 18788 35000 18844
rect 35048 18842 35104 18844
rect 35152 18842 35208 18844
rect 35048 18790 35068 18842
rect 35068 18790 35104 18842
rect 35152 18790 35192 18842
rect 35192 18790 35208 18842
rect 35048 18788 35104 18790
rect 35152 18788 35208 18790
rect 34008 17274 34064 17276
rect 34112 17274 34168 17276
rect 34008 17222 34024 17274
rect 34024 17222 34064 17274
rect 34112 17222 34148 17274
rect 34148 17222 34168 17274
rect 34008 17220 34064 17222
rect 34112 17220 34168 17222
rect 34216 17220 34272 17276
rect 34320 17274 34376 17276
rect 34424 17274 34480 17276
rect 34528 17274 34584 17276
rect 34320 17222 34324 17274
rect 34324 17222 34376 17274
rect 34424 17222 34448 17274
rect 34448 17222 34480 17274
rect 34528 17222 34572 17274
rect 34572 17222 34584 17274
rect 34320 17220 34376 17222
rect 34424 17220 34480 17222
rect 34528 17220 34584 17222
rect 34632 17274 34688 17276
rect 34736 17274 34792 17276
rect 34840 17274 34896 17276
rect 34632 17222 34644 17274
rect 34644 17222 34688 17274
rect 34736 17222 34768 17274
rect 34768 17222 34792 17274
rect 34840 17222 34892 17274
rect 34892 17222 34896 17274
rect 34632 17220 34688 17222
rect 34736 17220 34792 17222
rect 34840 17220 34896 17222
rect 34944 17220 35000 17276
rect 35048 17274 35104 17276
rect 35152 17274 35208 17276
rect 35048 17222 35068 17274
rect 35068 17222 35104 17274
rect 35152 17222 35192 17274
rect 35192 17222 35208 17274
rect 35048 17220 35104 17222
rect 35152 17220 35208 17222
rect 34008 15706 34064 15708
rect 34112 15706 34168 15708
rect 34008 15654 34024 15706
rect 34024 15654 34064 15706
rect 34112 15654 34148 15706
rect 34148 15654 34168 15706
rect 34008 15652 34064 15654
rect 34112 15652 34168 15654
rect 34216 15652 34272 15708
rect 34320 15706 34376 15708
rect 34424 15706 34480 15708
rect 34528 15706 34584 15708
rect 34320 15654 34324 15706
rect 34324 15654 34376 15706
rect 34424 15654 34448 15706
rect 34448 15654 34480 15706
rect 34528 15654 34572 15706
rect 34572 15654 34584 15706
rect 34320 15652 34376 15654
rect 34424 15652 34480 15654
rect 34528 15652 34584 15654
rect 34632 15706 34688 15708
rect 34736 15706 34792 15708
rect 34840 15706 34896 15708
rect 34632 15654 34644 15706
rect 34644 15654 34688 15706
rect 34736 15654 34768 15706
rect 34768 15654 34792 15706
rect 34840 15654 34892 15706
rect 34892 15654 34896 15706
rect 34632 15652 34688 15654
rect 34736 15652 34792 15654
rect 34840 15652 34896 15654
rect 34944 15652 35000 15708
rect 35048 15706 35104 15708
rect 35152 15706 35208 15708
rect 35048 15654 35068 15706
rect 35068 15654 35104 15706
rect 35152 15654 35192 15706
rect 35192 15654 35208 15706
rect 35048 15652 35104 15654
rect 35152 15652 35208 15654
rect 34008 14138 34064 14140
rect 34112 14138 34168 14140
rect 34008 14086 34024 14138
rect 34024 14086 34064 14138
rect 34112 14086 34148 14138
rect 34148 14086 34168 14138
rect 34008 14084 34064 14086
rect 34112 14084 34168 14086
rect 34216 14084 34272 14140
rect 34320 14138 34376 14140
rect 34424 14138 34480 14140
rect 34528 14138 34584 14140
rect 34320 14086 34324 14138
rect 34324 14086 34376 14138
rect 34424 14086 34448 14138
rect 34448 14086 34480 14138
rect 34528 14086 34572 14138
rect 34572 14086 34584 14138
rect 34320 14084 34376 14086
rect 34424 14084 34480 14086
rect 34528 14084 34584 14086
rect 34632 14138 34688 14140
rect 34736 14138 34792 14140
rect 34840 14138 34896 14140
rect 34632 14086 34644 14138
rect 34644 14086 34688 14138
rect 34736 14086 34768 14138
rect 34768 14086 34792 14138
rect 34840 14086 34892 14138
rect 34892 14086 34896 14138
rect 34632 14084 34688 14086
rect 34736 14084 34792 14086
rect 34840 14084 34896 14086
rect 34944 14084 35000 14140
rect 35048 14138 35104 14140
rect 35152 14138 35208 14140
rect 35048 14086 35068 14138
rect 35068 14086 35104 14138
rect 35152 14086 35192 14138
rect 35192 14086 35208 14138
rect 35048 14084 35104 14086
rect 35152 14084 35208 14086
rect 34008 12570 34064 12572
rect 34112 12570 34168 12572
rect 34008 12518 34024 12570
rect 34024 12518 34064 12570
rect 34112 12518 34148 12570
rect 34148 12518 34168 12570
rect 34008 12516 34064 12518
rect 34112 12516 34168 12518
rect 34216 12516 34272 12572
rect 34320 12570 34376 12572
rect 34424 12570 34480 12572
rect 34528 12570 34584 12572
rect 34320 12518 34324 12570
rect 34324 12518 34376 12570
rect 34424 12518 34448 12570
rect 34448 12518 34480 12570
rect 34528 12518 34572 12570
rect 34572 12518 34584 12570
rect 34320 12516 34376 12518
rect 34424 12516 34480 12518
rect 34528 12516 34584 12518
rect 34632 12570 34688 12572
rect 34736 12570 34792 12572
rect 34840 12570 34896 12572
rect 34632 12518 34644 12570
rect 34644 12518 34688 12570
rect 34736 12518 34768 12570
rect 34768 12518 34792 12570
rect 34840 12518 34892 12570
rect 34892 12518 34896 12570
rect 34632 12516 34688 12518
rect 34736 12516 34792 12518
rect 34840 12516 34896 12518
rect 34944 12516 35000 12572
rect 35048 12570 35104 12572
rect 35152 12570 35208 12572
rect 35048 12518 35068 12570
rect 35068 12518 35104 12570
rect 35152 12518 35192 12570
rect 35192 12518 35208 12570
rect 35048 12516 35104 12518
rect 35152 12516 35208 12518
rect 34008 11002 34064 11004
rect 34112 11002 34168 11004
rect 34008 10950 34024 11002
rect 34024 10950 34064 11002
rect 34112 10950 34148 11002
rect 34148 10950 34168 11002
rect 34008 10948 34064 10950
rect 34112 10948 34168 10950
rect 34216 10948 34272 11004
rect 34320 11002 34376 11004
rect 34424 11002 34480 11004
rect 34528 11002 34584 11004
rect 34320 10950 34324 11002
rect 34324 10950 34376 11002
rect 34424 10950 34448 11002
rect 34448 10950 34480 11002
rect 34528 10950 34572 11002
rect 34572 10950 34584 11002
rect 34320 10948 34376 10950
rect 34424 10948 34480 10950
rect 34528 10948 34584 10950
rect 34632 11002 34688 11004
rect 34736 11002 34792 11004
rect 34840 11002 34896 11004
rect 34632 10950 34644 11002
rect 34644 10950 34688 11002
rect 34736 10950 34768 11002
rect 34768 10950 34792 11002
rect 34840 10950 34892 11002
rect 34892 10950 34896 11002
rect 34632 10948 34688 10950
rect 34736 10948 34792 10950
rect 34840 10948 34896 10950
rect 34944 10948 35000 11004
rect 35048 11002 35104 11004
rect 35152 11002 35208 11004
rect 35048 10950 35068 11002
rect 35068 10950 35104 11002
rect 35152 10950 35192 11002
rect 35192 10950 35208 11002
rect 35048 10948 35104 10950
rect 35152 10948 35208 10950
rect 38220 43314 38276 43316
rect 38220 43262 38222 43314
rect 38222 43262 38274 43314
rect 38274 43262 38276 43314
rect 38220 43260 38276 43262
rect 37660 31554 37716 31556
rect 37660 31502 37662 31554
rect 37662 31502 37714 31554
rect 37714 31502 37716 31554
rect 37660 31500 37716 31502
rect 37436 10444 37492 10500
rect 38220 31554 38276 31556
rect 38220 31502 38222 31554
rect 38222 31502 38274 31554
rect 38274 31502 38276 31554
rect 38220 31500 38276 31502
rect 38220 30940 38276 30996
rect 38220 18620 38276 18676
rect 37884 9660 37940 9716
rect 34008 9434 34064 9436
rect 34112 9434 34168 9436
rect 34008 9382 34024 9434
rect 34024 9382 34064 9434
rect 34112 9382 34148 9434
rect 34148 9382 34168 9434
rect 34008 9380 34064 9382
rect 34112 9380 34168 9382
rect 34216 9380 34272 9436
rect 34320 9434 34376 9436
rect 34424 9434 34480 9436
rect 34528 9434 34584 9436
rect 34320 9382 34324 9434
rect 34324 9382 34376 9434
rect 34424 9382 34448 9434
rect 34448 9382 34480 9434
rect 34528 9382 34572 9434
rect 34572 9382 34584 9434
rect 34320 9380 34376 9382
rect 34424 9380 34480 9382
rect 34528 9380 34584 9382
rect 34632 9434 34688 9436
rect 34736 9434 34792 9436
rect 34840 9434 34896 9436
rect 34632 9382 34644 9434
rect 34644 9382 34688 9434
rect 34736 9382 34768 9434
rect 34768 9382 34792 9434
rect 34840 9382 34892 9434
rect 34892 9382 34896 9434
rect 34632 9380 34688 9382
rect 34736 9380 34792 9382
rect 34840 9380 34896 9382
rect 34944 9380 35000 9436
rect 35048 9434 35104 9436
rect 35152 9434 35208 9436
rect 35048 9382 35068 9434
rect 35068 9382 35104 9434
rect 35152 9382 35192 9434
rect 35192 9382 35208 9434
rect 35048 9380 35104 9382
rect 35152 9380 35208 9382
rect 28364 7980 28420 8036
rect 37884 8316 37940 8372
rect 14008 7866 14064 7868
rect 14112 7866 14168 7868
rect 14008 7814 14024 7866
rect 14024 7814 14064 7866
rect 14112 7814 14148 7866
rect 14148 7814 14168 7866
rect 14008 7812 14064 7814
rect 14112 7812 14168 7814
rect 14216 7812 14272 7868
rect 14320 7866 14376 7868
rect 14424 7866 14480 7868
rect 14528 7866 14584 7868
rect 14320 7814 14324 7866
rect 14324 7814 14376 7866
rect 14424 7814 14448 7866
rect 14448 7814 14480 7866
rect 14528 7814 14572 7866
rect 14572 7814 14584 7866
rect 14320 7812 14376 7814
rect 14424 7812 14480 7814
rect 14528 7812 14584 7814
rect 14632 7866 14688 7868
rect 14736 7866 14792 7868
rect 14840 7866 14896 7868
rect 14632 7814 14644 7866
rect 14644 7814 14688 7866
rect 14736 7814 14768 7866
rect 14768 7814 14792 7866
rect 14840 7814 14892 7866
rect 14892 7814 14896 7866
rect 14632 7812 14688 7814
rect 14736 7812 14792 7814
rect 14840 7812 14896 7814
rect 14944 7812 15000 7868
rect 15048 7866 15104 7868
rect 15152 7866 15208 7868
rect 15048 7814 15068 7866
rect 15068 7814 15104 7866
rect 15152 7814 15192 7866
rect 15192 7814 15208 7866
rect 15048 7812 15104 7814
rect 15152 7812 15208 7814
rect 34008 7866 34064 7868
rect 34112 7866 34168 7868
rect 34008 7814 34024 7866
rect 34024 7814 34064 7866
rect 34112 7814 34148 7866
rect 34148 7814 34168 7866
rect 34008 7812 34064 7814
rect 34112 7812 34168 7814
rect 34216 7812 34272 7868
rect 34320 7866 34376 7868
rect 34424 7866 34480 7868
rect 34528 7866 34584 7868
rect 34320 7814 34324 7866
rect 34324 7814 34376 7866
rect 34424 7814 34448 7866
rect 34448 7814 34480 7866
rect 34528 7814 34572 7866
rect 34572 7814 34584 7866
rect 34320 7812 34376 7814
rect 34424 7812 34480 7814
rect 34528 7812 34584 7814
rect 34632 7866 34688 7868
rect 34736 7866 34792 7868
rect 34840 7866 34896 7868
rect 34632 7814 34644 7866
rect 34644 7814 34688 7866
rect 34736 7814 34768 7866
rect 34768 7814 34792 7866
rect 34840 7814 34892 7866
rect 34892 7814 34896 7866
rect 34632 7812 34688 7814
rect 34736 7812 34792 7814
rect 34840 7812 34896 7814
rect 34944 7812 35000 7868
rect 35048 7866 35104 7868
rect 35152 7866 35208 7868
rect 35048 7814 35068 7866
rect 35068 7814 35104 7866
rect 35152 7814 35192 7866
rect 35192 7814 35208 7866
rect 35048 7812 35104 7814
rect 35152 7812 35208 7814
rect 13804 7532 13860 7588
rect 14700 7644 14756 7700
rect 13580 7084 13636 7140
rect 14700 7474 14756 7476
rect 14700 7422 14702 7474
rect 14702 7422 14754 7474
rect 14754 7422 14756 7474
rect 14700 7420 14756 7422
rect 17612 7532 17668 7588
rect 13692 7308 13748 7364
rect 13468 6690 13524 6692
rect 13468 6638 13470 6690
rect 13470 6638 13522 6690
rect 13522 6638 13524 6690
rect 13468 6636 13524 6638
rect 13356 6524 13412 6580
rect 13020 3612 13076 3668
rect 12460 3442 12516 3444
rect 12460 3390 12462 3442
rect 12462 3390 12514 3442
rect 12514 3390 12516 3442
rect 12460 3388 12516 3390
rect 13580 5180 13636 5236
rect 13580 4956 13636 5012
rect 13580 4396 13636 4452
rect 13804 7084 13860 7140
rect 24008 7082 24064 7084
rect 24112 7082 24168 7084
rect 24008 7030 24024 7082
rect 24024 7030 24064 7082
rect 24112 7030 24148 7082
rect 24148 7030 24168 7082
rect 24008 7028 24064 7030
rect 24112 7028 24168 7030
rect 24216 7028 24272 7084
rect 24320 7082 24376 7084
rect 24424 7082 24480 7084
rect 24528 7082 24584 7084
rect 24320 7030 24324 7082
rect 24324 7030 24376 7082
rect 24424 7030 24448 7082
rect 24448 7030 24480 7082
rect 24528 7030 24572 7082
rect 24572 7030 24584 7082
rect 24320 7028 24376 7030
rect 24424 7028 24480 7030
rect 24528 7028 24584 7030
rect 24632 7082 24688 7084
rect 24736 7082 24792 7084
rect 24840 7082 24896 7084
rect 24632 7030 24644 7082
rect 24644 7030 24688 7082
rect 24736 7030 24768 7082
rect 24768 7030 24792 7082
rect 24840 7030 24892 7082
rect 24892 7030 24896 7082
rect 24632 7028 24688 7030
rect 24736 7028 24792 7030
rect 24840 7028 24896 7030
rect 24944 7028 25000 7084
rect 25048 7082 25104 7084
rect 25152 7082 25208 7084
rect 25048 7030 25068 7082
rect 25068 7030 25104 7082
rect 25152 7030 25192 7082
rect 25192 7030 25208 7082
rect 25048 7028 25104 7030
rect 25152 7028 25208 7030
rect 15148 6524 15204 6580
rect 14008 6298 14064 6300
rect 14112 6298 14168 6300
rect 14008 6246 14024 6298
rect 14024 6246 14064 6298
rect 14112 6246 14148 6298
rect 14148 6246 14168 6298
rect 14008 6244 14064 6246
rect 14112 6244 14168 6246
rect 14216 6244 14272 6300
rect 14320 6298 14376 6300
rect 14424 6298 14480 6300
rect 14528 6298 14584 6300
rect 14320 6246 14324 6298
rect 14324 6246 14376 6298
rect 14424 6246 14448 6298
rect 14448 6246 14480 6298
rect 14528 6246 14572 6298
rect 14572 6246 14584 6298
rect 14320 6244 14376 6246
rect 14424 6244 14480 6246
rect 14528 6244 14584 6246
rect 14632 6298 14688 6300
rect 14736 6298 14792 6300
rect 14840 6298 14896 6300
rect 14632 6246 14644 6298
rect 14644 6246 14688 6298
rect 14736 6246 14768 6298
rect 14768 6246 14792 6298
rect 14840 6246 14892 6298
rect 14892 6246 14896 6298
rect 14632 6244 14688 6246
rect 14736 6244 14792 6246
rect 14840 6244 14896 6246
rect 14944 6244 15000 6300
rect 15048 6298 15104 6300
rect 15152 6298 15208 6300
rect 15048 6246 15068 6298
rect 15068 6246 15104 6298
rect 15152 6246 15192 6298
rect 15192 6246 15208 6298
rect 15048 6244 15104 6246
rect 15152 6244 15208 6246
rect 13692 4060 13748 4116
rect 13804 5740 13860 5796
rect 14812 5906 14868 5908
rect 14812 5854 14814 5906
rect 14814 5854 14866 5906
rect 14866 5854 14868 5906
rect 14812 5852 14868 5854
rect 15372 5906 15428 5908
rect 15372 5854 15374 5906
rect 15374 5854 15426 5906
rect 15426 5854 15428 5906
rect 15372 5852 15428 5854
rect 13916 4956 13972 5012
rect 14008 4730 14064 4732
rect 14112 4730 14168 4732
rect 14008 4678 14024 4730
rect 14024 4678 14064 4730
rect 14112 4678 14148 4730
rect 14148 4678 14168 4730
rect 14008 4676 14064 4678
rect 14112 4676 14168 4678
rect 14216 4676 14272 4732
rect 14320 4730 14376 4732
rect 14424 4730 14480 4732
rect 14528 4730 14584 4732
rect 14320 4678 14324 4730
rect 14324 4678 14376 4730
rect 14424 4678 14448 4730
rect 14448 4678 14480 4730
rect 14528 4678 14572 4730
rect 14572 4678 14584 4730
rect 14320 4676 14376 4678
rect 14424 4676 14480 4678
rect 14528 4676 14584 4678
rect 14632 4730 14688 4732
rect 14736 4730 14792 4732
rect 14840 4730 14896 4732
rect 14632 4678 14644 4730
rect 14644 4678 14688 4730
rect 14736 4678 14768 4730
rect 14768 4678 14792 4730
rect 14840 4678 14892 4730
rect 14892 4678 14896 4730
rect 14632 4676 14688 4678
rect 14736 4676 14792 4678
rect 14840 4676 14896 4678
rect 14944 4676 15000 4732
rect 15048 4730 15104 4732
rect 15152 4730 15208 4732
rect 15048 4678 15068 4730
rect 15068 4678 15104 4730
rect 15152 4678 15192 4730
rect 15192 4678 15208 4730
rect 15048 4676 15104 4678
rect 15152 4676 15208 4678
rect 14812 4508 14868 4564
rect 14700 4060 14756 4116
rect 14028 3724 14084 3780
rect 15484 4508 15540 4564
rect 20524 6690 20580 6692
rect 20524 6638 20526 6690
rect 20526 6638 20578 6690
rect 20578 6638 20580 6690
rect 20524 6636 20580 6638
rect 21420 6690 21476 6692
rect 21420 6638 21422 6690
rect 21422 6638 21474 6690
rect 21474 6638 21476 6690
rect 21420 6636 21476 6638
rect 36428 6636 36484 6692
rect 15708 4732 15764 4788
rect 17388 6524 17444 6580
rect 16380 5852 16436 5908
rect 16156 5794 16212 5796
rect 16156 5742 16158 5794
rect 16158 5742 16210 5794
rect 16210 5742 16212 5794
rect 16156 5740 16212 5742
rect 16044 4844 16100 4900
rect 16268 5068 16324 5124
rect 15708 4508 15764 4564
rect 15260 3554 15316 3556
rect 15260 3502 15262 3554
rect 15262 3502 15314 3554
rect 15314 3502 15316 3554
rect 15260 3500 15316 3502
rect 14812 3442 14868 3444
rect 14812 3390 14814 3442
rect 14814 3390 14866 3442
rect 14866 3390 14868 3442
rect 14812 3388 14868 3390
rect 14008 3162 14064 3164
rect 14112 3162 14168 3164
rect 14008 3110 14024 3162
rect 14024 3110 14064 3162
rect 14112 3110 14148 3162
rect 14148 3110 14168 3162
rect 14008 3108 14064 3110
rect 14112 3108 14168 3110
rect 14216 3108 14272 3164
rect 14320 3162 14376 3164
rect 14424 3162 14480 3164
rect 14528 3162 14584 3164
rect 14320 3110 14324 3162
rect 14324 3110 14376 3162
rect 14424 3110 14448 3162
rect 14448 3110 14480 3162
rect 14528 3110 14572 3162
rect 14572 3110 14584 3162
rect 14320 3108 14376 3110
rect 14424 3108 14480 3110
rect 14528 3108 14584 3110
rect 14632 3162 14688 3164
rect 14736 3162 14792 3164
rect 14840 3162 14896 3164
rect 14632 3110 14644 3162
rect 14644 3110 14688 3162
rect 14736 3110 14768 3162
rect 14768 3110 14792 3162
rect 14840 3110 14892 3162
rect 14892 3110 14896 3162
rect 14632 3108 14688 3110
rect 14736 3108 14792 3110
rect 14840 3108 14896 3110
rect 14944 3108 15000 3164
rect 15048 3162 15104 3164
rect 15152 3162 15208 3164
rect 15048 3110 15068 3162
rect 15068 3110 15104 3162
rect 15152 3110 15192 3162
rect 15192 3110 15208 3162
rect 15048 3108 15104 3110
rect 15152 3108 15208 3110
rect 16380 4844 16436 4900
rect 16492 4956 16548 5012
rect 16380 4562 16436 4564
rect 16380 4510 16382 4562
rect 16382 4510 16434 4562
rect 16434 4510 16436 4562
rect 16380 4508 16436 4510
rect 16716 4844 16772 4900
rect 16716 4172 16772 4228
rect 17052 5010 17108 5012
rect 17052 4958 17054 5010
rect 17054 4958 17106 5010
rect 17106 4958 17108 5010
rect 17052 4956 17108 4958
rect 16940 3836 16996 3892
rect 19740 6578 19796 6580
rect 19740 6526 19742 6578
rect 19742 6526 19794 6578
rect 19794 6526 19796 6578
rect 19740 6524 19796 6526
rect 20748 6524 20804 6580
rect 34008 6298 34064 6300
rect 34112 6298 34168 6300
rect 34008 6246 34024 6298
rect 34024 6246 34064 6298
rect 34112 6246 34148 6298
rect 34148 6246 34168 6298
rect 34008 6244 34064 6246
rect 34112 6244 34168 6246
rect 34216 6244 34272 6300
rect 34320 6298 34376 6300
rect 34424 6298 34480 6300
rect 34528 6298 34584 6300
rect 34320 6246 34324 6298
rect 34324 6246 34376 6298
rect 34424 6246 34448 6298
rect 34448 6246 34480 6298
rect 34528 6246 34572 6298
rect 34572 6246 34584 6298
rect 34320 6244 34376 6246
rect 34424 6244 34480 6246
rect 34528 6244 34584 6246
rect 34632 6298 34688 6300
rect 34736 6298 34792 6300
rect 34840 6298 34896 6300
rect 34632 6246 34644 6298
rect 34644 6246 34688 6298
rect 34736 6246 34768 6298
rect 34768 6246 34792 6298
rect 34840 6246 34892 6298
rect 34892 6246 34896 6298
rect 34632 6244 34688 6246
rect 34736 6244 34792 6246
rect 34840 6244 34896 6246
rect 34944 6244 35000 6300
rect 35048 6298 35104 6300
rect 35152 6298 35208 6300
rect 35048 6246 35068 6298
rect 35068 6246 35104 6298
rect 35152 6246 35192 6298
rect 35192 6246 35208 6298
rect 35048 6244 35104 6246
rect 35152 6244 35208 6246
rect 17500 5068 17556 5124
rect 17724 3836 17780 3892
rect 18620 3724 18676 3780
rect 20076 4396 20132 4452
rect 20860 4450 20916 4452
rect 20860 4398 20862 4450
rect 20862 4398 20914 4450
rect 20914 4398 20916 4450
rect 20860 4396 20916 4398
rect 22764 4114 22820 4116
rect 22764 4062 22766 4114
rect 22766 4062 22818 4114
rect 22818 4062 22820 4114
rect 22764 4060 22820 4062
rect 23660 4956 23716 5012
rect 23436 4060 23492 4116
rect 24008 5514 24064 5516
rect 24112 5514 24168 5516
rect 24008 5462 24024 5514
rect 24024 5462 24064 5514
rect 24112 5462 24148 5514
rect 24148 5462 24168 5514
rect 24008 5460 24064 5462
rect 24112 5460 24168 5462
rect 24216 5460 24272 5516
rect 24320 5514 24376 5516
rect 24424 5514 24480 5516
rect 24528 5514 24584 5516
rect 24320 5462 24324 5514
rect 24324 5462 24376 5514
rect 24424 5462 24448 5514
rect 24448 5462 24480 5514
rect 24528 5462 24572 5514
rect 24572 5462 24584 5514
rect 24320 5460 24376 5462
rect 24424 5460 24480 5462
rect 24528 5460 24584 5462
rect 24632 5514 24688 5516
rect 24736 5514 24792 5516
rect 24840 5514 24896 5516
rect 24632 5462 24644 5514
rect 24644 5462 24688 5514
rect 24736 5462 24768 5514
rect 24768 5462 24792 5514
rect 24840 5462 24892 5514
rect 24892 5462 24896 5514
rect 24632 5460 24688 5462
rect 24736 5460 24792 5462
rect 24840 5460 24896 5462
rect 24944 5460 25000 5516
rect 25048 5514 25104 5516
rect 25152 5514 25208 5516
rect 25048 5462 25068 5514
rect 25068 5462 25104 5514
rect 25152 5462 25192 5514
rect 25192 5462 25208 5514
rect 25048 5460 25104 5462
rect 25152 5460 25208 5462
rect 24892 5010 24948 5012
rect 24892 4958 24894 5010
rect 24894 4958 24946 5010
rect 24946 4958 24948 5010
rect 24892 4956 24948 4958
rect 24108 4508 24164 4564
rect 25340 4562 25396 4564
rect 25340 4510 25342 4562
rect 25342 4510 25394 4562
rect 25394 4510 25396 4562
rect 25340 4508 25396 4510
rect 24556 4060 24612 4116
rect 24008 3946 24064 3948
rect 24112 3946 24168 3948
rect 24008 3894 24024 3946
rect 24024 3894 24064 3946
rect 24112 3894 24148 3946
rect 24148 3894 24168 3946
rect 24008 3892 24064 3894
rect 24112 3892 24168 3894
rect 24216 3892 24272 3948
rect 24320 3946 24376 3948
rect 24424 3946 24480 3948
rect 24528 3946 24584 3948
rect 24320 3894 24324 3946
rect 24324 3894 24376 3946
rect 24424 3894 24448 3946
rect 24448 3894 24480 3946
rect 24528 3894 24572 3946
rect 24572 3894 24584 3946
rect 24320 3892 24376 3894
rect 24424 3892 24480 3894
rect 24528 3892 24584 3894
rect 24632 3946 24688 3948
rect 24736 3946 24792 3948
rect 24840 3946 24896 3948
rect 24632 3894 24644 3946
rect 24644 3894 24688 3946
rect 24736 3894 24768 3946
rect 24768 3894 24792 3946
rect 24840 3894 24892 3946
rect 24892 3894 24896 3946
rect 24632 3892 24688 3894
rect 24736 3892 24792 3894
rect 24840 3892 24896 3894
rect 24944 3892 25000 3948
rect 25048 3946 25104 3948
rect 25152 3946 25208 3948
rect 25048 3894 25068 3946
rect 25068 3894 25104 3946
rect 25152 3894 25192 3946
rect 25192 3894 25208 3946
rect 25048 3892 25104 3894
rect 25152 3892 25208 3894
rect 25116 3612 25172 3668
rect 24556 3442 24612 3444
rect 24556 3390 24558 3442
rect 24558 3390 24610 3442
rect 24610 3390 24612 3442
rect 24556 3388 24612 3390
rect 25788 3388 25844 3444
rect 26684 3388 26740 3444
rect 27692 3666 27748 3668
rect 27692 3614 27694 3666
rect 27694 3614 27746 3666
rect 27746 3614 27748 3666
rect 27692 3612 27748 3614
rect 27132 3388 27188 3444
rect 27580 3500 27636 3556
rect 28588 3554 28644 3556
rect 28588 3502 28590 3554
rect 28590 3502 28642 3554
rect 28642 3502 28644 3554
rect 28588 3500 28644 3502
rect 28476 3388 28532 3444
rect 29036 3442 29092 3444
rect 29036 3390 29038 3442
rect 29038 3390 29090 3442
rect 29090 3390 29092 3442
rect 29036 3388 29092 3390
rect 29484 3388 29540 3444
rect 30828 4956 30884 5012
rect 32844 5010 32900 5012
rect 32844 4958 32846 5010
rect 32846 4958 32898 5010
rect 32898 4958 32900 5010
rect 32844 4956 32900 4958
rect 32060 4284 32116 4340
rect 33180 4284 33236 4340
rect 33628 3612 33684 3668
rect 34412 4898 34468 4900
rect 34412 4846 34414 4898
rect 34414 4846 34466 4898
rect 34466 4846 34468 4898
rect 34412 4844 34468 4846
rect 34008 4730 34064 4732
rect 34112 4730 34168 4732
rect 34008 4678 34024 4730
rect 34024 4678 34064 4730
rect 34112 4678 34148 4730
rect 34148 4678 34168 4730
rect 34008 4676 34064 4678
rect 34112 4676 34168 4678
rect 34216 4676 34272 4732
rect 34320 4730 34376 4732
rect 34424 4730 34480 4732
rect 34528 4730 34584 4732
rect 34320 4678 34324 4730
rect 34324 4678 34376 4730
rect 34424 4678 34448 4730
rect 34448 4678 34480 4730
rect 34528 4678 34572 4730
rect 34572 4678 34584 4730
rect 34320 4676 34376 4678
rect 34424 4676 34480 4678
rect 34528 4676 34584 4678
rect 34632 4730 34688 4732
rect 34736 4730 34792 4732
rect 34840 4730 34896 4732
rect 34632 4678 34644 4730
rect 34644 4678 34688 4730
rect 34736 4678 34768 4730
rect 34768 4678 34792 4730
rect 34840 4678 34892 4730
rect 34892 4678 34896 4730
rect 34632 4676 34688 4678
rect 34736 4676 34792 4678
rect 34840 4676 34896 4678
rect 34944 4676 35000 4732
rect 35048 4730 35104 4732
rect 35152 4730 35208 4732
rect 35048 4678 35068 4730
rect 35068 4678 35104 4730
rect 35152 4678 35192 4730
rect 35192 4678 35208 4730
rect 35048 4676 35104 4678
rect 35152 4676 35208 4678
rect 33964 4338 34020 4340
rect 33964 4286 33966 4338
rect 33966 4286 34018 4338
rect 34018 4286 34020 4338
rect 33964 4284 34020 4286
rect 34412 4338 34468 4340
rect 34412 4286 34414 4338
rect 34414 4286 34466 4338
rect 34466 4286 34468 4338
rect 34412 4284 34468 4286
rect 35756 4284 35812 4340
rect 35308 3612 35364 3668
rect 35644 4172 35700 4228
rect 33852 3388 33908 3444
rect 34524 3442 34580 3444
rect 34524 3390 34526 3442
rect 34526 3390 34578 3442
rect 34578 3390 34580 3442
rect 34524 3388 34580 3390
rect 35308 3388 35364 3444
rect 34008 3162 34064 3164
rect 34112 3162 34168 3164
rect 34008 3110 34024 3162
rect 34024 3110 34064 3162
rect 34112 3110 34148 3162
rect 34148 3110 34168 3162
rect 34008 3108 34064 3110
rect 34112 3108 34168 3110
rect 34216 3108 34272 3164
rect 34320 3162 34376 3164
rect 34424 3162 34480 3164
rect 34528 3162 34584 3164
rect 34320 3110 34324 3162
rect 34324 3110 34376 3162
rect 34424 3110 34448 3162
rect 34448 3110 34480 3162
rect 34528 3110 34572 3162
rect 34572 3110 34584 3162
rect 34320 3108 34376 3110
rect 34424 3108 34480 3110
rect 34528 3108 34584 3110
rect 34632 3162 34688 3164
rect 34736 3162 34792 3164
rect 34840 3162 34896 3164
rect 34632 3110 34644 3162
rect 34644 3110 34688 3162
rect 34736 3110 34768 3162
rect 34768 3110 34792 3162
rect 34840 3110 34892 3162
rect 34892 3110 34896 3162
rect 34632 3108 34688 3110
rect 34736 3108 34792 3110
rect 34840 3108 34896 3110
rect 34944 3108 35000 3164
rect 35048 3162 35104 3164
rect 35152 3162 35208 3164
rect 35048 3110 35068 3162
rect 35068 3110 35104 3162
rect 35152 3110 35192 3162
rect 35192 3110 35208 3162
rect 35048 3108 35104 3110
rect 35152 3108 35208 3110
rect 36204 3388 36260 3444
rect 37660 6300 37716 6356
rect 38220 6300 38276 6356
rect 37212 4060 37268 4116
<< metal3 >>
rect 0 47124 800 47152
rect 0 47068 2100 47124
rect 0 47040 800 47068
rect 2044 47012 2100 47068
rect 2034 46956 2044 47012
rect 2100 46956 2110 47012
rect 3998 46228 4008 46284
rect 4064 46228 4112 46284
rect 4168 46228 4216 46284
rect 4272 46228 4320 46284
rect 4376 46228 4424 46284
rect 4480 46228 4528 46284
rect 4584 46228 4632 46284
rect 4688 46228 4736 46284
rect 4792 46228 4840 46284
rect 4896 46228 4944 46284
rect 5000 46228 5048 46284
rect 5104 46228 5152 46284
rect 5208 46228 5218 46284
rect 23998 46228 24008 46284
rect 24064 46228 24112 46284
rect 24168 46228 24216 46284
rect 24272 46228 24320 46284
rect 24376 46228 24424 46284
rect 24480 46228 24528 46284
rect 24584 46228 24632 46284
rect 24688 46228 24736 46284
rect 24792 46228 24840 46284
rect 24896 46228 24944 46284
rect 25000 46228 25048 46284
rect 25104 46228 25152 46284
rect 25208 46228 25218 46284
rect 27346 46060 27356 46116
rect 27412 46060 28812 46116
rect 28868 46060 28878 46116
rect 12562 45948 12572 46004
rect 12628 45948 13580 46004
rect 13636 45948 13646 46004
rect 0 45780 800 45808
rect 0 45724 2156 45780
rect 2212 45724 2222 45780
rect 0 45696 800 45724
rect 13998 45444 14008 45500
rect 14064 45444 14112 45500
rect 14168 45444 14216 45500
rect 14272 45444 14320 45500
rect 14376 45444 14424 45500
rect 14480 45444 14528 45500
rect 14584 45444 14632 45500
rect 14688 45444 14736 45500
rect 14792 45444 14840 45500
rect 14896 45444 14944 45500
rect 15000 45444 15048 45500
rect 15104 45444 15152 45500
rect 15208 45444 15218 45500
rect 33998 45444 34008 45500
rect 34064 45444 34112 45500
rect 34168 45444 34216 45500
rect 34272 45444 34320 45500
rect 34376 45444 34424 45500
rect 34480 45444 34528 45500
rect 34584 45444 34632 45500
rect 34688 45444 34736 45500
rect 34792 45444 34840 45500
rect 34896 45444 34944 45500
rect 35000 45444 35048 45500
rect 35104 45444 35152 45500
rect 35208 45444 35218 45500
rect 1810 44940 1820 44996
rect 1876 44940 2716 44996
rect 2772 44940 3500 44996
rect 3556 44940 3566 44996
rect 3998 44660 4008 44716
rect 4064 44660 4112 44716
rect 4168 44660 4216 44716
rect 4272 44660 4320 44716
rect 4376 44660 4424 44716
rect 4480 44660 4528 44716
rect 4584 44660 4632 44716
rect 4688 44660 4736 44716
rect 4792 44660 4840 44716
rect 4896 44660 4944 44716
rect 5000 44660 5048 44716
rect 5104 44660 5152 44716
rect 5208 44660 5218 44716
rect 23998 44660 24008 44716
rect 24064 44660 24112 44716
rect 24168 44660 24216 44716
rect 24272 44660 24320 44716
rect 24376 44660 24424 44716
rect 24480 44660 24528 44716
rect 24584 44660 24632 44716
rect 24688 44660 24736 44716
rect 24792 44660 24840 44716
rect 24896 44660 24944 44716
rect 25000 44660 25048 44716
rect 25104 44660 25152 44716
rect 25208 44660 25218 44716
rect 0 44436 800 44464
rect 0 44380 1708 44436
rect 1764 44380 1774 44436
rect 0 44352 800 44380
rect 13998 43876 14008 43932
rect 14064 43876 14112 43932
rect 14168 43876 14216 43932
rect 14272 43876 14320 43932
rect 14376 43876 14424 43932
rect 14480 43876 14528 43932
rect 14584 43876 14632 43932
rect 14688 43876 14736 43932
rect 14792 43876 14840 43932
rect 14896 43876 14944 43932
rect 15000 43876 15048 43932
rect 15104 43876 15152 43932
rect 15208 43876 15218 43932
rect 33998 43876 34008 43932
rect 34064 43876 34112 43932
rect 34168 43876 34216 43932
rect 34272 43876 34320 43932
rect 34376 43876 34424 43932
rect 34480 43876 34528 43932
rect 34584 43876 34632 43932
rect 34688 43876 34736 43932
rect 34792 43876 34840 43932
rect 34896 43876 34944 43932
rect 35000 43876 35048 43932
rect 35104 43876 35152 43932
rect 35208 43876 35218 43932
rect 39200 43316 40000 43344
rect 38210 43260 38220 43316
rect 38276 43260 40000 43316
rect 39200 43232 40000 43260
rect 0 43092 800 43120
rect 3998 43092 4008 43148
rect 4064 43092 4112 43148
rect 4168 43092 4216 43148
rect 4272 43092 4320 43148
rect 4376 43092 4424 43148
rect 4480 43092 4528 43148
rect 4584 43092 4632 43148
rect 4688 43092 4736 43148
rect 4792 43092 4840 43148
rect 4896 43092 4944 43148
rect 5000 43092 5048 43148
rect 5104 43092 5152 43148
rect 5208 43092 5218 43148
rect 23998 43092 24008 43148
rect 24064 43092 24112 43148
rect 24168 43092 24216 43148
rect 24272 43092 24320 43148
rect 24376 43092 24424 43148
rect 24480 43092 24528 43148
rect 24584 43092 24632 43148
rect 24688 43092 24736 43148
rect 24792 43092 24840 43148
rect 24896 43092 24944 43148
rect 25000 43092 25048 43148
rect 25104 43092 25152 43148
rect 25208 43092 25218 43148
rect 0 43036 1708 43092
rect 1764 43036 1774 43092
rect 0 43008 800 43036
rect 13998 42308 14008 42364
rect 14064 42308 14112 42364
rect 14168 42308 14216 42364
rect 14272 42308 14320 42364
rect 14376 42308 14424 42364
rect 14480 42308 14528 42364
rect 14584 42308 14632 42364
rect 14688 42308 14736 42364
rect 14792 42308 14840 42364
rect 14896 42308 14944 42364
rect 15000 42308 15048 42364
rect 15104 42308 15152 42364
rect 15208 42308 15218 42364
rect 33998 42308 34008 42364
rect 34064 42308 34112 42364
rect 34168 42308 34216 42364
rect 34272 42308 34320 42364
rect 34376 42308 34424 42364
rect 34480 42308 34528 42364
rect 34584 42308 34632 42364
rect 34688 42308 34736 42364
rect 34792 42308 34840 42364
rect 34896 42308 34944 42364
rect 35000 42308 35048 42364
rect 35104 42308 35152 42364
rect 35208 42308 35218 42364
rect 0 41748 800 41776
rect 0 41692 1708 41748
rect 1764 41692 1774 41748
rect 0 41664 800 41692
rect 3998 41524 4008 41580
rect 4064 41524 4112 41580
rect 4168 41524 4216 41580
rect 4272 41524 4320 41580
rect 4376 41524 4424 41580
rect 4480 41524 4528 41580
rect 4584 41524 4632 41580
rect 4688 41524 4736 41580
rect 4792 41524 4840 41580
rect 4896 41524 4944 41580
rect 5000 41524 5048 41580
rect 5104 41524 5152 41580
rect 5208 41524 5218 41580
rect 23998 41524 24008 41580
rect 24064 41524 24112 41580
rect 24168 41524 24216 41580
rect 24272 41524 24320 41580
rect 24376 41524 24424 41580
rect 24480 41524 24528 41580
rect 24584 41524 24632 41580
rect 24688 41524 24736 41580
rect 24792 41524 24840 41580
rect 24896 41524 24944 41580
rect 25000 41524 25048 41580
rect 25104 41524 25152 41580
rect 25208 41524 25218 41580
rect 13998 40740 14008 40796
rect 14064 40740 14112 40796
rect 14168 40740 14216 40796
rect 14272 40740 14320 40796
rect 14376 40740 14424 40796
rect 14480 40740 14528 40796
rect 14584 40740 14632 40796
rect 14688 40740 14736 40796
rect 14792 40740 14840 40796
rect 14896 40740 14944 40796
rect 15000 40740 15048 40796
rect 15104 40740 15152 40796
rect 15208 40740 15218 40796
rect 33998 40740 34008 40796
rect 34064 40740 34112 40796
rect 34168 40740 34216 40796
rect 34272 40740 34320 40796
rect 34376 40740 34424 40796
rect 34480 40740 34528 40796
rect 34584 40740 34632 40796
rect 34688 40740 34736 40796
rect 34792 40740 34840 40796
rect 34896 40740 34944 40796
rect 35000 40740 35048 40796
rect 35104 40740 35152 40796
rect 35208 40740 35218 40796
rect 0 40404 800 40432
rect 0 40348 1708 40404
rect 1764 40348 1774 40404
rect 0 40320 800 40348
rect 3998 39956 4008 40012
rect 4064 39956 4112 40012
rect 4168 39956 4216 40012
rect 4272 39956 4320 40012
rect 4376 39956 4424 40012
rect 4480 39956 4528 40012
rect 4584 39956 4632 40012
rect 4688 39956 4736 40012
rect 4792 39956 4840 40012
rect 4896 39956 4944 40012
rect 5000 39956 5048 40012
rect 5104 39956 5152 40012
rect 5208 39956 5218 40012
rect 23998 39956 24008 40012
rect 24064 39956 24112 40012
rect 24168 39956 24216 40012
rect 24272 39956 24320 40012
rect 24376 39956 24424 40012
rect 24480 39956 24528 40012
rect 24584 39956 24632 40012
rect 24688 39956 24736 40012
rect 24792 39956 24840 40012
rect 24896 39956 24944 40012
rect 25000 39956 25048 40012
rect 25104 39956 25152 40012
rect 25208 39956 25218 40012
rect 13998 39172 14008 39228
rect 14064 39172 14112 39228
rect 14168 39172 14216 39228
rect 14272 39172 14320 39228
rect 14376 39172 14424 39228
rect 14480 39172 14528 39228
rect 14584 39172 14632 39228
rect 14688 39172 14736 39228
rect 14792 39172 14840 39228
rect 14896 39172 14944 39228
rect 15000 39172 15048 39228
rect 15104 39172 15152 39228
rect 15208 39172 15218 39228
rect 33998 39172 34008 39228
rect 34064 39172 34112 39228
rect 34168 39172 34216 39228
rect 34272 39172 34320 39228
rect 34376 39172 34424 39228
rect 34480 39172 34528 39228
rect 34584 39172 34632 39228
rect 34688 39172 34736 39228
rect 34792 39172 34840 39228
rect 34896 39172 34944 39228
rect 35000 39172 35048 39228
rect 35104 39172 35152 39228
rect 35208 39172 35218 39228
rect 0 39060 800 39088
rect 0 39004 1708 39060
rect 1764 39004 1774 39060
rect 0 38976 800 39004
rect 3998 38388 4008 38444
rect 4064 38388 4112 38444
rect 4168 38388 4216 38444
rect 4272 38388 4320 38444
rect 4376 38388 4424 38444
rect 4480 38388 4528 38444
rect 4584 38388 4632 38444
rect 4688 38388 4736 38444
rect 4792 38388 4840 38444
rect 4896 38388 4944 38444
rect 5000 38388 5048 38444
rect 5104 38388 5152 38444
rect 5208 38388 5218 38444
rect 23998 38388 24008 38444
rect 24064 38388 24112 38444
rect 24168 38388 24216 38444
rect 24272 38388 24320 38444
rect 24376 38388 24424 38444
rect 24480 38388 24528 38444
rect 24584 38388 24632 38444
rect 24688 38388 24736 38444
rect 24792 38388 24840 38444
rect 24896 38388 24944 38444
rect 25000 38388 25048 38444
rect 25104 38388 25152 38444
rect 25208 38388 25218 38444
rect 1698 37772 1708 37828
rect 1764 37772 1774 37828
rect 0 37716 800 37744
rect 1708 37716 1764 37772
rect 0 37660 1764 37716
rect 0 37632 800 37660
rect 13998 37604 14008 37660
rect 14064 37604 14112 37660
rect 14168 37604 14216 37660
rect 14272 37604 14320 37660
rect 14376 37604 14424 37660
rect 14480 37604 14528 37660
rect 14584 37604 14632 37660
rect 14688 37604 14736 37660
rect 14792 37604 14840 37660
rect 14896 37604 14944 37660
rect 15000 37604 15048 37660
rect 15104 37604 15152 37660
rect 15208 37604 15218 37660
rect 33998 37604 34008 37660
rect 34064 37604 34112 37660
rect 34168 37604 34216 37660
rect 34272 37604 34320 37660
rect 34376 37604 34424 37660
rect 34480 37604 34528 37660
rect 34584 37604 34632 37660
rect 34688 37604 34736 37660
rect 34792 37604 34840 37660
rect 34896 37604 34944 37660
rect 35000 37604 35048 37660
rect 35104 37604 35152 37660
rect 35208 37604 35218 37660
rect 3998 36820 4008 36876
rect 4064 36820 4112 36876
rect 4168 36820 4216 36876
rect 4272 36820 4320 36876
rect 4376 36820 4424 36876
rect 4480 36820 4528 36876
rect 4584 36820 4632 36876
rect 4688 36820 4736 36876
rect 4792 36820 4840 36876
rect 4896 36820 4944 36876
rect 5000 36820 5048 36876
rect 5104 36820 5152 36876
rect 5208 36820 5218 36876
rect 23998 36820 24008 36876
rect 24064 36820 24112 36876
rect 24168 36820 24216 36876
rect 24272 36820 24320 36876
rect 24376 36820 24424 36876
rect 24480 36820 24528 36876
rect 24584 36820 24632 36876
rect 24688 36820 24736 36876
rect 24792 36820 24840 36876
rect 24896 36820 24944 36876
rect 25000 36820 25048 36876
rect 25104 36820 25152 36876
rect 25208 36820 25218 36876
rect 0 36372 800 36400
rect 0 36316 1708 36372
rect 1764 36316 1774 36372
rect 0 36288 800 36316
rect 13998 36036 14008 36092
rect 14064 36036 14112 36092
rect 14168 36036 14216 36092
rect 14272 36036 14320 36092
rect 14376 36036 14424 36092
rect 14480 36036 14528 36092
rect 14584 36036 14632 36092
rect 14688 36036 14736 36092
rect 14792 36036 14840 36092
rect 14896 36036 14944 36092
rect 15000 36036 15048 36092
rect 15104 36036 15152 36092
rect 15208 36036 15218 36092
rect 33998 36036 34008 36092
rect 34064 36036 34112 36092
rect 34168 36036 34216 36092
rect 34272 36036 34320 36092
rect 34376 36036 34424 36092
rect 34480 36036 34528 36092
rect 34584 36036 34632 36092
rect 34688 36036 34736 36092
rect 34792 36036 34840 36092
rect 34896 36036 34944 36092
rect 35000 36036 35048 36092
rect 35104 36036 35152 36092
rect 35208 36036 35218 36092
rect 3998 35252 4008 35308
rect 4064 35252 4112 35308
rect 4168 35252 4216 35308
rect 4272 35252 4320 35308
rect 4376 35252 4424 35308
rect 4480 35252 4528 35308
rect 4584 35252 4632 35308
rect 4688 35252 4736 35308
rect 4792 35252 4840 35308
rect 4896 35252 4944 35308
rect 5000 35252 5048 35308
rect 5104 35252 5152 35308
rect 5208 35252 5218 35308
rect 23998 35252 24008 35308
rect 24064 35252 24112 35308
rect 24168 35252 24216 35308
rect 24272 35252 24320 35308
rect 24376 35252 24424 35308
rect 24480 35252 24528 35308
rect 24584 35252 24632 35308
rect 24688 35252 24736 35308
rect 24792 35252 24840 35308
rect 24896 35252 24944 35308
rect 25000 35252 25048 35308
rect 25104 35252 25152 35308
rect 25208 35252 25218 35308
rect 0 35028 800 35056
rect 0 34972 1708 35028
rect 1764 34972 1774 35028
rect 0 34944 800 34972
rect 13998 34468 14008 34524
rect 14064 34468 14112 34524
rect 14168 34468 14216 34524
rect 14272 34468 14320 34524
rect 14376 34468 14424 34524
rect 14480 34468 14528 34524
rect 14584 34468 14632 34524
rect 14688 34468 14736 34524
rect 14792 34468 14840 34524
rect 14896 34468 14944 34524
rect 15000 34468 15048 34524
rect 15104 34468 15152 34524
rect 15208 34468 15218 34524
rect 33998 34468 34008 34524
rect 34064 34468 34112 34524
rect 34168 34468 34216 34524
rect 34272 34468 34320 34524
rect 34376 34468 34424 34524
rect 34480 34468 34528 34524
rect 34584 34468 34632 34524
rect 34688 34468 34736 34524
rect 34792 34468 34840 34524
rect 34896 34468 34944 34524
rect 35000 34468 35048 34524
rect 35104 34468 35152 34524
rect 35208 34468 35218 34524
rect 0 33684 800 33712
rect 3998 33684 4008 33740
rect 4064 33684 4112 33740
rect 4168 33684 4216 33740
rect 4272 33684 4320 33740
rect 4376 33684 4424 33740
rect 4480 33684 4528 33740
rect 4584 33684 4632 33740
rect 4688 33684 4736 33740
rect 4792 33684 4840 33740
rect 4896 33684 4944 33740
rect 5000 33684 5048 33740
rect 5104 33684 5152 33740
rect 5208 33684 5218 33740
rect 23998 33684 24008 33740
rect 24064 33684 24112 33740
rect 24168 33684 24216 33740
rect 24272 33684 24320 33740
rect 24376 33684 24424 33740
rect 24480 33684 24528 33740
rect 24584 33684 24632 33740
rect 24688 33684 24736 33740
rect 24792 33684 24840 33740
rect 24896 33684 24944 33740
rect 25000 33684 25048 33740
rect 25104 33684 25152 33740
rect 25208 33684 25218 33740
rect 0 33628 1708 33684
rect 1764 33628 1774 33684
rect 0 33600 800 33628
rect 13998 32900 14008 32956
rect 14064 32900 14112 32956
rect 14168 32900 14216 32956
rect 14272 32900 14320 32956
rect 14376 32900 14424 32956
rect 14480 32900 14528 32956
rect 14584 32900 14632 32956
rect 14688 32900 14736 32956
rect 14792 32900 14840 32956
rect 14896 32900 14944 32956
rect 15000 32900 15048 32956
rect 15104 32900 15152 32956
rect 15208 32900 15218 32956
rect 33998 32900 34008 32956
rect 34064 32900 34112 32956
rect 34168 32900 34216 32956
rect 34272 32900 34320 32956
rect 34376 32900 34424 32956
rect 34480 32900 34528 32956
rect 34584 32900 34632 32956
rect 34688 32900 34736 32956
rect 34792 32900 34840 32956
rect 34896 32900 34944 32956
rect 35000 32900 35048 32956
rect 35104 32900 35152 32956
rect 35208 32900 35218 32956
rect 0 32340 800 32368
rect 0 32284 1708 32340
rect 1764 32284 1774 32340
rect 0 32256 800 32284
rect 3998 32116 4008 32172
rect 4064 32116 4112 32172
rect 4168 32116 4216 32172
rect 4272 32116 4320 32172
rect 4376 32116 4424 32172
rect 4480 32116 4528 32172
rect 4584 32116 4632 32172
rect 4688 32116 4736 32172
rect 4792 32116 4840 32172
rect 4896 32116 4944 32172
rect 5000 32116 5048 32172
rect 5104 32116 5152 32172
rect 5208 32116 5218 32172
rect 23998 32116 24008 32172
rect 24064 32116 24112 32172
rect 24168 32116 24216 32172
rect 24272 32116 24320 32172
rect 24376 32116 24424 32172
rect 24480 32116 24528 32172
rect 24584 32116 24632 32172
rect 24688 32116 24736 32172
rect 24792 32116 24840 32172
rect 24896 32116 24944 32172
rect 25000 32116 25048 32172
rect 25104 32116 25152 32172
rect 25208 32116 25218 32172
rect 37650 31500 37660 31556
rect 37716 31500 38220 31556
rect 38276 31500 38286 31556
rect 13998 31332 14008 31388
rect 14064 31332 14112 31388
rect 14168 31332 14216 31388
rect 14272 31332 14320 31388
rect 14376 31332 14424 31388
rect 14480 31332 14528 31388
rect 14584 31332 14632 31388
rect 14688 31332 14736 31388
rect 14792 31332 14840 31388
rect 14896 31332 14944 31388
rect 15000 31332 15048 31388
rect 15104 31332 15152 31388
rect 15208 31332 15218 31388
rect 33998 31332 34008 31388
rect 34064 31332 34112 31388
rect 34168 31332 34216 31388
rect 34272 31332 34320 31388
rect 34376 31332 34424 31388
rect 34480 31332 34528 31388
rect 34584 31332 34632 31388
rect 34688 31332 34736 31388
rect 34792 31332 34840 31388
rect 34896 31332 34944 31388
rect 35000 31332 35048 31388
rect 35104 31332 35152 31388
rect 35208 31332 35218 31388
rect 0 30996 800 31024
rect 39200 30996 40000 31024
rect 0 30940 1708 30996
rect 1764 30940 1774 30996
rect 38210 30940 38220 30996
rect 38276 30940 40000 30996
rect 0 30912 800 30940
rect 39200 30912 40000 30940
rect 3998 30548 4008 30604
rect 4064 30548 4112 30604
rect 4168 30548 4216 30604
rect 4272 30548 4320 30604
rect 4376 30548 4424 30604
rect 4480 30548 4528 30604
rect 4584 30548 4632 30604
rect 4688 30548 4736 30604
rect 4792 30548 4840 30604
rect 4896 30548 4944 30604
rect 5000 30548 5048 30604
rect 5104 30548 5152 30604
rect 5208 30548 5218 30604
rect 23998 30548 24008 30604
rect 24064 30548 24112 30604
rect 24168 30548 24216 30604
rect 24272 30548 24320 30604
rect 24376 30548 24424 30604
rect 24480 30548 24528 30604
rect 24584 30548 24632 30604
rect 24688 30548 24736 30604
rect 24792 30548 24840 30604
rect 24896 30548 24944 30604
rect 25000 30548 25048 30604
rect 25104 30548 25152 30604
rect 25208 30548 25218 30604
rect 13998 29764 14008 29820
rect 14064 29764 14112 29820
rect 14168 29764 14216 29820
rect 14272 29764 14320 29820
rect 14376 29764 14424 29820
rect 14480 29764 14528 29820
rect 14584 29764 14632 29820
rect 14688 29764 14736 29820
rect 14792 29764 14840 29820
rect 14896 29764 14944 29820
rect 15000 29764 15048 29820
rect 15104 29764 15152 29820
rect 15208 29764 15218 29820
rect 33998 29764 34008 29820
rect 34064 29764 34112 29820
rect 34168 29764 34216 29820
rect 34272 29764 34320 29820
rect 34376 29764 34424 29820
rect 34480 29764 34528 29820
rect 34584 29764 34632 29820
rect 34688 29764 34736 29820
rect 34792 29764 34840 29820
rect 34896 29764 34944 29820
rect 35000 29764 35048 29820
rect 35104 29764 35152 29820
rect 35208 29764 35218 29820
rect 0 29652 800 29680
rect 0 29596 1708 29652
rect 1764 29596 1774 29652
rect 0 29568 800 29596
rect 3998 28980 4008 29036
rect 4064 28980 4112 29036
rect 4168 28980 4216 29036
rect 4272 28980 4320 29036
rect 4376 28980 4424 29036
rect 4480 28980 4528 29036
rect 4584 28980 4632 29036
rect 4688 28980 4736 29036
rect 4792 28980 4840 29036
rect 4896 28980 4944 29036
rect 5000 28980 5048 29036
rect 5104 28980 5152 29036
rect 5208 28980 5218 29036
rect 23998 28980 24008 29036
rect 24064 28980 24112 29036
rect 24168 28980 24216 29036
rect 24272 28980 24320 29036
rect 24376 28980 24424 29036
rect 24480 28980 24528 29036
rect 24584 28980 24632 29036
rect 24688 28980 24736 29036
rect 24792 28980 24840 29036
rect 24896 28980 24944 29036
rect 25000 28980 25048 29036
rect 25104 28980 25152 29036
rect 25208 28980 25218 29036
rect 1698 28364 1708 28420
rect 1764 28364 1774 28420
rect 0 28308 800 28336
rect 1708 28308 1764 28364
rect 0 28252 1764 28308
rect 0 28224 800 28252
rect 13998 28196 14008 28252
rect 14064 28196 14112 28252
rect 14168 28196 14216 28252
rect 14272 28196 14320 28252
rect 14376 28196 14424 28252
rect 14480 28196 14528 28252
rect 14584 28196 14632 28252
rect 14688 28196 14736 28252
rect 14792 28196 14840 28252
rect 14896 28196 14944 28252
rect 15000 28196 15048 28252
rect 15104 28196 15152 28252
rect 15208 28196 15218 28252
rect 33998 28196 34008 28252
rect 34064 28196 34112 28252
rect 34168 28196 34216 28252
rect 34272 28196 34320 28252
rect 34376 28196 34424 28252
rect 34480 28196 34528 28252
rect 34584 28196 34632 28252
rect 34688 28196 34736 28252
rect 34792 28196 34840 28252
rect 34896 28196 34944 28252
rect 35000 28196 35048 28252
rect 35104 28196 35152 28252
rect 35208 28196 35218 28252
rect 3998 27412 4008 27468
rect 4064 27412 4112 27468
rect 4168 27412 4216 27468
rect 4272 27412 4320 27468
rect 4376 27412 4424 27468
rect 4480 27412 4528 27468
rect 4584 27412 4632 27468
rect 4688 27412 4736 27468
rect 4792 27412 4840 27468
rect 4896 27412 4944 27468
rect 5000 27412 5048 27468
rect 5104 27412 5152 27468
rect 5208 27412 5218 27468
rect 23998 27412 24008 27468
rect 24064 27412 24112 27468
rect 24168 27412 24216 27468
rect 24272 27412 24320 27468
rect 24376 27412 24424 27468
rect 24480 27412 24528 27468
rect 24584 27412 24632 27468
rect 24688 27412 24736 27468
rect 24792 27412 24840 27468
rect 24896 27412 24944 27468
rect 25000 27412 25048 27468
rect 25104 27412 25152 27468
rect 25208 27412 25218 27468
rect 0 26964 800 26992
rect 0 26908 1708 26964
rect 1764 26908 1774 26964
rect 0 26880 800 26908
rect 13998 26628 14008 26684
rect 14064 26628 14112 26684
rect 14168 26628 14216 26684
rect 14272 26628 14320 26684
rect 14376 26628 14424 26684
rect 14480 26628 14528 26684
rect 14584 26628 14632 26684
rect 14688 26628 14736 26684
rect 14792 26628 14840 26684
rect 14896 26628 14944 26684
rect 15000 26628 15048 26684
rect 15104 26628 15152 26684
rect 15208 26628 15218 26684
rect 33998 26628 34008 26684
rect 34064 26628 34112 26684
rect 34168 26628 34216 26684
rect 34272 26628 34320 26684
rect 34376 26628 34424 26684
rect 34480 26628 34528 26684
rect 34584 26628 34632 26684
rect 34688 26628 34736 26684
rect 34792 26628 34840 26684
rect 34896 26628 34944 26684
rect 35000 26628 35048 26684
rect 35104 26628 35152 26684
rect 35208 26628 35218 26684
rect 3998 25844 4008 25900
rect 4064 25844 4112 25900
rect 4168 25844 4216 25900
rect 4272 25844 4320 25900
rect 4376 25844 4424 25900
rect 4480 25844 4528 25900
rect 4584 25844 4632 25900
rect 4688 25844 4736 25900
rect 4792 25844 4840 25900
rect 4896 25844 4944 25900
rect 5000 25844 5048 25900
rect 5104 25844 5152 25900
rect 5208 25844 5218 25900
rect 23998 25844 24008 25900
rect 24064 25844 24112 25900
rect 24168 25844 24216 25900
rect 24272 25844 24320 25900
rect 24376 25844 24424 25900
rect 24480 25844 24528 25900
rect 24584 25844 24632 25900
rect 24688 25844 24736 25900
rect 24792 25844 24840 25900
rect 24896 25844 24944 25900
rect 25000 25844 25048 25900
rect 25104 25844 25152 25900
rect 25208 25844 25218 25900
rect 0 25620 800 25648
rect 0 25564 1708 25620
rect 1764 25564 1774 25620
rect 0 25536 800 25564
rect 13998 25060 14008 25116
rect 14064 25060 14112 25116
rect 14168 25060 14216 25116
rect 14272 25060 14320 25116
rect 14376 25060 14424 25116
rect 14480 25060 14528 25116
rect 14584 25060 14632 25116
rect 14688 25060 14736 25116
rect 14792 25060 14840 25116
rect 14896 25060 14944 25116
rect 15000 25060 15048 25116
rect 15104 25060 15152 25116
rect 15208 25060 15218 25116
rect 33998 25060 34008 25116
rect 34064 25060 34112 25116
rect 34168 25060 34216 25116
rect 34272 25060 34320 25116
rect 34376 25060 34424 25116
rect 34480 25060 34528 25116
rect 34584 25060 34632 25116
rect 34688 25060 34736 25116
rect 34792 25060 34840 25116
rect 34896 25060 34944 25116
rect 35000 25060 35048 25116
rect 35104 25060 35152 25116
rect 35208 25060 35218 25116
rect 0 24276 800 24304
rect 3998 24276 4008 24332
rect 4064 24276 4112 24332
rect 4168 24276 4216 24332
rect 4272 24276 4320 24332
rect 4376 24276 4424 24332
rect 4480 24276 4528 24332
rect 4584 24276 4632 24332
rect 4688 24276 4736 24332
rect 4792 24276 4840 24332
rect 4896 24276 4944 24332
rect 5000 24276 5048 24332
rect 5104 24276 5152 24332
rect 5208 24276 5218 24332
rect 23998 24276 24008 24332
rect 24064 24276 24112 24332
rect 24168 24276 24216 24332
rect 24272 24276 24320 24332
rect 24376 24276 24424 24332
rect 24480 24276 24528 24332
rect 24584 24276 24632 24332
rect 24688 24276 24736 24332
rect 24792 24276 24840 24332
rect 24896 24276 24944 24332
rect 25000 24276 25048 24332
rect 25104 24276 25152 24332
rect 25208 24276 25218 24332
rect 0 24220 1708 24276
rect 1764 24220 1774 24276
rect 0 24192 800 24220
rect 13998 23492 14008 23548
rect 14064 23492 14112 23548
rect 14168 23492 14216 23548
rect 14272 23492 14320 23548
rect 14376 23492 14424 23548
rect 14480 23492 14528 23548
rect 14584 23492 14632 23548
rect 14688 23492 14736 23548
rect 14792 23492 14840 23548
rect 14896 23492 14944 23548
rect 15000 23492 15048 23548
rect 15104 23492 15152 23548
rect 15208 23492 15218 23548
rect 33998 23492 34008 23548
rect 34064 23492 34112 23548
rect 34168 23492 34216 23548
rect 34272 23492 34320 23548
rect 34376 23492 34424 23548
rect 34480 23492 34528 23548
rect 34584 23492 34632 23548
rect 34688 23492 34736 23548
rect 34792 23492 34840 23548
rect 34896 23492 34944 23548
rect 35000 23492 35048 23548
rect 35104 23492 35152 23548
rect 35208 23492 35218 23548
rect 0 22932 800 22960
rect 0 22876 1708 22932
rect 1764 22876 1774 22932
rect 0 22848 800 22876
rect 3998 22708 4008 22764
rect 4064 22708 4112 22764
rect 4168 22708 4216 22764
rect 4272 22708 4320 22764
rect 4376 22708 4424 22764
rect 4480 22708 4528 22764
rect 4584 22708 4632 22764
rect 4688 22708 4736 22764
rect 4792 22708 4840 22764
rect 4896 22708 4944 22764
rect 5000 22708 5048 22764
rect 5104 22708 5152 22764
rect 5208 22708 5218 22764
rect 23998 22708 24008 22764
rect 24064 22708 24112 22764
rect 24168 22708 24216 22764
rect 24272 22708 24320 22764
rect 24376 22708 24424 22764
rect 24480 22708 24528 22764
rect 24584 22708 24632 22764
rect 24688 22708 24736 22764
rect 24792 22708 24840 22764
rect 24896 22708 24944 22764
rect 25000 22708 25048 22764
rect 25104 22708 25152 22764
rect 25208 22708 25218 22764
rect 13998 21924 14008 21980
rect 14064 21924 14112 21980
rect 14168 21924 14216 21980
rect 14272 21924 14320 21980
rect 14376 21924 14424 21980
rect 14480 21924 14528 21980
rect 14584 21924 14632 21980
rect 14688 21924 14736 21980
rect 14792 21924 14840 21980
rect 14896 21924 14944 21980
rect 15000 21924 15048 21980
rect 15104 21924 15152 21980
rect 15208 21924 15218 21980
rect 33998 21924 34008 21980
rect 34064 21924 34112 21980
rect 34168 21924 34216 21980
rect 34272 21924 34320 21980
rect 34376 21924 34424 21980
rect 34480 21924 34528 21980
rect 34584 21924 34632 21980
rect 34688 21924 34736 21980
rect 34792 21924 34840 21980
rect 34896 21924 34944 21980
rect 35000 21924 35048 21980
rect 35104 21924 35152 21980
rect 35208 21924 35218 21980
rect 0 21588 800 21616
rect 0 21532 1708 21588
rect 1764 21532 1774 21588
rect 0 21504 800 21532
rect 3998 21140 4008 21196
rect 4064 21140 4112 21196
rect 4168 21140 4216 21196
rect 4272 21140 4320 21196
rect 4376 21140 4424 21196
rect 4480 21140 4528 21196
rect 4584 21140 4632 21196
rect 4688 21140 4736 21196
rect 4792 21140 4840 21196
rect 4896 21140 4944 21196
rect 5000 21140 5048 21196
rect 5104 21140 5152 21196
rect 5208 21140 5218 21196
rect 23998 21140 24008 21196
rect 24064 21140 24112 21196
rect 24168 21140 24216 21196
rect 24272 21140 24320 21196
rect 24376 21140 24424 21196
rect 24480 21140 24528 21196
rect 24584 21140 24632 21196
rect 24688 21140 24736 21196
rect 24792 21140 24840 21196
rect 24896 21140 24944 21196
rect 25000 21140 25048 21196
rect 25104 21140 25152 21196
rect 25208 21140 25218 21196
rect 13998 20356 14008 20412
rect 14064 20356 14112 20412
rect 14168 20356 14216 20412
rect 14272 20356 14320 20412
rect 14376 20356 14424 20412
rect 14480 20356 14528 20412
rect 14584 20356 14632 20412
rect 14688 20356 14736 20412
rect 14792 20356 14840 20412
rect 14896 20356 14944 20412
rect 15000 20356 15048 20412
rect 15104 20356 15152 20412
rect 15208 20356 15218 20412
rect 33998 20356 34008 20412
rect 34064 20356 34112 20412
rect 34168 20356 34216 20412
rect 34272 20356 34320 20412
rect 34376 20356 34424 20412
rect 34480 20356 34528 20412
rect 34584 20356 34632 20412
rect 34688 20356 34736 20412
rect 34792 20356 34840 20412
rect 34896 20356 34944 20412
rect 35000 20356 35048 20412
rect 35104 20356 35152 20412
rect 35208 20356 35218 20412
rect 0 20244 800 20272
rect 0 20188 1708 20244
rect 1764 20188 1774 20244
rect 0 20160 800 20188
rect 3998 19572 4008 19628
rect 4064 19572 4112 19628
rect 4168 19572 4216 19628
rect 4272 19572 4320 19628
rect 4376 19572 4424 19628
rect 4480 19572 4528 19628
rect 4584 19572 4632 19628
rect 4688 19572 4736 19628
rect 4792 19572 4840 19628
rect 4896 19572 4944 19628
rect 5000 19572 5048 19628
rect 5104 19572 5152 19628
rect 5208 19572 5218 19628
rect 23998 19572 24008 19628
rect 24064 19572 24112 19628
rect 24168 19572 24216 19628
rect 24272 19572 24320 19628
rect 24376 19572 24424 19628
rect 24480 19572 24528 19628
rect 24584 19572 24632 19628
rect 24688 19572 24736 19628
rect 24792 19572 24840 19628
rect 24896 19572 24944 19628
rect 25000 19572 25048 19628
rect 25104 19572 25152 19628
rect 25208 19572 25218 19628
rect 1698 18956 1708 19012
rect 1764 18956 1774 19012
rect 0 18900 800 18928
rect 1708 18900 1764 18956
rect 0 18844 1764 18900
rect 0 18816 800 18844
rect 13998 18788 14008 18844
rect 14064 18788 14112 18844
rect 14168 18788 14216 18844
rect 14272 18788 14320 18844
rect 14376 18788 14424 18844
rect 14480 18788 14528 18844
rect 14584 18788 14632 18844
rect 14688 18788 14736 18844
rect 14792 18788 14840 18844
rect 14896 18788 14944 18844
rect 15000 18788 15048 18844
rect 15104 18788 15152 18844
rect 15208 18788 15218 18844
rect 33998 18788 34008 18844
rect 34064 18788 34112 18844
rect 34168 18788 34216 18844
rect 34272 18788 34320 18844
rect 34376 18788 34424 18844
rect 34480 18788 34528 18844
rect 34584 18788 34632 18844
rect 34688 18788 34736 18844
rect 34792 18788 34840 18844
rect 34896 18788 34944 18844
rect 35000 18788 35048 18844
rect 35104 18788 35152 18844
rect 35208 18788 35218 18844
rect 39200 18676 40000 18704
rect 38210 18620 38220 18676
rect 38276 18620 40000 18676
rect 39200 18592 40000 18620
rect 3998 18004 4008 18060
rect 4064 18004 4112 18060
rect 4168 18004 4216 18060
rect 4272 18004 4320 18060
rect 4376 18004 4424 18060
rect 4480 18004 4528 18060
rect 4584 18004 4632 18060
rect 4688 18004 4736 18060
rect 4792 18004 4840 18060
rect 4896 18004 4944 18060
rect 5000 18004 5048 18060
rect 5104 18004 5152 18060
rect 5208 18004 5218 18060
rect 23998 18004 24008 18060
rect 24064 18004 24112 18060
rect 24168 18004 24216 18060
rect 24272 18004 24320 18060
rect 24376 18004 24424 18060
rect 24480 18004 24528 18060
rect 24584 18004 24632 18060
rect 24688 18004 24736 18060
rect 24792 18004 24840 18060
rect 24896 18004 24944 18060
rect 25000 18004 25048 18060
rect 25104 18004 25152 18060
rect 25208 18004 25218 18060
rect 0 17556 800 17584
rect 0 17500 1708 17556
rect 1764 17500 1774 17556
rect 0 17472 800 17500
rect 13998 17220 14008 17276
rect 14064 17220 14112 17276
rect 14168 17220 14216 17276
rect 14272 17220 14320 17276
rect 14376 17220 14424 17276
rect 14480 17220 14528 17276
rect 14584 17220 14632 17276
rect 14688 17220 14736 17276
rect 14792 17220 14840 17276
rect 14896 17220 14944 17276
rect 15000 17220 15048 17276
rect 15104 17220 15152 17276
rect 15208 17220 15218 17276
rect 33998 17220 34008 17276
rect 34064 17220 34112 17276
rect 34168 17220 34216 17276
rect 34272 17220 34320 17276
rect 34376 17220 34424 17276
rect 34480 17220 34528 17276
rect 34584 17220 34632 17276
rect 34688 17220 34736 17276
rect 34792 17220 34840 17276
rect 34896 17220 34944 17276
rect 35000 17220 35048 17276
rect 35104 17220 35152 17276
rect 35208 17220 35218 17276
rect 3998 16436 4008 16492
rect 4064 16436 4112 16492
rect 4168 16436 4216 16492
rect 4272 16436 4320 16492
rect 4376 16436 4424 16492
rect 4480 16436 4528 16492
rect 4584 16436 4632 16492
rect 4688 16436 4736 16492
rect 4792 16436 4840 16492
rect 4896 16436 4944 16492
rect 5000 16436 5048 16492
rect 5104 16436 5152 16492
rect 5208 16436 5218 16492
rect 23998 16436 24008 16492
rect 24064 16436 24112 16492
rect 24168 16436 24216 16492
rect 24272 16436 24320 16492
rect 24376 16436 24424 16492
rect 24480 16436 24528 16492
rect 24584 16436 24632 16492
rect 24688 16436 24736 16492
rect 24792 16436 24840 16492
rect 24896 16436 24944 16492
rect 25000 16436 25048 16492
rect 25104 16436 25152 16492
rect 25208 16436 25218 16492
rect 0 16212 800 16240
rect 0 16156 1708 16212
rect 1764 16156 1774 16212
rect 0 16128 800 16156
rect 13998 15652 14008 15708
rect 14064 15652 14112 15708
rect 14168 15652 14216 15708
rect 14272 15652 14320 15708
rect 14376 15652 14424 15708
rect 14480 15652 14528 15708
rect 14584 15652 14632 15708
rect 14688 15652 14736 15708
rect 14792 15652 14840 15708
rect 14896 15652 14944 15708
rect 15000 15652 15048 15708
rect 15104 15652 15152 15708
rect 15208 15652 15218 15708
rect 33998 15652 34008 15708
rect 34064 15652 34112 15708
rect 34168 15652 34216 15708
rect 34272 15652 34320 15708
rect 34376 15652 34424 15708
rect 34480 15652 34528 15708
rect 34584 15652 34632 15708
rect 34688 15652 34736 15708
rect 34792 15652 34840 15708
rect 34896 15652 34944 15708
rect 35000 15652 35048 15708
rect 35104 15652 35152 15708
rect 35208 15652 35218 15708
rect 0 14868 800 14896
rect 3998 14868 4008 14924
rect 4064 14868 4112 14924
rect 4168 14868 4216 14924
rect 4272 14868 4320 14924
rect 4376 14868 4424 14924
rect 4480 14868 4528 14924
rect 4584 14868 4632 14924
rect 4688 14868 4736 14924
rect 4792 14868 4840 14924
rect 4896 14868 4944 14924
rect 5000 14868 5048 14924
rect 5104 14868 5152 14924
rect 5208 14868 5218 14924
rect 23998 14868 24008 14924
rect 24064 14868 24112 14924
rect 24168 14868 24216 14924
rect 24272 14868 24320 14924
rect 24376 14868 24424 14924
rect 24480 14868 24528 14924
rect 24584 14868 24632 14924
rect 24688 14868 24736 14924
rect 24792 14868 24840 14924
rect 24896 14868 24944 14924
rect 25000 14868 25048 14924
rect 25104 14868 25152 14924
rect 25208 14868 25218 14924
rect 0 14812 1708 14868
rect 1764 14812 1774 14868
rect 0 14784 800 14812
rect 13998 14084 14008 14140
rect 14064 14084 14112 14140
rect 14168 14084 14216 14140
rect 14272 14084 14320 14140
rect 14376 14084 14424 14140
rect 14480 14084 14528 14140
rect 14584 14084 14632 14140
rect 14688 14084 14736 14140
rect 14792 14084 14840 14140
rect 14896 14084 14944 14140
rect 15000 14084 15048 14140
rect 15104 14084 15152 14140
rect 15208 14084 15218 14140
rect 33998 14084 34008 14140
rect 34064 14084 34112 14140
rect 34168 14084 34216 14140
rect 34272 14084 34320 14140
rect 34376 14084 34424 14140
rect 34480 14084 34528 14140
rect 34584 14084 34632 14140
rect 34688 14084 34736 14140
rect 34792 14084 34840 14140
rect 34896 14084 34944 14140
rect 35000 14084 35048 14140
rect 35104 14084 35152 14140
rect 35208 14084 35218 14140
rect 0 13524 800 13552
rect 0 13468 1708 13524
rect 1764 13468 1774 13524
rect 0 13440 800 13468
rect 3998 13300 4008 13356
rect 4064 13300 4112 13356
rect 4168 13300 4216 13356
rect 4272 13300 4320 13356
rect 4376 13300 4424 13356
rect 4480 13300 4528 13356
rect 4584 13300 4632 13356
rect 4688 13300 4736 13356
rect 4792 13300 4840 13356
rect 4896 13300 4944 13356
rect 5000 13300 5048 13356
rect 5104 13300 5152 13356
rect 5208 13300 5218 13356
rect 23998 13300 24008 13356
rect 24064 13300 24112 13356
rect 24168 13300 24216 13356
rect 24272 13300 24320 13356
rect 24376 13300 24424 13356
rect 24480 13300 24528 13356
rect 24584 13300 24632 13356
rect 24688 13300 24736 13356
rect 24792 13300 24840 13356
rect 24896 13300 24944 13356
rect 25000 13300 25048 13356
rect 25104 13300 25152 13356
rect 25208 13300 25218 13356
rect 13998 12516 14008 12572
rect 14064 12516 14112 12572
rect 14168 12516 14216 12572
rect 14272 12516 14320 12572
rect 14376 12516 14424 12572
rect 14480 12516 14528 12572
rect 14584 12516 14632 12572
rect 14688 12516 14736 12572
rect 14792 12516 14840 12572
rect 14896 12516 14944 12572
rect 15000 12516 15048 12572
rect 15104 12516 15152 12572
rect 15208 12516 15218 12572
rect 33998 12516 34008 12572
rect 34064 12516 34112 12572
rect 34168 12516 34216 12572
rect 34272 12516 34320 12572
rect 34376 12516 34424 12572
rect 34480 12516 34528 12572
rect 34584 12516 34632 12572
rect 34688 12516 34736 12572
rect 34792 12516 34840 12572
rect 34896 12516 34944 12572
rect 35000 12516 35048 12572
rect 35104 12516 35152 12572
rect 35208 12516 35218 12572
rect 0 12180 800 12208
rect 0 12124 1708 12180
rect 1764 12124 1774 12180
rect 0 12096 800 12124
rect 3998 11732 4008 11788
rect 4064 11732 4112 11788
rect 4168 11732 4216 11788
rect 4272 11732 4320 11788
rect 4376 11732 4424 11788
rect 4480 11732 4528 11788
rect 4584 11732 4632 11788
rect 4688 11732 4736 11788
rect 4792 11732 4840 11788
rect 4896 11732 4944 11788
rect 5000 11732 5048 11788
rect 5104 11732 5152 11788
rect 5208 11732 5218 11788
rect 23998 11732 24008 11788
rect 24064 11732 24112 11788
rect 24168 11732 24216 11788
rect 24272 11732 24320 11788
rect 24376 11732 24424 11788
rect 24480 11732 24528 11788
rect 24584 11732 24632 11788
rect 24688 11732 24736 11788
rect 24792 11732 24840 11788
rect 24896 11732 24944 11788
rect 25000 11732 25048 11788
rect 25104 11732 25152 11788
rect 25208 11732 25218 11788
rect 13998 10948 14008 11004
rect 14064 10948 14112 11004
rect 14168 10948 14216 11004
rect 14272 10948 14320 11004
rect 14376 10948 14424 11004
rect 14480 10948 14528 11004
rect 14584 10948 14632 11004
rect 14688 10948 14736 11004
rect 14792 10948 14840 11004
rect 14896 10948 14944 11004
rect 15000 10948 15048 11004
rect 15104 10948 15152 11004
rect 15208 10948 15218 11004
rect 33998 10948 34008 11004
rect 34064 10948 34112 11004
rect 34168 10948 34216 11004
rect 34272 10948 34320 11004
rect 34376 10948 34424 11004
rect 34480 10948 34528 11004
rect 34584 10948 34632 11004
rect 34688 10948 34736 11004
rect 34792 10948 34840 11004
rect 34896 10948 34944 11004
rect 35000 10948 35048 11004
rect 35104 10948 35152 11004
rect 35208 10948 35218 11004
rect 0 10836 800 10864
rect 0 10780 1708 10836
rect 1764 10780 1774 10836
rect 0 10752 800 10780
rect 10322 10556 10332 10612
rect 10388 10556 11900 10612
rect 11956 10556 11966 10612
rect 12114 10556 12124 10612
rect 12180 10556 12908 10612
rect 12964 10556 12974 10612
rect 12908 10500 12964 10556
rect 10770 10444 10780 10500
rect 10836 10444 12012 10500
rect 12068 10444 12078 10500
rect 12908 10444 37436 10500
rect 37492 10444 37502 10500
rect 3998 10164 4008 10220
rect 4064 10164 4112 10220
rect 4168 10164 4216 10220
rect 4272 10164 4320 10220
rect 4376 10164 4424 10220
rect 4480 10164 4528 10220
rect 4584 10164 4632 10220
rect 4688 10164 4736 10220
rect 4792 10164 4840 10220
rect 4896 10164 4944 10220
rect 5000 10164 5048 10220
rect 5104 10164 5152 10220
rect 5208 10164 5218 10220
rect 23998 10164 24008 10220
rect 24064 10164 24112 10220
rect 24168 10164 24216 10220
rect 24272 10164 24320 10220
rect 24376 10164 24424 10220
rect 24480 10164 24528 10220
rect 24584 10164 24632 10220
rect 24688 10164 24736 10220
rect 24792 10164 24840 10220
rect 24896 10164 24944 10220
rect 25000 10164 25048 10220
rect 25104 10164 25152 10220
rect 25208 10164 25218 10220
rect 7746 9660 7756 9716
rect 7812 9660 8316 9716
rect 8372 9660 37884 9716
rect 37940 9660 37950 9716
rect 1698 9548 1708 9604
rect 1764 9548 1774 9604
rect 0 9492 800 9520
rect 1708 9492 1764 9548
rect 0 9436 1764 9492
rect 0 9408 800 9436
rect 13998 9380 14008 9436
rect 14064 9380 14112 9436
rect 14168 9380 14216 9436
rect 14272 9380 14320 9436
rect 14376 9380 14424 9436
rect 14480 9380 14528 9436
rect 14584 9380 14632 9436
rect 14688 9380 14736 9436
rect 14792 9380 14840 9436
rect 14896 9380 14944 9436
rect 15000 9380 15048 9436
rect 15104 9380 15152 9436
rect 15208 9380 15218 9436
rect 33998 9380 34008 9436
rect 34064 9380 34112 9436
rect 34168 9380 34216 9436
rect 34272 9380 34320 9436
rect 34376 9380 34424 9436
rect 34480 9380 34528 9436
rect 34584 9380 34632 9436
rect 34688 9380 34736 9436
rect 34792 9380 34840 9436
rect 34896 9380 34944 9436
rect 35000 9380 35048 9436
rect 35104 9380 35152 9436
rect 35208 9380 35218 9436
rect 8866 8876 8876 8932
rect 8932 8876 9660 8932
rect 9716 8876 12684 8932
rect 12740 8876 12750 8932
rect 7382 8652 7420 8708
rect 7476 8652 7868 8708
rect 7924 8652 7934 8708
rect 3998 8596 4008 8652
rect 4064 8596 4112 8652
rect 4168 8596 4216 8652
rect 4272 8596 4320 8652
rect 4376 8596 4424 8652
rect 4480 8596 4528 8652
rect 4584 8596 4632 8652
rect 4688 8596 4736 8652
rect 4792 8596 4840 8652
rect 4896 8596 4944 8652
rect 5000 8596 5048 8652
rect 5104 8596 5152 8652
rect 5208 8596 5218 8652
rect 23998 8596 24008 8652
rect 24064 8596 24112 8652
rect 24168 8596 24216 8652
rect 24272 8596 24320 8652
rect 24376 8596 24424 8652
rect 24480 8596 24528 8652
rect 24584 8596 24632 8652
rect 24688 8596 24736 8652
rect 24792 8596 24840 8652
rect 24896 8596 24944 8652
rect 25000 8596 25048 8652
rect 25104 8596 25152 8652
rect 25208 8596 25218 8652
rect 7186 8540 7196 8596
rect 7252 8540 9772 8596
rect 9828 8540 13468 8596
rect 13524 8540 13534 8596
rect 7410 8316 7420 8372
rect 7476 8316 7756 8372
rect 7812 8316 37884 8372
rect 37940 8316 37950 8372
rect 5618 8204 5628 8260
rect 5684 8204 5964 8260
rect 6020 8204 6030 8260
rect 8194 8204 8204 8260
rect 8260 8204 8764 8260
rect 8820 8204 11564 8260
rect 11620 8204 11630 8260
rect 0 8148 800 8176
rect 0 8092 1708 8148
rect 1764 8092 1774 8148
rect 9314 8092 9324 8148
rect 9380 8092 14252 8148
rect 14308 8092 14318 8148
rect 0 8064 800 8092
rect 6486 7980 6524 8036
rect 6580 7980 6590 8036
rect 6934 7980 6972 8036
rect 7028 7980 7038 8036
rect 8306 7980 8316 8036
rect 8372 7980 8988 8036
rect 9044 7980 9054 8036
rect 16482 7980 16492 8036
rect 16548 7980 28364 8036
rect 28420 7980 28430 8036
rect 13998 7812 14008 7868
rect 14064 7812 14112 7868
rect 14168 7812 14216 7868
rect 14272 7812 14320 7868
rect 14376 7812 14424 7868
rect 14480 7812 14528 7868
rect 14584 7812 14632 7868
rect 14688 7812 14736 7868
rect 14792 7812 14840 7868
rect 14896 7812 14944 7868
rect 15000 7812 15048 7868
rect 15104 7812 15152 7868
rect 15208 7812 15218 7868
rect 16492 7700 16548 7980
rect 33998 7812 34008 7868
rect 34064 7812 34112 7868
rect 34168 7812 34216 7868
rect 34272 7812 34320 7868
rect 34376 7812 34424 7868
rect 34480 7812 34528 7868
rect 34584 7812 34632 7868
rect 34688 7812 34736 7868
rect 34792 7812 34840 7868
rect 34896 7812 34944 7868
rect 35000 7812 35048 7868
rect 35104 7812 35152 7868
rect 35208 7812 35218 7868
rect 5954 7644 5964 7700
rect 6020 7644 7980 7700
rect 8036 7644 8046 7700
rect 14690 7644 14700 7700
rect 14756 7644 16548 7700
rect 6514 7532 6524 7588
rect 6580 7532 10108 7588
rect 10164 7532 10174 7588
rect 13794 7532 13804 7588
rect 13860 7532 17612 7588
rect 17668 7532 17678 7588
rect 7074 7420 7084 7476
rect 7140 7420 7756 7476
rect 7812 7420 7822 7476
rect 8194 7420 8204 7476
rect 8260 7420 8652 7476
rect 8708 7420 8718 7476
rect 11554 7420 11564 7476
rect 11620 7420 14700 7476
rect 14756 7420 14766 7476
rect 6402 7308 6412 7364
rect 6468 7308 7980 7364
rect 8036 7308 8046 7364
rect 8306 7308 8316 7364
rect 8372 7308 10444 7364
rect 10500 7308 10510 7364
rect 12898 7308 12908 7364
rect 12964 7308 13692 7364
rect 13748 7308 13758 7364
rect 2930 7196 2940 7252
rect 2996 7196 4284 7252
rect 4340 7196 5796 7252
rect 5740 7140 5796 7196
rect 5730 7084 5740 7140
rect 5796 7084 5806 7140
rect 10770 7084 10780 7140
rect 10836 7084 11676 7140
rect 11732 7084 13580 7140
rect 13636 7084 13804 7140
rect 13860 7084 13870 7140
rect 3998 7028 4008 7084
rect 4064 7028 4112 7084
rect 4168 7028 4216 7084
rect 4272 7028 4320 7084
rect 4376 7028 4424 7084
rect 4480 7028 4528 7084
rect 4584 7028 4632 7084
rect 4688 7028 4736 7084
rect 4792 7028 4840 7084
rect 4896 7028 4944 7084
rect 5000 7028 5048 7084
rect 5104 7028 5152 7084
rect 5208 7028 5218 7084
rect 23998 7028 24008 7084
rect 24064 7028 24112 7084
rect 24168 7028 24216 7084
rect 24272 7028 24320 7084
rect 24376 7028 24424 7084
rect 24480 7028 24528 7084
rect 24584 7028 24632 7084
rect 24688 7028 24736 7084
rect 24792 7028 24840 7084
rect 24896 7028 24944 7084
rect 25000 7028 25048 7084
rect 25104 7028 25152 7084
rect 25208 7028 25218 7084
rect 6738 6860 6748 6916
rect 6804 6860 7420 6916
rect 7476 6860 7486 6916
rect 0 6804 800 6832
rect 0 6748 1932 6804
rect 1988 6748 1998 6804
rect 0 6720 800 6748
rect 7942 6636 7980 6692
rect 8036 6636 8046 6692
rect 10770 6636 10780 6692
rect 10836 6636 13468 6692
rect 13524 6636 13534 6692
rect 20514 6636 20524 6692
rect 20580 6636 21420 6692
rect 21476 6636 36428 6692
rect 36484 6636 36494 6692
rect 6300 6524 8652 6580
rect 8708 6524 9436 6580
rect 9492 6524 9502 6580
rect 12114 6524 12124 6580
rect 12180 6524 13356 6580
rect 13412 6524 15148 6580
rect 15204 6524 17388 6580
rect 17444 6524 19740 6580
rect 19796 6524 20748 6580
rect 20804 6524 20814 6580
rect 6300 6468 6356 6524
rect 12124 6468 12180 6524
rect 2258 6412 2268 6468
rect 2324 6412 5516 6468
rect 5572 6412 5582 6468
rect 6290 6412 6300 6468
rect 6356 6412 6366 6468
rect 6626 6412 6636 6468
rect 6692 6412 7868 6468
rect 7924 6412 7934 6468
rect 8194 6412 8204 6468
rect 8260 6412 12180 6468
rect 8204 6356 8260 6412
rect 39200 6356 40000 6384
rect 3490 6300 3500 6356
rect 3556 6300 3948 6356
rect 4004 6300 5852 6356
rect 5908 6300 7420 6356
rect 7476 6300 8260 6356
rect 37650 6300 37660 6356
rect 37716 6300 38220 6356
rect 38276 6300 40000 6356
rect 13998 6244 14008 6300
rect 14064 6244 14112 6300
rect 14168 6244 14216 6300
rect 14272 6244 14320 6300
rect 14376 6244 14424 6300
rect 14480 6244 14528 6300
rect 14584 6244 14632 6300
rect 14688 6244 14736 6300
rect 14792 6244 14840 6300
rect 14896 6244 14944 6300
rect 15000 6244 15048 6300
rect 15104 6244 15152 6300
rect 15208 6244 15218 6300
rect 33998 6244 34008 6300
rect 34064 6244 34112 6300
rect 34168 6244 34216 6300
rect 34272 6244 34320 6300
rect 34376 6244 34424 6300
rect 34480 6244 34528 6300
rect 34584 6244 34632 6300
rect 34688 6244 34736 6300
rect 34792 6244 34840 6300
rect 34896 6244 34944 6300
rect 35000 6244 35048 6300
rect 35104 6244 35152 6300
rect 35208 6244 35218 6300
rect 39200 6272 40000 6300
rect 6150 6188 6188 6244
rect 6244 6188 6254 6244
rect 6850 6188 6860 6244
rect 6916 6188 7084 6244
rect 7140 6188 7150 6244
rect 7298 6188 7308 6244
rect 7364 6188 7756 6244
rect 7812 6188 7822 6244
rect 7970 6188 7980 6244
rect 8036 6188 8046 6244
rect 7980 6132 8036 6188
rect 2594 6076 2604 6132
rect 2660 6076 8036 6132
rect 8978 6076 8988 6132
rect 9044 6076 10220 6132
rect 10276 6076 11452 6132
rect 11508 6076 11518 6132
rect 4722 5964 4732 6020
rect 4788 5964 5516 6020
rect 5572 5964 5582 6020
rect 5730 5964 5740 6020
rect 5796 5964 7084 6020
rect 7140 5964 7150 6020
rect 7634 5964 7644 6020
rect 7700 5964 11788 6020
rect 11844 5964 11854 6020
rect 1922 5852 1932 5908
rect 1988 5852 7756 5908
rect 7812 5852 7822 5908
rect 8530 5852 8540 5908
rect 8596 5852 11564 5908
rect 11620 5852 11630 5908
rect 14802 5852 14812 5908
rect 14868 5852 15372 5908
rect 15428 5852 16380 5908
rect 16436 5852 16446 5908
rect 4722 5740 4732 5796
rect 4788 5740 6076 5796
rect 6132 5740 6142 5796
rect 13794 5740 13804 5796
rect 13860 5740 16156 5796
rect 16212 5740 16222 5796
rect 5618 5628 5628 5684
rect 5684 5628 7084 5684
rect 7140 5628 7150 5684
rect 0 5460 800 5488
rect 3998 5460 4008 5516
rect 4064 5460 4112 5516
rect 4168 5460 4216 5516
rect 4272 5460 4320 5516
rect 4376 5460 4424 5516
rect 4480 5460 4528 5516
rect 4584 5460 4632 5516
rect 4688 5460 4736 5516
rect 4792 5460 4840 5516
rect 4896 5460 4944 5516
rect 5000 5460 5048 5516
rect 5104 5460 5152 5516
rect 5208 5460 5218 5516
rect 23998 5460 24008 5516
rect 24064 5460 24112 5516
rect 24168 5460 24216 5516
rect 24272 5460 24320 5516
rect 24376 5460 24424 5516
rect 24480 5460 24528 5516
rect 24584 5460 24632 5516
rect 24688 5460 24736 5516
rect 24792 5460 24840 5516
rect 24896 5460 24944 5516
rect 25000 5460 25048 5516
rect 25104 5460 25152 5516
rect 25208 5460 25218 5516
rect 0 5404 2212 5460
rect 0 5376 800 5404
rect 2156 5348 2212 5404
rect 2146 5292 2156 5348
rect 2212 5292 2222 5348
rect 3714 5292 3724 5348
rect 3780 5292 5404 5348
rect 5460 5292 5470 5348
rect 9650 5292 9660 5348
rect 9716 5292 12236 5348
rect 12292 5292 12302 5348
rect 4610 5180 4620 5236
rect 4676 5180 5516 5236
rect 5572 5180 5582 5236
rect 8866 5180 8876 5236
rect 8932 5180 13580 5236
rect 13636 5180 13646 5236
rect 2482 5068 2492 5124
rect 2548 5068 3052 5124
rect 3108 5068 4060 5124
rect 4116 5068 4126 5124
rect 4386 5068 4396 5124
rect 4452 5068 6188 5124
rect 6244 5068 6254 5124
rect 8642 5068 8652 5124
rect 8708 5068 11228 5124
rect 11284 5068 11294 5124
rect 16258 5068 16268 5124
rect 16324 5068 17500 5124
rect 17556 5068 17566 5124
rect 5618 4956 5628 5012
rect 5684 4956 5694 5012
rect 5842 4956 5852 5012
rect 5908 4956 6412 5012
rect 6468 4956 6478 5012
rect 10210 4956 10220 5012
rect 10276 4956 10892 5012
rect 10948 4956 10958 5012
rect 13570 4956 13580 5012
rect 13636 4956 13916 5012
rect 13972 4956 13982 5012
rect 16482 4956 16492 5012
rect 16548 4956 17052 5012
rect 17108 4956 17118 5012
rect 23650 4956 23660 5012
rect 23716 4956 24892 5012
rect 24948 4956 24958 5012
rect 30818 4956 30828 5012
rect 30884 4956 32844 5012
rect 32900 4956 32910 5012
rect 5628 4900 5684 4956
rect 5058 4844 5068 4900
rect 5124 4844 5684 4900
rect 6178 4844 6188 4900
rect 6244 4844 6254 4900
rect 6850 4844 6860 4900
rect 6916 4844 7980 4900
rect 8036 4844 8046 4900
rect 9426 4844 9436 4900
rect 9492 4844 12460 4900
rect 12516 4844 12526 4900
rect 13804 4844 16044 4900
rect 16100 4844 16110 4900
rect 16370 4844 16380 4900
rect 16436 4844 16716 4900
rect 16772 4844 16782 4900
rect 33852 4844 34412 4900
rect 34468 4844 34478 4900
rect 6188 4788 6244 4844
rect 6188 4732 9884 4788
rect 9940 4732 12572 4788
rect 12628 4732 12638 4788
rect 13804 4676 13860 4844
rect 15670 4732 15708 4788
rect 15764 4732 15774 4788
rect 13998 4676 14008 4732
rect 14064 4676 14112 4732
rect 14168 4676 14216 4732
rect 14272 4676 14320 4732
rect 14376 4676 14424 4732
rect 14480 4676 14528 4732
rect 14584 4676 14632 4732
rect 14688 4676 14736 4732
rect 14792 4676 14840 4732
rect 14896 4676 14944 4732
rect 15000 4676 15048 4732
rect 15104 4676 15152 4732
rect 15208 4676 15218 4732
rect 4946 4620 4956 4676
rect 5012 4620 7308 4676
rect 7364 4620 7374 4676
rect 10210 4620 10220 4676
rect 10276 4620 13860 4676
rect 6290 4508 6300 4564
rect 6356 4508 6860 4564
rect 6916 4508 6926 4564
rect 14802 4508 14812 4564
rect 14868 4508 15484 4564
rect 15540 4508 15550 4564
rect 15698 4508 15708 4564
rect 15764 4508 16380 4564
rect 16436 4508 16446 4564
rect 24098 4508 24108 4564
rect 24164 4508 25340 4564
rect 25396 4508 25406 4564
rect 1698 4396 1708 4452
rect 1764 4396 1774 4452
rect 2034 4396 2044 4452
rect 2100 4396 3836 4452
rect 3892 4396 3902 4452
rect 13570 4396 13580 4452
rect 13636 4396 19908 4452
rect 20066 4396 20076 4452
rect 20132 4396 20860 4452
rect 20916 4396 20926 4452
rect 26852 4396 31948 4452
rect 0 4116 800 4144
rect 1708 4116 1764 4396
rect 19852 4340 19908 4396
rect 26852 4340 26908 4396
rect 6402 4284 6412 4340
rect 6468 4284 12012 4340
rect 12068 4284 12078 4340
rect 19852 4284 26908 4340
rect 31892 4340 31948 4396
rect 33852 4340 33908 4844
rect 33998 4676 34008 4732
rect 34064 4676 34112 4732
rect 34168 4676 34216 4732
rect 34272 4676 34320 4732
rect 34376 4676 34424 4732
rect 34480 4676 34528 4732
rect 34584 4676 34632 4732
rect 34688 4676 34736 4732
rect 34792 4676 34840 4732
rect 34896 4676 34944 4732
rect 35000 4676 35048 4732
rect 35104 4676 35152 4732
rect 35208 4676 35218 4732
rect 31892 4284 32060 4340
rect 32116 4284 32126 4340
rect 33170 4284 33180 4340
rect 33236 4284 33964 4340
rect 34020 4284 34030 4340
rect 34402 4284 34412 4340
rect 34468 4284 35756 4340
rect 35812 4284 35822 4340
rect 3332 4172 8428 4228
rect 8484 4172 12348 4228
rect 12404 4172 12414 4228
rect 16706 4172 16716 4228
rect 16772 4172 35644 4228
rect 35700 4172 35710 4228
rect 3332 4116 3388 4172
rect 0 4060 1764 4116
rect 3042 4060 3052 4116
rect 3108 4060 3388 4116
rect 3602 4060 3612 4116
rect 3668 4060 4844 4116
rect 4900 4060 5404 4116
rect 5460 4060 6860 4116
rect 6916 4060 6926 4116
rect 7868 4060 9884 4116
rect 9940 4060 10668 4116
rect 10724 4060 10734 4116
rect 13682 4060 13692 4116
rect 13748 4060 14700 4116
rect 14756 4060 22764 4116
rect 22820 4060 22830 4116
rect 23426 4060 23436 4116
rect 23492 4060 24556 4116
rect 24612 4060 24622 4116
rect 26852 4060 37212 4116
rect 37268 4060 37278 4116
rect 0 4032 800 4060
rect 7868 4004 7924 4060
rect 5852 3948 7924 4004
rect 8082 3948 8092 4004
rect 8148 3948 15708 4004
rect 15764 3948 15774 4004
rect 3998 3892 4008 3948
rect 4064 3892 4112 3948
rect 4168 3892 4216 3948
rect 4272 3892 4320 3948
rect 4376 3892 4424 3948
rect 4480 3892 4528 3948
rect 4584 3892 4632 3948
rect 4688 3892 4736 3948
rect 4792 3892 4840 3948
rect 4896 3892 4944 3948
rect 5000 3892 5048 3948
rect 5104 3892 5152 3948
rect 5208 3892 5218 3948
rect 5852 3780 5908 3948
rect 23998 3892 24008 3948
rect 24064 3892 24112 3948
rect 24168 3892 24216 3948
rect 24272 3892 24320 3948
rect 24376 3892 24424 3948
rect 24480 3892 24528 3948
rect 24584 3892 24632 3948
rect 24688 3892 24736 3948
rect 24792 3892 24840 3948
rect 24896 3892 24944 3948
rect 25000 3892 25048 3948
rect 25104 3892 25152 3948
rect 25208 3892 25218 3948
rect 6066 3836 6076 3892
rect 6132 3836 10108 3892
rect 10164 3836 10174 3892
rect 16930 3836 16940 3892
rect 16996 3836 17724 3892
rect 17780 3836 18900 3892
rect 18844 3780 18900 3836
rect 26852 3780 26908 4060
rect 4274 3724 4284 3780
rect 4340 3724 5908 3780
rect 6486 3724 6524 3780
rect 6580 3724 6590 3780
rect 7858 3724 7868 3780
rect 7924 3724 8316 3780
rect 8372 3724 9884 3780
rect 9940 3724 9950 3780
rect 12562 3724 12572 3780
rect 12628 3724 14028 3780
rect 14084 3724 18620 3780
rect 18676 3724 18686 3780
rect 18844 3724 26908 3780
rect 3490 3612 3500 3668
rect 3556 3612 4060 3668
rect 4116 3612 4126 3668
rect 8316 3612 9996 3668
rect 10052 3612 10062 3668
rect 10546 3612 10556 3668
rect 10612 3612 13020 3668
rect 13076 3612 13086 3668
rect 25106 3612 25116 3668
rect 25172 3612 27692 3668
rect 27748 3612 27758 3668
rect 33618 3612 33628 3668
rect 33684 3612 35308 3668
rect 35364 3612 35374 3668
rect 8316 3556 8372 3612
rect 3938 3500 3948 3556
rect 4004 3500 5180 3556
rect 5236 3500 5246 3556
rect 5730 3500 5740 3556
rect 5796 3500 6972 3556
rect 7028 3500 7038 3556
rect 7410 3500 7420 3556
rect 7476 3500 8372 3556
rect 9762 3500 9772 3556
rect 9828 3500 11452 3556
rect 11508 3500 11518 3556
rect 11666 3500 11676 3556
rect 11732 3500 15260 3556
rect 15316 3500 15326 3556
rect 27570 3500 27580 3556
rect 27636 3500 28588 3556
rect 28644 3500 28654 3556
rect 4946 3388 4956 3444
rect 5012 3388 11228 3444
rect 11284 3388 11294 3444
rect 12450 3388 12460 3444
rect 12516 3388 14812 3444
rect 14868 3388 14878 3444
rect 24546 3388 24556 3444
rect 24612 3388 25788 3444
rect 25844 3388 25854 3444
rect 26674 3388 26684 3444
rect 26740 3388 27132 3444
rect 27188 3388 27198 3444
rect 28466 3388 28476 3444
rect 28532 3388 29036 3444
rect 29092 3388 29484 3444
rect 29540 3388 29550 3444
rect 33842 3388 33852 3444
rect 33908 3388 34524 3444
rect 34580 3388 34590 3444
rect 35298 3388 35308 3444
rect 35364 3388 36204 3444
rect 36260 3388 36270 3444
rect 6962 3276 6972 3332
rect 7028 3276 7084 3332
rect 7140 3276 7150 3332
rect 13998 3108 14008 3164
rect 14064 3108 14112 3164
rect 14168 3108 14216 3164
rect 14272 3108 14320 3164
rect 14376 3108 14424 3164
rect 14480 3108 14528 3164
rect 14584 3108 14632 3164
rect 14688 3108 14736 3164
rect 14792 3108 14840 3164
rect 14896 3108 14944 3164
rect 15000 3108 15048 3164
rect 15104 3108 15152 3164
rect 15208 3108 15218 3164
rect 33998 3108 34008 3164
rect 34064 3108 34112 3164
rect 34168 3108 34216 3164
rect 34272 3108 34320 3164
rect 34376 3108 34424 3164
rect 34480 3108 34528 3164
rect 34584 3108 34632 3164
rect 34688 3108 34736 3164
rect 34792 3108 34840 3164
rect 34896 3108 34944 3164
rect 35000 3108 35048 3164
rect 35104 3108 35152 3164
rect 35208 3108 35218 3164
rect 0 2772 800 2800
rect 0 2716 2156 2772
rect 2212 2716 2222 2772
rect 0 2688 800 2716
rect 6514 924 6524 980
rect 6580 924 7868 980
rect 7924 924 7934 980
<< via3 >>
rect 4008 46228 4064 46284
rect 4112 46228 4168 46284
rect 4216 46228 4272 46284
rect 4320 46228 4376 46284
rect 4424 46228 4480 46284
rect 4528 46228 4584 46284
rect 4632 46228 4688 46284
rect 4736 46228 4792 46284
rect 4840 46228 4896 46284
rect 4944 46228 5000 46284
rect 5048 46228 5104 46284
rect 5152 46228 5208 46284
rect 24008 46228 24064 46284
rect 24112 46228 24168 46284
rect 24216 46228 24272 46284
rect 24320 46228 24376 46284
rect 24424 46228 24480 46284
rect 24528 46228 24584 46284
rect 24632 46228 24688 46284
rect 24736 46228 24792 46284
rect 24840 46228 24896 46284
rect 24944 46228 25000 46284
rect 25048 46228 25104 46284
rect 25152 46228 25208 46284
rect 14008 45444 14064 45500
rect 14112 45444 14168 45500
rect 14216 45444 14272 45500
rect 14320 45444 14376 45500
rect 14424 45444 14480 45500
rect 14528 45444 14584 45500
rect 14632 45444 14688 45500
rect 14736 45444 14792 45500
rect 14840 45444 14896 45500
rect 14944 45444 15000 45500
rect 15048 45444 15104 45500
rect 15152 45444 15208 45500
rect 34008 45444 34064 45500
rect 34112 45444 34168 45500
rect 34216 45444 34272 45500
rect 34320 45444 34376 45500
rect 34424 45444 34480 45500
rect 34528 45444 34584 45500
rect 34632 45444 34688 45500
rect 34736 45444 34792 45500
rect 34840 45444 34896 45500
rect 34944 45444 35000 45500
rect 35048 45444 35104 45500
rect 35152 45444 35208 45500
rect 4008 44660 4064 44716
rect 4112 44660 4168 44716
rect 4216 44660 4272 44716
rect 4320 44660 4376 44716
rect 4424 44660 4480 44716
rect 4528 44660 4584 44716
rect 4632 44660 4688 44716
rect 4736 44660 4792 44716
rect 4840 44660 4896 44716
rect 4944 44660 5000 44716
rect 5048 44660 5104 44716
rect 5152 44660 5208 44716
rect 24008 44660 24064 44716
rect 24112 44660 24168 44716
rect 24216 44660 24272 44716
rect 24320 44660 24376 44716
rect 24424 44660 24480 44716
rect 24528 44660 24584 44716
rect 24632 44660 24688 44716
rect 24736 44660 24792 44716
rect 24840 44660 24896 44716
rect 24944 44660 25000 44716
rect 25048 44660 25104 44716
rect 25152 44660 25208 44716
rect 14008 43876 14064 43932
rect 14112 43876 14168 43932
rect 14216 43876 14272 43932
rect 14320 43876 14376 43932
rect 14424 43876 14480 43932
rect 14528 43876 14584 43932
rect 14632 43876 14688 43932
rect 14736 43876 14792 43932
rect 14840 43876 14896 43932
rect 14944 43876 15000 43932
rect 15048 43876 15104 43932
rect 15152 43876 15208 43932
rect 34008 43876 34064 43932
rect 34112 43876 34168 43932
rect 34216 43876 34272 43932
rect 34320 43876 34376 43932
rect 34424 43876 34480 43932
rect 34528 43876 34584 43932
rect 34632 43876 34688 43932
rect 34736 43876 34792 43932
rect 34840 43876 34896 43932
rect 34944 43876 35000 43932
rect 35048 43876 35104 43932
rect 35152 43876 35208 43932
rect 4008 43092 4064 43148
rect 4112 43092 4168 43148
rect 4216 43092 4272 43148
rect 4320 43092 4376 43148
rect 4424 43092 4480 43148
rect 4528 43092 4584 43148
rect 4632 43092 4688 43148
rect 4736 43092 4792 43148
rect 4840 43092 4896 43148
rect 4944 43092 5000 43148
rect 5048 43092 5104 43148
rect 5152 43092 5208 43148
rect 24008 43092 24064 43148
rect 24112 43092 24168 43148
rect 24216 43092 24272 43148
rect 24320 43092 24376 43148
rect 24424 43092 24480 43148
rect 24528 43092 24584 43148
rect 24632 43092 24688 43148
rect 24736 43092 24792 43148
rect 24840 43092 24896 43148
rect 24944 43092 25000 43148
rect 25048 43092 25104 43148
rect 25152 43092 25208 43148
rect 14008 42308 14064 42364
rect 14112 42308 14168 42364
rect 14216 42308 14272 42364
rect 14320 42308 14376 42364
rect 14424 42308 14480 42364
rect 14528 42308 14584 42364
rect 14632 42308 14688 42364
rect 14736 42308 14792 42364
rect 14840 42308 14896 42364
rect 14944 42308 15000 42364
rect 15048 42308 15104 42364
rect 15152 42308 15208 42364
rect 34008 42308 34064 42364
rect 34112 42308 34168 42364
rect 34216 42308 34272 42364
rect 34320 42308 34376 42364
rect 34424 42308 34480 42364
rect 34528 42308 34584 42364
rect 34632 42308 34688 42364
rect 34736 42308 34792 42364
rect 34840 42308 34896 42364
rect 34944 42308 35000 42364
rect 35048 42308 35104 42364
rect 35152 42308 35208 42364
rect 4008 41524 4064 41580
rect 4112 41524 4168 41580
rect 4216 41524 4272 41580
rect 4320 41524 4376 41580
rect 4424 41524 4480 41580
rect 4528 41524 4584 41580
rect 4632 41524 4688 41580
rect 4736 41524 4792 41580
rect 4840 41524 4896 41580
rect 4944 41524 5000 41580
rect 5048 41524 5104 41580
rect 5152 41524 5208 41580
rect 24008 41524 24064 41580
rect 24112 41524 24168 41580
rect 24216 41524 24272 41580
rect 24320 41524 24376 41580
rect 24424 41524 24480 41580
rect 24528 41524 24584 41580
rect 24632 41524 24688 41580
rect 24736 41524 24792 41580
rect 24840 41524 24896 41580
rect 24944 41524 25000 41580
rect 25048 41524 25104 41580
rect 25152 41524 25208 41580
rect 14008 40740 14064 40796
rect 14112 40740 14168 40796
rect 14216 40740 14272 40796
rect 14320 40740 14376 40796
rect 14424 40740 14480 40796
rect 14528 40740 14584 40796
rect 14632 40740 14688 40796
rect 14736 40740 14792 40796
rect 14840 40740 14896 40796
rect 14944 40740 15000 40796
rect 15048 40740 15104 40796
rect 15152 40740 15208 40796
rect 34008 40740 34064 40796
rect 34112 40740 34168 40796
rect 34216 40740 34272 40796
rect 34320 40740 34376 40796
rect 34424 40740 34480 40796
rect 34528 40740 34584 40796
rect 34632 40740 34688 40796
rect 34736 40740 34792 40796
rect 34840 40740 34896 40796
rect 34944 40740 35000 40796
rect 35048 40740 35104 40796
rect 35152 40740 35208 40796
rect 4008 39956 4064 40012
rect 4112 39956 4168 40012
rect 4216 39956 4272 40012
rect 4320 39956 4376 40012
rect 4424 39956 4480 40012
rect 4528 39956 4584 40012
rect 4632 39956 4688 40012
rect 4736 39956 4792 40012
rect 4840 39956 4896 40012
rect 4944 39956 5000 40012
rect 5048 39956 5104 40012
rect 5152 39956 5208 40012
rect 24008 39956 24064 40012
rect 24112 39956 24168 40012
rect 24216 39956 24272 40012
rect 24320 39956 24376 40012
rect 24424 39956 24480 40012
rect 24528 39956 24584 40012
rect 24632 39956 24688 40012
rect 24736 39956 24792 40012
rect 24840 39956 24896 40012
rect 24944 39956 25000 40012
rect 25048 39956 25104 40012
rect 25152 39956 25208 40012
rect 14008 39172 14064 39228
rect 14112 39172 14168 39228
rect 14216 39172 14272 39228
rect 14320 39172 14376 39228
rect 14424 39172 14480 39228
rect 14528 39172 14584 39228
rect 14632 39172 14688 39228
rect 14736 39172 14792 39228
rect 14840 39172 14896 39228
rect 14944 39172 15000 39228
rect 15048 39172 15104 39228
rect 15152 39172 15208 39228
rect 34008 39172 34064 39228
rect 34112 39172 34168 39228
rect 34216 39172 34272 39228
rect 34320 39172 34376 39228
rect 34424 39172 34480 39228
rect 34528 39172 34584 39228
rect 34632 39172 34688 39228
rect 34736 39172 34792 39228
rect 34840 39172 34896 39228
rect 34944 39172 35000 39228
rect 35048 39172 35104 39228
rect 35152 39172 35208 39228
rect 4008 38388 4064 38444
rect 4112 38388 4168 38444
rect 4216 38388 4272 38444
rect 4320 38388 4376 38444
rect 4424 38388 4480 38444
rect 4528 38388 4584 38444
rect 4632 38388 4688 38444
rect 4736 38388 4792 38444
rect 4840 38388 4896 38444
rect 4944 38388 5000 38444
rect 5048 38388 5104 38444
rect 5152 38388 5208 38444
rect 24008 38388 24064 38444
rect 24112 38388 24168 38444
rect 24216 38388 24272 38444
rect 24320 38388 24376 38444
rect 24424 38388 24480 38444
rect 24528 38388 24584 38444
rect 24632 38388 24688 38444
rect 24736 38388 24792 38444
rect 24840 38388 24896 38444
rect 24944 38388 25000 38444
rect 25048 38388 25104 38444
rect 25152 38388 25208 38444
rect 14008 37604 14064 37660
rect 14112 37604 14168 37660
rect 14216 37604 14272 37660
rect 14320 37604 14376 37660
rect 14424 37604 14480 37660
rect 14528 37604 14584 37660
rect 14632 37604 14688 37660
rect 14736 37604 14792 37660
rect 14840 37604 14896 37660
rect 14944 37604 15000 37660
rect 15048 37604 15104 37660
rect 15152 37604 15208 37660
rect 34008 37604 34064 37660
rect 34112 37604 34168 37660
rect 34216 37604 34272 37660
rect 34320 37604 34376 37660
rect 34424 37604 34480 37660
rect 34528 37604 34584 37660
rect 34632 37604 34688 37660
rect 34736 37604 34792 37660
rect 34840 37604 34896 37660
rect 34944 37604 35000 37660
rect 35048 37604 35104 37660
rect 35152 37604 35208 37660
rect 4008 36820 4064 36876
rect 4112 36820 4168 36876
rect 4216 36820 4272 36876
rect 4320 36820 4376 36876
rect 4424 36820 4480 36876
rect 4528 36820 4584 36876
rect 4632 36820 4688 36876
rect 4736 36820 4792 36876
rect 4840 36820 4896 36876
rect 4944 36820 5000 36876
rect 5048 36820 5104 36876
rect 5152 36820 5208 36876
rect 24008 36820 24064 36876
rect 24112 36820 24168 36876
rect 24216 36820 24272 36876
rect 24320 36820 24376 36876
rect 24424 36820 24480 36876
rect 24528 36820 24584 36876
rect 24632 36820 24688 36876
rect 24736 36820 24792 36876
rect 24840 36820 24896 36876
rect 24944 36820 25000 36876
rect 25048 36820 25104 36876
rect 25152 36820 25208 36876
rect 14008 36036 14064 36092
rect 14112 36036 14168 36092
rect 14216 36036 14272 36092
rect 14320 36036 14376 36092
rect 14424 36036 14480 36092
rect 14528 36036 14584 36092
rect 14632 36036 14688 36092
rect 14736 36036 14792 36092
rect 14840 36036 14896 36092
rect 14944 36036 15000 36092
rect 15048 36036 15104 36092
rect 15152 36036 15208 36092
rect 34008 36036 34064 36092
rect 34112 36036 34168 36092
rect 34216 36036 34272 36092
rect 34320 36036 34376 36092
rect 34424 36036 34480 36092
rect 34528 36036 34584 36092
rect 34632 36036 34688 36092
rect 34736 36036 34792 36092
rect 34840 36036 34896 36092
rect 34944 36036 35000 36092
rect 35048 36036 35104 36092
rect 35152 36036 35208 36092
rect 4008 35252 4064 35308
rect 4112 35252 4168 35308
rect 4216 35252 4272 35308
rect 4320 35252 4376 35308
rect 4424 35252 4480 35308
rect 4528 35252 4584 35308
rect 4632 35252 4688 35308
rect 4736 35252 4792 35308
rect 4840 35252 4896 35308
rect 4944 35252 5000 35308
rect 5048 35252 5104 35308
rect 5152 35252 5208 35308
rect 24008 35252 24064 35308
rect 24112 35252 24168 35308
rect 24216 35252 24272 35308
rect 24320 35252 24376 35308
rect 24424 35252 24480 35308
rect 24528 35252 24584 35308
rect 24632 35252 24688 35308
rect 24736 35252 24792 35308
rect 24840 35252 24896 35308
rect 24944 35252 25000 35308
rect 25048 35252 25104 35308
rect 25152 35252 25208 35308
rect 14008 34468 14064 34524
rect 14112 34468 14168 34524
rect 14216 34468 14272 34524
rect 14320 34468 14376 34524
rect 14424 34468 14480 34524
rect 14528 34468 14584 34524
rect 14632 34468 14688 34524
rect 14736 34468 14792 34524
rect 14840 34468 14896 34524
rect 14944 34468 15000 34524
rect 15048 34468 15104 34524
rect 15152 34468 15208 34524
rect 34008 34468 34064 34524
rect 34112 34468 34168 34524
rect 34216 34468 34272 34524
rect 34320 34468 34376 34524
rect 34424 34468 34480 34524
rect 34528 34468 34584 34524
rect 34632 34468 34688 34524
rect 34736 34468 34792 34524
rect 34840 34468 34896 34524
rect 34944 34468 35000 34524
rect 35048 34468 35104 34524
rect 35152 34468 35208 34524
rect 4008 33684 4064 33740
rect 4112 33684 4168 33740
rect 4216 33684 4272 33740
rect 4320 33684 4376 33740
rect 4424 33684 4480 33740
rect 4528 33684 4584 33740
rect 4632 33684 4688 33740
rect 4736 33684 4792 33740
rect 4840 33684 4896 33740
rect 4944 33684 5000 33740
rect 5048 33684 5104 33740
rect 5152 33684 5208 33740
rect 24008 33684 24064 33740
rect 24112 33684 24168 33740
rect 24216 33684 24272 33740
rect 24320 33684 24376 33740
rect 24424 33684 24480 33740
rect 24528 33684 24584 33740
rect 24632 33684 24688 33740
rect 24736 33684 24792 33740
rect 24840 33684 24896 33740
rect 24944 33684 25000 33740
rect 25048 33684 25104 33740
rect 25152 33684 25208 33740
rect 14008 32900 14064 32956
rect 14112 32900 14168 32956
rect 14216 32900 14272 32956
rect 14320 32900 14376 32956
rect 14424 32900 14480 32956
rect 14528 32900 14584 32956
rect 14632 32900 14688 32956
rect 14736 32900 14792 32956
rect 14840 32900 14896 32956
rect 14944 32900 15000 32956
rect 15048 32900 15104 32956
rect 15152 32900 15208 32956
rect 34008 32900 34064 32956
rect 34112 32900 34168 32956
rect 34216 32900 34272 32956
rect 34320 32900 34376 32956
rect 34424 32900 34480 32956
rect 34528 32900 34584 32956
rect 34632 32900 34688 32956
rect 34736 32900 34792 32956
rect 34840 32900 34896 32956
rect 34944 32900 35000 32956
rect 35048 32900 35104 32956
rect 35152 32900 35208 32956
rect 4008 32116 4064 32172
rect 4112 32116 4168 32172
rect 4216 32116 4272 32172
rect 4320 32116 4376 32172
rect 4424 32116 4480 32172
rect 4528 32116 4584 32172
rect 4632 32116 4688 32172
rect 4736 32116 4792 32172
rect 4840 32116 4896 32172
rect 4944 32116 5000 32172
rect 5048 32116 5104 32172
rect 5152 32116 5208 32172
rect 24008 32116 24064 32172
rect 24112 32116 24168 32172
rect 24216 32116 24272 32172
rect 24320 32116 24376 32172
rect 24424 32116 24480 32172
rect 24528 32116 24584 32172
rect 24632 32116 24688 32172
rect 24736 32116 24792 32172
rect 24840 32116 24896 32172
rect 24944 32116 25000 32172
rect 25048 32116 25104 32172
rect 25152 32116 25208 32172
rect 14008 31332 14064 31388
rect 14112 31332 14168 31388
rect 14216 31332 14272 31388
rect 14320 31332 14376 31388
rect 14424 31332 14480 31388
rect 14528 31332 14584 31388
rect 14632 31332 14688 31388
rect 14736 31332 14792 31388
rect 14840 31332 14896 31388
rect 14944 31332 15000 31388
rect 15048 31332 15104 31388
rect 15152 31332 15208 31388
rect 34008 31332 34064 31388
rect 34112 31332 34168 31388
rect 34216 31332 34272 31388
rect 34320 31332 34376 31388
rect 34424 31332 34480 31388
rect 34528 31332 34584 31388
rect 34632 31332 34688 31388
rect 34736 31332 34792 31388
rect 34840 31332 34896 31388
rect 34944 31332 35000 31388
rect 35048 31332 35104 31388
rect 35152 31332 35208 31388
rect 4008 30548 4064 30604
rect 4112 30548 4168 30604
rect 4216 30548 4272 30604
rect 4320 30548 4376 30604
rect 4424 30548 4480 30604
rect 4528 30548 4584 30604
rect 4632 30548 4688 30604
rect 4736 30548 4792 30604
rect 4840 30548 4896 30604
rect 4944 30548 5000 30604
rect 5048 30548 5104 30604
rect 5152 30548 5208 30604
rect 24008 30548 24064 30604
rect 24112 30548 24168 30604
rect 24216 30548 24272 30604
rect 24320 30548 24376 30604
rect 24424 30548 24480 30604
rect 24528 30548 24584 30604
rect 24632 30548 24688 30604
rect 24736 30548 24792 30604
rect 24840 30548 24896 30604
rect 24944 30548 25000 30604
rect 25048 30548 25104 30604
rect 25152 30548 25208 30604
rect 14008 29764 14064 29820
rect 14112 29764 14168 29820
rect 14216 29764 14272 29820
rect 14320 29764 14376 29820
rect 14424 29764 14480 29820
rect 14528 29764 14584 29820
rect 14632 29764 14688 29820
rect 14736 29764 14792 29820
rect 14840 29764 14896 29820
rect 14944 29764 15000 29820
rect 15048 29764 15104 29820
rect 15152 29764 15208 29820
rect 34008 29764 34064 29820
rect 34112 29764 34168 29820
rect 34216 29764 34272 29820
rect 34320 29764 34376 29820
rect 34424 29764 34480 29820
rect 34528 29764 34584 29820
rect 34632 29764 34688 29820
rect 34736 29764 34792 29820
rect 34840 29764 34896 29820
rect 34944 29764 35000 29820
rect 35048 29764 35104 29820
rect 35152 29764 35208 29820
rect 4008 28980 4064 29036
rect 4112 28980 4168 29036
rect 4216 28980 4272 29036
rect 4320 28980 4376 29036
rect 4424 28980 4480 29036
rect 4528 28980 4584 29036
rect 4632 28980 4688 29036
rect 4736 28980 4792 29036
rect 4840 28980 4896 29036
rect 4944 28980 5000 29036
rect 5048 28980 5104 29036
rect 5152 28980 5208 29036
rect 24008 28980 24064 29036
rect 24112 28980 24168 29036
rect 24216 28980 24272 29036
rect 24320 28980 24376 29036
rect 24424 28980 24480 29036
rect 24528 28980 24584 29036
rect 24632 28980 24688 29036
rect 24736 28980 24792 29036
rect 24840 28980 24896 29036
rect 24944 28980 25000 29036
rect 25048 28980 25104 29036
rect 25152 28980 25208 29036
rect 14008 28196 14064 28252
rect 14112 28196 14168 28252
rect 14216 28196 14272 28252
rect 14320 28196 14376 28252
rect 14424 28196 14480 28252
rect 14528 28196 14584 28252
rect 14632 28196 14688 28252
rect 14736 28196 14792 28252
rect 14840 28196 14896 28252
rect 14944 28196 15000 28252
rect 15048 28196 15104 28252
rect 15152 28196 15208 28252
rect 34008 28196 34064 28252
rect 34112 28196 34168 28252
rect 34216 28196 34272 28252
rect 34320 28196 34376 28252
rect 34424 28196 34480 28252
rect 34528 28196 34584 28252
rect 34632 28196 34688 28252
rect 34736 28196 34792 28252
rect 34840 28196 34896 28252
rect 34944 28196 35000 28252
rect 35048 28196 35104 28252
rect 35152 28196 35208 28252
rect 4008 27412 4064 27468
rect 4112 27412 4168 27468
rect 4216 27412 4272 27468
rect 4320 27412 4376 27468
rect 4424 27412 4480 27468
rect 4528 27412 4584 27468
rect 4632 27412 4688 27468
rect 4736 27412 4792 27468
rect 4840 27412 4896 27468
rect 4944 27412 5000 27468
rect 5048 27412 5104 27468
rect 5152 27412 5208 27468
rect 24008 27412 24064 27468
rect 24112 27412 24168 27468
rect 24216 27412 24272 27468
rect 24320 27412 24376 27468
rect 24424 27412 24480 27468
rect 24528 27412 24584 27468
rect 24632 27412 24688 27468
rect 24736 27412 24792 27468
rect 24840 27412 24896 27468
rect 24944 27412 25000 27468
rect 25048 27412 25104 27468
rect 25152 27412 25208 27468
rect 14008 26628 14064 26684
rect 14112 26628 14168 26684
rect 14216 26628 14272 26684
rect 14320 26628 14376 26684
rect 14424 26628 14480 26684
rect 14528 26628 14584 26684
rect 14632 26628 14688 26684
rect 14736 26628 14792 26684
rect 14840 26628 14896 26684
rect 14944 26628 15000 26684
rect 15048 26628 15104 26684
rect 15152 26628 15208 26684
rect 34008 26628 34064 26684
rect 34112 26628 34168 26684
rect 34216 26628 34272 26684
rect 34320 26628 34376 26684
rect 34424 26628 34480 26684
rect 34528 26628 34584 26684
rect 34632 26628 34688 26684
rect 34736 26628 34792 26684
rect 34840 26628 34896 26684
rect 34944 26628 35000 26684
rect 35048 26628 35104 26684
rect 35152 26628 35208 26684
rect 4008 25844 4064 25900
rect 4112 25844 4168 25900
rect 4216 25844 4272 25900
rect 4320 25844 4376 25900
rect 4424 25844 4480 25900
rect 4528 25844 4584 25900
rect 4632 25844 4688 25900
rect 4736 25844 4792 25900
rect 4840 25844 4896 25900
rect 4944 25844 5000 25900
rect 5048 25844 5104 25900
rect 5152 25844 5208 25900
rect 24008 25844 24064 25900
rect 24112 25844 24168 25900
rect 24216 25844 24272 25900
rect 24320 25844 24376 25900
rect 24424 25844 24480 25900
rect 24528 25844 24584 25900
rect 24632 25844 24688 25900
rect 24736 25844 24792 25900
rect 24840 25844 24896 25900
rect 24944 25844 25000 25900
rect 25048 25844 25104 25900
rect 25152 25844 25208 25900
rect 14008 25060 14064 25116
rect 14112 25060 14168 25116
rect 14216 25060 14272 25116
rect 14320 25060 14376 25116
rect 14424 25060 14480 25116
rect 14528 25060 14584 25116
rect 14632 25060 14688 25116
rect 14736 25060 14792 25116
rect 14840 25060 14896 25116
rect 14944 25060 15000 25116
rect 15048 25060 15104 25116
rect 15152 25060 15208 25116
rect 34008 25060 34064 25116
rect 34112 25060 34168 25116
rect 34216 25060 34272 25116
rect 34320 25060 34376 25116
rect 34424 25060 34480 25116
rect 34528 25060 34584 25116
rect 34632 25060 34688 25116
rect 34736 25060 34792 25116
rect 34840 25060 34896 25116
rect 34944 25060 35000 25116
rect 35048 25060 35104 25116
rect 35152 25060 35208 25116
rect 4008 24276 4064 24332
rect 4112 24276 4168 24332
rect 4216 24276 4272 24332
rect 4320 24276 4376 24332
rect 4424 24276 4480 24332
rect 4528 24276 4584 24332
rect 4632 24276 4688 24332
rect 4736 24276 4792 24332
rect 4840 24276 4896 24332
rect 4944 24276 5000 24332
rect 5048 24276 5104 24332
rect 5152 24276 5208 24332
rect 24008 24276 24064 24332
rect 24112 24276 24168 24332
rect 24216 24276 24272 24332
rect 24320 24276 24376 24332
rect 24424 24276 24480 24332
rect 24528 24276 24584 24332
rect 24632 24276 24688 24332
rect 24736 24276 24792 24332
rect 24840 24276 24896 24332
rect 24944 24276 25000 24332
rect 25048 24276 25104 24332
rect 25152 24276 25208 24332
rect 14008 23492 14064 23548
rect 14112 23492 14168 23548
rect 14216 23492 14272 23548
rect 14320 23492 14376 23548
rect 14424 23492 14480 23548
rect 14528 23492 14584 23548
rect 14632 23492 14688 23548
rect 14736 23492 14792 23548
rect 14840 23492 14896 23548
rect 14944 23492 15000 23548
rect 15048 23492 15104 23548
rect 15152 23492 15208 23548
rect 34008 23492 34064 23548
rect 34112 23492 34168 23548
rect 34216 23492 34272 23548
rect 34320 23492 34376 23548
rect 34424 23492 34480 23548
rect 34528 23492 34584 23548
rect 34632 23492 34688 23548
rect 34736 23492 34792 23548
rect 34840 23492 34896 23548
rect 34944 23492 35000 23548
rect 35048 23492 35104 23548
rect 35152 23492 35208 23548
rect 4008 22708 4064 22764
rect 4112 22708 4168 22764
rect 4216 22708 4272 22764
rect 4320 22708 4376 22764
rect 4424 22708 4480 22764
rect 4528 22708 4584 22764
rect 4632 22708 4688 22764
rect 4736 22708 4792 22764
rect 4840 22708 4896 22764
rect 4944 22708 5000 22764
rect 5048 22708 5104 22764
rect 5152 22708 5208 22764
rect 24008 22708 24064 22764
rect 24112 22708 24168 22764
rect 24216 22708 24272 22764
rect 24320 22708 24376 22764
rect 24424 22708 24480 22764
rect 24528 22708 24584 22764
rect 24632 22708 24688 22764
rect 24736 22708 24792 22764
rect 24840 22708 24896 22764
rect 24944 22708 25000 22764
rect 25048 22708 25104 22764
rect 25152 22708 25208 22764
rect 14008 21924 14064 21980
rect 14112 21924 14168 21980
rect 14216 21924 14272 21980
rect 14320 21924 14376 21980
rect 14424 21924 14480 21980
rect 14528 21924 14584 21980
rect 14632 21924 14688 21980
rect 14736 21924 14792 21980
rect 14840 21924 14896 21980
rect 14944 21924 15000 21980
rect 15048 21924 15104 21980
rect 15152 21924 15208 21980
rect 34008 21924 34064 21980
rect 34112 21924 34168 21980
rect 34216 21924 34272 21980
rect 34320 21924 34376 21980
rect 34424 21924 34480 21980
rect 34528 21924 34584 21980
rect 34632 21924 34688 21980
rect 34736 21924 34792 21980
rect 34840 21924 34896 21980
rect 34944 21924 35000 21980
rect 35048 21924 35104 21980
rect 35152 21924 35208 21980
rect 4008 21140 4064 21196
rect 4112 21140 4168 21196
rect 4216 21140 4272 21196
rect 4320 21140 4376 21196
rect 4424 21140 4480 21196
rect 4528 21140 4584 21196
rect 4632 21140 4688 21196
rect 4736 21140 4792 21196
rect 4840 21140 4896 21196
rect 4944 21140 5000 21196
rect 5048 21140 5104 21196
rect 5152 21140 5208 21196
rect 24008 21140 24064 21196
rect 24112 21140 24168 21196
rect 24216 21140 24272 21196
rect 24320 21140 24376 21196
rect 24424 21140 24480 21196
rect 24528 21140 24584 21196
rect 24632 21140 24688 21196
rect 24736 21140 24792 21196
rect 24840 21140 24896 21196
rect 24944 21140 25000 21196
rect 25048 21140 25104 21196
rect 25152 21140 25208 21196
rect 14008 20356 14064 20412
rect 14112 20356 14168 20412
rect 14216 20356 14272 20412
rect 14320 20356 14376 20412
rect 14424 20356 14480 20412
rect 14528 20356 14584 20412
rect 14632 20356 14688 20412
rect 14736 20356 14792 20412
rect 14840 20356 14896 20412
rect 14944 20356 15000 20412
rect 15048 20356 15104 20412
rect 15152 20356 15208 20412
rect 34008 20356 34064 20412
rect 34112 20356 34168 20412
rect 34216 20356 34272 20412
rect 34320 20356 34376 20412
rect 34424 20356 34480 20412
rect 34528 20356 34584 20412
rect 34632 20356 34688 20412
rect 34736 20356 34792 20412
rect 34840 20356 34896 20412
rect 34944 20356 35000 20412
rect 35048 20356 35104 20412
rect 35152 20356 35208 20412
rect 4008 19572 4064 19628
rect 4112 19572 4168 19628
rect 4216 19572 4272 19628
rect 4320 19572 4376 19628
rect 4424 19572 4480 19628
rect 4528 19572 4584 19628
rect 4632 19572 4688 19628
rect 4736 19572 4792 19628
rect 4840 19572 4896 19628
rect 4944 19572 5000 19628
rect 5048 19572 5104 19628
rect 5152 19572 5208 19628
rect 24008 19572 24064 19628
rect 24112 19572 24168 19628
rect 24216 19572 24272 19628
rect 24320 19572 24376 19628
rect 24424 19572 24480 19628
rect 24528 19572 24584 19628
rect 24632 19572 24688 19628
rect 24736 19572 24792 19628
rect 24840 19572 24896 19628
rect 24944 19572 25000 19628
rect 25048 19572 25104 19628
rect 25152 19572 25208 19628
rect 14008 18788 14064 18844
rect 14112 18788 14168 18844
rect 14216 18788 14272 18844
rect 14320 18788 14376 18844
rect 14424 18788 14480 18844
rect 14528 18788 14584 18844
rect 14632 18788 14688 18844
rect 14736 18788 14792 18844
rect 14840 18788 14896 18844
rect 14944 18788 15000 18844
rect 15048 18788 15104 18844
rect 15152 18788 15208 18844
rect 34008 18788 34064 18844
rect 34112 18788 34168 18844
rect 34216 18788 34272 18844
rect 34320 18788 34376 18844
rect 34424 18788 34480 18844
rect 34528 18788 34584 18844
rect 34632 18788 34688 18844
rect 34736 18788 34792 18844
rect 34840 18788 34896 18844
rect 34944 18788 35000 18844
rect 35048 18788 35104 18844
rect 35152 18788 35208 18844
rect 4008 18004 4064 18060
rect 4112 18004 4168 18060
rect 4216 18004 4272 18060
rect 4320 18004 4376 18060
rect 4424 18004 4480 18060
rect 4528 18004 4584 18060
rect 4632 18004 4688 18060
rect 4736 18004 4792 18060
rect 4840 18004 4896 18060
rect 4944 18004 5000 18060
rect 5048 18004 5104 18060
rect 5152 18004 5208 18060
rect 24008 18004 24064 18060
rect 24112 18004 24168 18060
rect 24216 18004 24272 18060
rect 24320 18004 24376 18060
rect 24424 18004 24480 18060
rect 24528 18004 24584 18060
rect 24632 18004 24688 18060
rect 24736 18004 24792 18060
rect 24840 18004 24896 18060
rect 24944 18004 25000 18060
rect 25048 18004 25104 18060
rect 25152 18004 25208 18060
rect 14008 17220 14064 17276
rect 14112 17220 14168 17276
rect 14216 17220 14272 17276
rect 14320 17220 14376 17276
rect 14424 17220 14480 17276
rect 14528 17220 14584 17276
rect 14632 17220 14688 17276
rect 14736 17220 14792 17276
rect 14840 17220 14896 17276
rect 14944 17220 15000 17276
rect 15048 17220 15104 17276
rect 15152 17220 15208 17276
rect 34008 17220 34064 17276
rect 34112 17220 34168 17276
rect 34216 17220 34272 17276
rect 34320 17220 34376 17276
rect 34424 17220 34480 17276
rect 34528 17220 34584 17276
rect 34632 17220 34688 17276
rect 34736 17220 34792 17276
rect 34840 17220 34896 17276
rect 34944 17220 35000 17276
rect 35048 17220 35104 17276
rect 35152 17220 35208 17276
rect 4008 16436 4064 16492
rect 4112 16436 4168 16492
rect 4216 16436 4272 16492
rect 4320 16436 4376 16492
rect 4424 16436 4480 16492
rect 4528 16436 4584 16492
rect 4632 16436 4688 16492
rect 4736 16436 4792 16492
rect 4840 16436 4896 16492
rect 4944 16436 5000 16492
rect 5048 16436 5104 16492
rect 5152 16436 5208 16492
rect 24008 16436 24064 16492
rect 24112 16436 24168 16492
rect 24216 16436 24272 16492
rect 24320 16436 24376 16492
rect 24424 16436 24480 16492
rect 24528 16436 24584 16492
rect 24632 16436 24688 16492
rect 24736 16436 24792 16492
rect 24840 16436 24896 16492
rect 24944 16436 25000 16492
rect 25048 16436 25104 16492
rect 25152 16436 25208 16492
rect 14008 15652 14064 15708
rect 14112 15652 14168 15708
rect 14216 15652 14272 15708
rect 14320 15652 14376 15708
rect 14424 15652 14480 15708
rect 14528 15652 14584 15708
rect 14632 15652 14688 15708
rect 14736 15652 14792 15708
rect 14840 15652 14896 15708
rect 14944 15652 15000 15708
rect 15048 15652 15104 15708
rect 15152 15652 15208 15708
rect 34008 15652 34064 15708
rect 34112 15652 34168 15708
rect 34216 15652 34272 15708
rect 34320 15652 34376 15708
rect 34424 15652 34480 15708
rect 34528 15652 34584 15708
rect 34632 15652 34688 15708
rect 34736 15652 34792 15708
rect 34840 15652 34896 15708
rect 34944 15652 35000 15708
rect 35048 15652 35104 15708
rect 35152 15652 35208 15708
rect 4008 14868 4064 14924
rect 4112 14868 4168 14924
rect 4216 14868 4272 14924
rect 4320 14868 4376 14924
rect 4424 14868 4480 14924
rect 4528 14868 4584 14924
rect 4632 14868 4688 14924
rect 4736 14868 4792 14924
rect 4840 14868 4896 14924
rect 4944 14868 5000 14924
rect 5048 14868 5104 14924
rect 5152 14868 5208 14924
rect 24008 14868 24064 14924
rect 24112 14868 24168 14924
rect 24216 14868 24272 14924
rect 24320 14868 24376 14924
rect 24424 14868 24480 14924
rect 24528 14868 24584 14924
rect 24632 14868 24688 14924
rect 24736 14868 24792 14924
rect 24840 14868 24896 14924
rect 24944 14868 25000 14924
rect 25048 14868 25104 14924
rect 25152 14868 25208 14924
rect 14008 14084 14064 14140
rect 14112 14084 14168 14140
rect 14216 14084 14272 14140
rect 14320 14084 14376 14140
rect 14424 14084 14480 14140
rect 14528 14084 14584 14140
rect 14632 14084 14688 14140
rect 14736 14084 14792 14140
rect 14840 14084 14896 14140
rect 14944 14084 15000 14140
rect 15048 14084 15104 14140
rect 15152 14084 15208 14140
rect 34008 14084 34064 14140
rect 34112 14084 34168 14140
rect 34216 14084 34272 14140
rect 34320 14084 34376 14140
rect 34424 14084 34480 14140
rect 34528 14084 34584 14140
rect 34632 14084 34688 14140
rect 34736 14084 34792 14140
rect 34840 14084 34896 14140
rect 34944 14084 35000 14140
rect 35048 14084 35104 14140
rect 35152 14084 35208 14140
rect 4008 13300 4064 13356
rect 4112 13300 4168 13356
rect 4216 13300 4272 13356
rect 4320 13300 4376 13356
rect 4424 13300 4480 13356
rect 4528 13300 4584 13356
rect 4632 13300 4688 13356
rect 4736 13300 4792 13356
rect 4840 13300 4896 13356
rect 4944 13300 5000 13356
rect 5048 13300 5104 13356
rect 5152 13300 5208 13356
rect 24008 13300 24064 13356
rect 24112 13300 24168 13356
rect 24216 13300 24272 13356
rect 24320 13300 24376 13356
rect 24424 13300 24480 13356
rect 24528 13300 24584 13356
rect 24632 13300 24688 13356
rect 24736 13300 24792 13356
rect 24840 13300 24896 13356
rect 24944 13300 25000 13356
rect 25048 13300 25104 13356
rect 25152 13300 25208 13356
rect 14008 12516 14064 12572
rect 14112 12516 14168 12572
rect 14216 12516 14272 12572
rect 14320 12516 14376 12572
rect 14424 12516 14480 12572
rect 14528 12516 14584 12572
rect 14632 12516 14688 12572
rect 14736 12516 14792 12572
rect 14840 12516 14896 12572
rect 14944 12516 15000 12572
rect 15048 12516 15104 12572
rect 15152 12516 15208 12572
rect 34008 12516 34064 12572
rect 34112 12516 34168 12572
rect 34216 12516 34272 12572
rect 34320 12516 34376 12572
rect 34424 12516 34480 12572
rect 34528 12516 34584 12572
rect 34632 12516 34688 12572
rect 34736 12516 34792 12572
rect 34840 12516 34896 12572
rect 34944 12516 35000 12572
rect 35048 12516 35104 12572
rect 35152 12516 35208 12572
rect 4008 11732 4064 11788
rect 4112 11732 4168 11788
rect 4216 11732 4272 11788
rect 4320 11732 4376 11788
rect 4424 11732 4480 11788
rect 4528 11732 4584 11788
rect 4632 11732 4688 11788
rect 4736 11732 4792 11788
rect 4840 11732 4896 11788
rect 4944 11732 5000 11788
rect 5048 11732 5104 11788
rect 5152 11732 5208 11788
rect 24008 11732 24064 11788
rect 24112 11732 24168 11788
rect 24216 11732 24272 11788
rect 24320 11732 24376 11788
rect 24424 11732 24480 11788
rect 24528 11732 24584 11788
rect 24632 11732 24688 11788
rect 24736 11732 24792 11788
rect 24840 11732 24896 11788
rect 24944 11732 25000 11788
rect 25048 11732 25104 11788
rect 25152 11732 25208 11788
rect 14008 10948 14064 11004
rect 14112 10948 14168 11004
rect 14216 10948 14272 11004
rect 14320 10948 14376 11004
rect 14424 10948 14480 11004
rect 14528 10948 14584 11004
rect 14632 10948 14688 11004
rect 14736 10948 14792 11004
rect 14840 10948 14896 11004
rect 14944 10948 15000 11004
rect 15048 10948 15104 11004
rect 15152 10948 15208 11004
rect 34008 10948 34064 11004
rect 34112 10948 34168 11004
rect 34216 10948 34272 11004
rect 34320 10948 34376 11004
rect 34424 10948 34480 11004
rect 34528 10948 34584 11004
rect 34632 10948 34688 11004
rect 34736 10948 34792 11004
rect 34840 10948 34896 11004
rect 34944 10948 35000 11004
rect 35048 10948 35104 11004
rect 35152 10948 35208 11004
rect 4008 10164 4064 10220
rect 4112 10164 4168 10220
rect 4216 10164 4272 10220
rect 4320 10164 4376 10220
rect 4424 10164 4480 10220
rect 4528 10164 4584 10220
rect 4632 10164 4688 10220
rect 4736 10164 4792 10220
rect 4840 10164 4896 10220
rect 4944 10164 5000 10220
rect 5048 10164 5104 10220
rect 5152 10164 5208 10220
rect 24008 10164 24064 10220
rect 24112 10164 24168 10220
rect 24216 10164 24272 10220
rect 24320 10164 24376 10220
rect 24424 10164 24480 10220
rect 24528 10164 24584 10220
rect 24632 10164 24688 10220
rect 24736 10164 24792 10220
rect 24840 10164 24896 10220
rect 24944 10164 25000 10220
rect 25048 10164 25104 10220
rect 25152 10164 25208 10220
rect 14008 9380 14064 9436
rect 14112 9380 14168 9436
rect 14216 9380 14272 9436
rect 14320 9380 14376 9436
rect 14424 9380 14480 9436
rect 14528 9380 14584 9436
rect 14632 9380 14688 9436
rect 14736 9380 14792 9436
rect 14840 9380 14896 9436
rect 14944 9380 15000 9436
rect 15048 9380 15104 9436
rect 15152 9380 15208 9436
rect 34008 9380 34064 9436
rect 34112 9380 34168 9436
rect 34216 9380 34272 9436
rect 34320 9380 34376 9436
rect 34424 9380 34480 9436
rect 34528 9380 34584 9436
rect 34632 9380 34688 9436
rect 34736 9380 34792 9436
rect 34840 9380 34896 9436
rect 34944 9380 35000 9436
rect 35048 9380 35104 9436
rect 35152 9380 35208 9436
rect 7420 8652 7476 8708
rect 4008 8596 4064 8652
rect 4112 8596 4168 8652
rect 4216 8596 4272 8652
rect 4320 8596 4376 8652
rect 4424 8596 4480 8652
rect 4528 8596 4584 8652
rect 4632 8596 4688 8652
rect 4736 8596 4792 8652
rect 4840 8596 4896 8652
rect 4944 8596 5000 8652
rect 5048 8596 5104 8652
rect 5152 8596 5208 8652
rect 24008 8596 24064 8652
rect 24112 8596 24168 8652
rect 24216 8596 24272 8652
rect 24320 8596 24376 8652
rect 24424 8596 24480 8652
rect 24528 8596 24584 8652
rect 24632 8596 24688 8652
rect 24736 8596 24792 8652
rect 24840 8596 24896 8652
rect 24944 8596 25000 8652
rect 25048 8596 25104 8652
rect 25152 8596 25208 8652
rect 5628 8204 5684 8260
rect 6524 7980 6580 8036
rect 6972 7980 7028 8036
rect 14008 7812 14064 7868
rect 14112 7812 14168 7868
rect 14216 7812 14272 7868
rect 14320 7812 14376 7868
rect 14424 7812 14480 7868
rect 14528 7812 14584 7868
rect 14632 7812 14688 7868
rect 14736 7812 14792 7868
rect 14840 7812 14896 7868
rect 14944 7812 15000 7868
rect 15048 7812 15104 7868
rect 15152 7812 15208 7868
rect 34008 7812 34064 7868
rect 34112 7812 34168 7868
rect 34216 7812 34272 7868
rect 34320 7812 34376 7868
rect 34424 7812 34480 7868
rect 34528 7812 34584 7868
rect 34632 7812 34688 7868
rect 34736 7812 34792 7868
rect 34840 7812 34896 7868
rect 34944 7812 35000 7868
rect 35048 7812 35104 7868
rect 35152 7812 35208 7868
rect 7084 7420 7140 7476
rect 5740 7084 5796 7140
rect 4008 7028 4064 7084
rect 4112 7028 4168 7084
rect 4216 7028 4272 7084
rect 4320 7028 4376 7084
rect 4424 7028 4480 7084
rect 4528 7028 4584 7084
rect 4632 7028 4688 7084
rect 4736 7028 4792 7084
rect 4840 7028 4896 7084
rect 4944 7028 5000 7084
rect 5048 7028 5104 7084
rect 5152 7028 5208 7084
rect 24008 7028 24064 7084
rect 24112 7028 24168 7084
rect 24216 7028 24272 7084
rect 24320 7028 24376 7084
rect 24424 7028 24480 7084
rect 24528 7028 24584 7084
rect 24632 7028 24688 7084
rect 24736 7028 24792 7084
rect 24840 7028 24896 7084
rect 24944 7028 25000 7084
rect 25048 7028 25104 7084
rect 25152 7028 25208 7084
rect 7420 6860 7476 6916
rect 7980 6636 8036 6692
rect 7420 6300 7476 6356
rect 14008 6244 14064 6300
rect 14112 6244 14168 6300
rect 14216 6244 14272 6300
rect 14320 6244 14376 6300
rect 14424 6244 14480 6300
rect 14528 6244 14584 6300
rect 14632 6244 14688 6300
rect 14736 6244 14792 6300
rect 14840 6244 14896 6300
rect 14944 6244 15000 6300
rect 15048 6244 15104 6300
rect 15152 6244 15208 6300
rect 34008 6244 34064 6300
rect 34112 6244 34168 6300
rect 34216 6244 34272 6300
rect 34320 6244 34376 6300
rect 34424 6244 34480 6300
rect 34528 6244 34584 6300
rect 34632 6244 34688 6300
rect 34736 6244 34792 6300
rect 34840 6244 34896 6300
rect 34944 6244 35000 6300
rect 35048 6244 35104 6300
rect 35152 6244 35208 6300
rect 6188 6188 6244 6244
rect 7084 6188 7140 6244
rect 7980 6188 8036 6244
rect 5740 5964 5796 6020
rect 5628 5628 5684 5684
rect 4008 5460 4064 5516
rect 4112 5460 4168 5516
rect 4216 5460 4272 5516
rect 4320 5460 4376 5516
rect 4424 5460 4480 5516
rect 4528 5460 4584 5516
rect 4632 5460 4688 5516
rect 4736 5460 4792 5516
rect 4840 5460 4896 5516
rect 4944 5460 5000 5516
rect 5048 5460 5104 5516
rect 5152 5460 5208 5516
rect 24008 5460 24064 5516
rect 24112 5460 24168 5516
rect 24216 5460 24272 5516
rect 24320 5460 24376 5516
rect 24424 5460 24480 5516
rect 24528 5460 24584 5516
rect 24632 5460 24688 5516
rect 24736 5460 24792 5516
rect 24840 5460 24896 5516
rect 24944 5460 25000 5516
rect 25048 5460 25104 5516
rect 25152 5460 25208 5516
rect 5628 4956 5684 5012
rect 6188 4844 6244 4900
rect 15708 4732 15764 4788
rect 14008 4676 14064 4732
rect 14112 4676 14168 4732
rect 14216 4676 14272 4732
rect 14320 4676 14376 4732
rect 14424 4676 14480 4732
rect 14528 4676 14584 4732
rect 14632 4676 14688 4732
rect 14736 4676 14792 4732
rect 14840 4676 14896 4732
rect 14944 4676 15000 4732
rect 15048 4676 15104 4732
rect 15152 4676 15208 4732
rect 34008 4676 34064 4732
rect 34112 4676 34168 4732
rect 34216 4676 34272 4732
rect 34320 4676 34376 4732
rect 34424 4676 34480 4732
rect 34528 4676 34584 4732
rect 34632 4676 34688 4732
rect 34736 4676 34792 4732
rect 34840 4676 34896 4732
rect 34944 4676 35000 4732
rect 35048 4676 35104 4732
rect 35152 4676 35208 4732
rect 15708 3948 15764 4004
rect 4008 3892 4064 3948
rect 4112 3892 4168 3948
rect 4216 3892 4272 3948
rect 4320 3892 4376 3948
rect 4424 3892 4480 3948
rect 4528 3892 4584 3948
rect 4632 3892 4688 3948
rect 4736 3892 4792 3948
rect 4840 3892 4896 3948
rect 4944 3892 5000 3948
rect 5048 3892 5104 3948
rect 5152 3892 5208 3948
rect 24008 3892 24064 3948
rect 24112 3892 24168 3948
rect 24216 3892 24272 3948
rect 24320 3892 24376 3948
rect 24424 3892 24480 3948
rect 24528 3892 24584 3948
rect 24632 3892 24688 3948
rect 24736 3892 24792 3948
rect 24840 3892 24896 3948
rect 24944 3892 25000 3948
rect 25048 3892 25104 3948
rect 25152 3892 25208 3948
rect 6524 3724 6580 3780
rect 6972 3276 7028 3332
rect 14008 3108 14064 3164
rect 14112 3108 14168 3164
rect 14216 3108 14272 3164
rect 14320 3108 14376 3164
rect 14424 3108 14480 3164
rect 14528 3108 14584 3164
rect 14632 3108 14688 3164
rect 14736 3108 14792 3164
rect 14840 3108 14896 3164
rect 14944 3108 15000 3164
rect 15048 3108 15104 3164
rect 15152 3108 15208 3164
rect 34008 3108 34064 3164
rect 34112 3108 34168 3164
rect 34216 3108 34272 3164
rect 34320 3108 34376 3164
rect 34424 3108 34480 3164
rect 34528 3108 34584 3164
rect 34632 3108 34688 3164
rect 34736 3108 34792 3164
rect 34840 3108 34896 3164
rect 34944 3108 35000 3164
rect 35048 3108 35104 3164
rect 35152 3108 35208 3164
<< metal4 >>
rect 3988 46284 5228 46316
rect 3988 46228 4008 46284
rect 4064 46228 4112 46284
rect 4168 46228 4216 46284
rect 4272 46228 4320 46284
rect 4376 46228 4424 46284
rect 4480 46228 4528 46284
rect 4584 46228 4632 46284
rect 4688 46228 4736 46284
rect 4792 46228 4840 46284
rect 4896 46228 4944 46284
rect 5000 46228 5048 46284
rect 5104 46228 5152 46284
rect 5208 46228 5228 46284
rect 3988 44716 5228 46228
rect 3988 44660 4008 44716
rect 4064 44660 4112 44716
rect 4168 44660 4216 44716
rect 4272 44660 4320 44716
rect 4376 44660 4424 44716
rect 4480 44660 4528 44716
rect 4584 44660 4632 44716
rect 4688 44660 4736 44716
rect 4792 44660 4840 44716
rect 4896 44660 4944 44716
rect 5000 44660 5048 44716
rect 5104 44660 5152 44716
rect 5208 44660 5228 44716
rect 3988 43148 5228 44660
rect 3988 43092 4008 43148
rect 4064 43092 4112 43148
rect 4168 43092 4216 43148
rect 4272 43092 4320 43148
rect 4376 43092 4424 43148
rect 4480 43092 4528 43148
rect 4584 43092 4632 43148
rect 4688 43092 4736 43148
rect 4792 43092 4840 43148
rect 4896 43092 4944 43148
rect 5000 43092 5048 43148
rect 5104 43092 5152 43148
rect 5208 43092 5228 43148
rect 3988 41580 5228 43092
rect 3988 41524 4008 41580
rect 4064 41524 4112 41580
rect 4168 41524 4216 41580
rect 4272 41524 4320 41580
rect 4376 41524 4424 41580
rect 4480 41524 4528 41580
rect 4584 41524 4632 41580
rect 4688 41524 4736 41580
rect 4792 41524 4840 41580
rect 4896 41524 4944 41580
rect 5000 41524 5048 41580
rect 5104 41524 5152 41580
rect 5208 41524 5228 41580
rect 3988 40012 5228 41524
rect 3988 39956 4008 40012
rect 4064 39956 4112 40012
rect 4168 39956 4216 40012
rect 4272 39956 4320 40012
rect 4376 39956 4424 40012
rect 4480 39956 4528 40012
rect 4584 39956 4632 40012
rect 4688 39956 4736 40012
rect 4792 39956 4840 40012
rect 4896 39956 4944 40012
rect 5000 39956 5048 40012
rect 5104 39956 5152 40012
rect 5208 39956 5228 40012
rect 3988 38444 5228 39956
rect 3988 38388 4008 38444
rect 4064 38388 4112 38444
rect 4168 38388 4216 38444
rect 4272 38388 4320 38444
rect 4376 38388 4424 38444
rect 4480 38388 4528 38444
rect 4584 38388 4632 38444
rect 4688 38388 4736 38444
rect 4792 38388 4840 38444
rect 4896 38388 4944 38444
rect 5000 38388 5048 38444
rect 5104 38388 5152 38444
rect 5208 38388 5228 38444
rect 3988 36876 5228 38388
rect 3988 36820 4008 36876
rect 4064 36820 4112 36876
rect 4168 36820 4216 36876
rect 4272 36820 4320 36876
rect 4376 36820 4424 36876
rect 4480 36820 4528 36876
rect 4584 36820 4632 36876
rect 4688 36820 4736 36876
rect 4792 36820 4840 36876
rect 4896 36820 4944 36876
rect 5000 36820 5048 36876
rect 5104 36820 5152 36876
rect 5208 36820 5228 36876
rect 3988 35308 5228 36820
rect 3988 35252 4008 35308
rect 4064 35252 4112 35308
rect 4168 35252 4216 35308
rect 4272 35252 4320 35308
rect 4376 35252 4424 35308
rect 4480 35252 4528 35308
rect 4584 35252 4632 35308
rect 4688 35252 4736 35308
rect 4792 35252 4840 35308
rect 4896 35252 4944 35308
rect 5000 35252 5048 35308
rect 5104 35252 5152 35308
rect 5208 35252 5228 35308
rect 3988 33740 5228 35252
rect 3988 33684 4008 33740
rect 4064 33684 4112 33740
rect 4168 33684 4216 33740
rect 4272 33684 4320 33740
rect 4376 33684 4424 33740
rect 4480 33684 4528 33740
rect 4584 33684 4632 33740
rect 4688 33684 4736 33740
rect 4792 33684 4840 33740
rect 4896 33684 4944 33740
rect 5000 33684 5048 33740
rect 5104 33684 5152 33740
rect 5208 33684 5228 33740
rect 3988 32172 5228 33684
rect 3988 32116 4008 32172
rect 4064 32116 4112 32172
rect 4168 32116 4216 32172
rect 4272 32116 4320 32172
rect 4376 32116 4424 32172
rect 4480 32116 4528 32172
rect 4584 32116 4632 32172
rect 4688 32116 4736 32172
rect 4792 32116 4840 32172
rect 4896 32116 4944 32172
rect 5000 32116 5048 32172
rect 5104 32116 5152 32172
rect 5208 32116 5228 32172
rect 3988 30604 5228 32116
rect 3988 30548 4008 30604
rect 4064 30548 4112 30604
rect 4168 30548 4216 30604
rect 4272 30548 4320 30604
rect 4376 30548 4424 30604
rect 4480 30548 4528 30604
rect 4584 30548 4632 30604
rect 4688 30548 4736 30604
rect 4792 30548 4840 30604
rect 4896 30548 4944 30604
rect 5000 30548 5048 30604
rect 5104 30548 5152 30604
rect 5208 30548 5228 30604
rect 3988 29036 5228 30548
rect 3988 28980 4008 29036
rect 4064 28980 4112 29036
rect 4168 28980 4216 29036
rect 4272 28980 4320 29036
rect 4376 28980 4424 29036
rect 4480 28980 4528 29036
rect 4584 28980 4632 29036
rect 4688 28980 4736 29036
rect 4792 28980 4840 29036
rect 4896 28980 4944 29036
rect 5000 28980 5048 29036
rect 5104 28980 5152 29036
rect 5208 28980 5228 29036
rect 3988 27468 5228 28980
rect 3988 27412 4008 27468
rect 4064 27412 4112 27468
rect 4168 27412 4216 27468
rect 4272 27412 4320 27468
rect 4376 27412 4424 27468
rect 4480 27412 4528 27468
rect 4584 27412 4632 27468
rect 4688 27412 4736 27468
rect 4792 27412 4840 27468
rect 4896 27412 4944 27468
rect 5000 27412 5048 27468
rect 5104 27412 5152 27468
rect 5208 27412 5228 27468
rect 3988 25900 5228 27412
rect 3988 25844 4008 25900
rect 4064 25844 4112 25900
rect 4168 25844 4216 25900
rect 4272 25844 4320 25900
rect 4376 25844 4424 25900
rect 4480 25844 4528 25900
rect 4584 25844 4632 25900
rect 4688 25844 4736 25900
rect 4792 25844 4840 25900
rect 4896 25844 4944 25900
rect 5000 25844 5048 25900
rect 5104 25844 5152 25900
rect 5208 25844 5228 25900
rect 3988 24332 5228 25844
rect 3988 24276 4008 24332
rect 4064 24276 4112 24332
rect 4168 24276 4216 24332
rect 4272 24276 4320 24332
rect 4376 24276 4424 24332
rect 4480 24276 4528 24332
rect 4584 24276 4632 24332
rect 4688 24276 4736 24332
rect 4792 24276 4840 24332
rect 4896 24276 4944 24332
rect 5000 24276 5048 24332
rect 5104 24276 5152 24332
rect 5208 24276 5228 24332
rect 3988 22764 5228 24276
rect 3988 22708 4008 22764
rect 4064 22708 4112 22764
rect 4168 22708 4216 22764
rect 4272 22708 4320 22764
rect 4376 22708 4424 22764
rect 4480 22708 4528 22764
rect 4584 22708 4632 22764
rect 4688 22708 4736 22764
rect 4792 22708 4840 22764
rect 4896 22708 4944 22764
rect 5000 22708 5048 22764
rect 5104 22708 5152 22764
rect 5208 22708 5228 22764
rect 3988 21196 5228 22708
rect 3988 21140 4008 21196
rect 4064 21140 4112 21196
rect 4168 21140 4216 21196
rect 4272 21140 4320 21196
rect 4376 21140 4424 21196
rect 4480 21140 4528 21196
rect 4584 21140 4632 21196
rect 4688 21140 4736 21196
rect 4792 21140 4840 21196
rect 4896 21140 4944 21196
rect 5000 21140 5048 21196
rect 5104 21140 5152 21196
rect 5208 21140 5228 21196
rect 3988 19628 5228 21140
rect 3988 19572 4008 19628
rect 4064 19572 4112 19628
rect 4168 19572 4216 19628
rect 4272 19572 4320 19628
rect 4376 19572 4424 19628
rect 4480 19572 4528 19628
rect 4584 19572 4632 19628
rect 4688 19572 4736 19628
rect 4792 19572 4840 19628
rect 4896 19572 4944 19628
rect 5000 19572 5048 19628
rect 5104 19572 5152 19628
rect 5208 19572 5228 19628
rect 3988 18060 5228 19572
rect 3988 18004 4008 18060
rect 4064 18004 4112 18060
rect 4168 18004 4216 18060
rect 4272 18004 4320 18060
rect 4376 18004 4424 18060
rect 4480 18004 4528 18060
rect 4584 18004 4632 18060
rect 4688 18004 4736 18060
rect 4792 18004 4840 18060
rect 4896 18004 4944 18060
rect 5000 18004 5048 18060
rect 5104 18004 5152 18060
rect 5208 18004 5228 18060
rect 3988 16492 5228 18004
rect 3988 16436 4008 16492
rect 4064 16436 4112 16492
rect 4168 16436 4216 16492
rect 4272 16436 4320 16492
rect 4376 16436 4424 16492
rect 4480 16436 4528 16492
rect 4584 16436 4632 16492
rect 4688 16436 4736 16492
rect 4792 16436 4840 16492
rect 4896 16436 4944 16492
rect 5000 16436 5048 16492
rect 5104 16436 5152 16492
rect 5208 16436 5228 16492
rect 3988 14924 5228 16436
rect 3988 14868 4008 14924
rect 4064 14868 4112 14924
rect 4168 14868 4216 14924
rect 4272 14868 4320 14924
rect 4376 14868 4424 14924
rect 4480 14868 4528 14924
rect 4584 14868 4632 14924
rect 4688 14868 4736 14924
rect 4792 14868 4840 14924
rect 4896 14868 4944 14924
rect 5000 14868 5048 14924
rect 5104 14868 5152 14924
rect 5208 14868 5228 14924
rect 3988 13356 5228 14868
rect 3988 13300 4008 13356
rect 4064 13300 4112 13356
rect 4168 13300 4216 13356
rect 4272 13300 4320 13356
rect 4376 13300 4424 13356
rect 4480 13300 4528 13356
rect 4584 13300 4632 13356
rect 4688 13300 4736 13356
rect 4792 13300 4840 13356
rect 4896 13300 4944 13356
rect 5000 13300 5048 13356
rect 5104 13300 5152 13356
rect 5208 13300 5228 13356
rect 3988 11788 5228 13300
rect 3988 11732 4008 11788
rect 4064 11732 4112 11788
rect 4168 11732 4216 11788
rect 4272 11732 4320 11788
rect 4376 11732 4424 11788
rect 4480 11732 4528 11788
rect 4584 11732 4632 11788
rect 4688 11732 4736 11788
rect 4792 11732 4840 11788
rect 4896 11732 4944 11788
rect 5000 11732 5048 11788
rect 5104 11732 5152 11788
rect 5208 11732 5228 11788
rect 3988 10220 5228 11732
rect 3988 10164 4008 10220
rect 4064 10164 4112 10220
rect 4168 10164 4216 10220
rect 4272 10164 4320 10220
rect 4376 10164 4424 10220
rect 4480 10164 4528 10220
rect 4584 10164 4632 10220
rect 4688 10164 4736 10220
rect 4792 10164 4840 10220
rect 4896 10164 4944 10220
rect 5000 10164 5048 10220
rect 5104 10164 5152 10220
rect 5208 10164 5228 10220
rect 3988 8652 5228 10164
rect 13988 45500 15228 46316
rect 13988 45444 14008 45500
rect 14064 45444 14112 45500
rect 14168 45444 14216 45500
rect 14272 45444 14320 45500
rect 14376 45444 14424 45500
rect 14480 45444 14528 45500
rect 14584 45444 14632 45500
rect 14688 45444 14736 45500
rect 14792 45444 14840 45500
rect 14896 45444 14944 45500
rect 15000 45444 15048 45500
rect 15104 45444 15152 45500
rect 15208 45444 15228 45500
rect 13988 43932 15228 45444
rect 13988 43876 14008 43932
rect 14064 43876 14112 43932
rect 14168 43876 14216 43932
rect 14272 43876 14320 43932
rect 14376 43876 14424 43932
rect 14480 43876 14528 43932
rect 14584 43876 14632 43932
rect 14688 43876 14736 43932
rect 14792 43876 14840 43932
rect 14896 43876 14944 43932
rect 15000 43876 15048 43932
rect 15104 43876 15152 43932
rect 15208 43876 15228 43932
rect 13988 42364 15228 43876
rect 13988 42308 14008 42364
rect 14064 42308 14112 42364
rect 14168 42308 14216 42364
rect 14272 42308 14320 42364
rect 14376 42308 14424 42364
rect 14480 42308 14528 42364
rect 14584 42308 14632 42364
rect 14688 42308 14736 42364
rect 14792 42308 14840 42364
rect 14896 42308 14944 42364
rect 15000 42308 15048 42364
rect 15104 42308 15152 42364
rect 15208 42308 15228 42364
rect 13988 40796 15228 42308
rect 13988 40740 14008 40796
rect 14064 40740 14112 40796
rect 14168 40740 14216 40796
rect 14272 40740 14320 40796
rect 14376 40740 14424 40796
rect 14480 40740 14528 40796
rect 14584 40740 14632 40796
rect 14688 40740 14736 40796
rect 14792 40740 14840 40796
rect 14896 40740 14944 40796
rect 15000 40740 15048 40796
rect 15104 40740 15152 40796
rect 15208 40740 15228 40796
rect 13988 39228 15228 40740
rect 13988 39172 14008 39228
rect 14064 39172 14112 39228
rect 14168 39172 14216 39228
rect 14272 39172 14320 39228
rect 14376 39172 14424 39228
rect 14480 39172 14528 39228
rect 14584 39172 14632 39228
rect 14688 39172 14736 39228
rect 14792 39172 14840 39228
rect 14896 39172 14944 39228
rect 15000 39172 15048 39228
rect 15104 39172 15152 39228
rect 15208 39172 15228 39228
rect 13988 37660 15228 39172
rect 13988 37604 14008 37660
rect 14064 37604 14112 37660
rect 14168 37604 14216 37660
rect 14272 37604 14320 37660
rect 14376 37604 14424 37660
rect 14480 37604 14528 37660
rect 14584 37604 14632 37660
rect 14688 37604 14736 37660
rect 14792 37604 14840 37660
rect 14896 37604 14944 37660
rect 15000 37604 15048 37660
rect 15104 37604 15152 37660
rect 15208 37604 15228 37660
rect 13988 36092 15228 37604
rect 13988 36036 14008 36092
rect 14064 36036 14112 36092
rect 14168 36036 14216 36092
rect 14272 36036 14320 36092
rect 14376 36036 14424 36092
rect 14480 36036 14528 36092
rect 14584 36036 14632 36092
rect 14688 36036 14736 36092
rect 14792 36036 14840 36092
rect 14896 36036 14944 36092
rect 15000 36036 15048 36092
rect 15104 36036 15152 36092
rect 15208 36036 15228 36092
rect 13988 34524 15228 36036
rect 13988 34468 14008 34524
rect 14064 34468 14112 34524
rect 14168 34468 14216 34524
rect 14272 34468 14320 34524
rect 14376 34468 14424 34524
rect 14480 34468 14528 34524
rect 14584 34468 14632 34524
rect 14688 34468 14736 34524
rect 14792 34468 14840 34524
rect 14896 34468 14944 34524
rect 15000 34468 15048 34524
rect 15104 34468 15152 34524
rect 15208 34468 15228 34524
rect 13988 32956 15228 34468
rect 13988 32900 14008 32956
rect 14064 32900 14112 32956
rect 14168 32900 14216 32956
rect 14272 32900 14320 32956
rect 14376 32900 14424 32956
rect 14480 32900 14528 32956
rect 14584 32900 14632 32956
rect 14688 32900 14736 32956
rect 14792 32900 14840 32956
rect 14896 32900 14944 32956
rect 15000 32900 15048 32956
rect 15104 32900 15152 32956
rect 15208 32900 15228 32956
rect 13988 31388 15228 32900
rect 13988 31332 14008 31388
rect 14064 31332 14112 31388
rect 14168 31332 14216 31388
rect 14272 31332 14320 31388
rect 14376 31332 14424 31388
rect 14480 31332 14528 31388
rect 14584 31332 14632 31388
rect 14688 31332 14736 31388
rect 14792 31332 14840 31388
rect 14896 31332 14944 31388
rect 15000 31332 15048 31388
rect 15104 31332 15152 31388
rect 15208 31332 15228 31388
rect 13988 29820 15228 31332
rect 13988 29764 14008 29820
rect 14064 29764 14112 29820
rect 14168 29764 14216 29820
rect 14272 29764 14320 29820
rect 14376 29764 14424 29820
rect 14480 29764 14528 29820
rect 14584 29764 14632 29820
rect 14688 29764 14736 29820
rect 14792 29764 14840 29820
rect 14896 29764 14944 29820
rect 15000 29764 15048 29820
rect 15104 29764 15152 29820
rect 15208 29764 15228 29820
rect 13988 28252 15228 29764
rect 13988 28196 14008 28252
rect 14064 28196 14112 28252
rect 14168 28196 14216 28252
rect 14272 28196 14320 28252
rect 14376 28196 14424 28252
rect 14480 28196 14528 28252
rect 14584 28196 14632 28252
rect 14688 28196 14736 28252
rect 14792 28196 14840 28252
rect 14896 28196 14944 28252
rect 15000 28196 15048 28252
rect 15104 28196 15152 28252
rect 15208 28196 15228 28252
rect 13988 26684 15228 28196
rect 13988 26628 14008 26684
rect 14064 26628 14112 26684
rect 14168 26628 14216 26684
rect 14272 26628 14320 26684
rect 14376 26628 14424 26684
rect 14480 26628 14528 26684
rect 14584 26628 14632 26684
rect 14688 26628 14736 26684
rect 14792 26628 14840 26684
rect 14896 26628 14944 26684
rect 15000 26628 15048 26684
rect 15104 26628 15152 26684
rect 15208 26628 15228 26684
rect 13988 25116 15228 26628
rect 13988 25060 14008 25116
rect 14064 25060 14112 25116
rect 14168 25060 14216 25116
rect 14272 25060 14320 25116
rect 14376 25060 14424 25116
rect 14480 25060 14528 25116
rect 14584 25060 14632 25116
rect 14688 25060 14736 25116
rect 14792 25060 14840 25116
rect 14896 25060 14944 25116
rect 15000 25060 15048 25116
rect 15104 25060 15152 25116
rect 15208 25060 15228 25116
rect 13988 23548 15228 25060
rect 13988 23492 14008 23548
rect 14064 23492 14112 23548
rect 14168 23492 14216 23548
rect 14272 23492 14320 23548
rect 14376 23492 14424 23548
rect 14480 23492 14528 23548
rect 14584 23492 14632 23548
rect 14688 23492 14736 23548
rect 14792 23492 14840 23548
rect 14896 23492 14944 23548
rect 15000 23492 15048 23548
rect 15104 23492 15152 23548
rect 15208 23492 15228 23548
rect 13988 21980 15228 23492
rect 13988 21924 14008 21980
rect 14064 21924 14112 21980
rect 14168 21924 14216 21980
rect 14272 21924 14320 21980
rect 14376 21924 14424 21980
rect 14480 21924 14528 21980
rect 14584 21924 14632 21980
rect 14688 21924 14736 21980
rect 14792 21924 14840 21980
rect 14896 21924 14944 21980
rect 15000 21924 15048 21980
rect 15104 21924 15152 21980
rect 15208 21924 15228 21980
rect 13988 20412 15228 21924
rect 13988 20356 14008 20412
rect 14064 20356 14112 20412
rect 14168 20356 14216 20412
rect 14272 20356 14320 20412
rect 14376 20356 14424 20412
rect 14480 20356 14528 20412
rect 14584 20356 14632 20412
rect 14688 20356 14736 20412
rect 14792 20356 14840 20412
rect 14896 20356 14944 20412
rect 15000 20356 15048 20412
rect 15104 20356 15152 20412
rect 15208 20356 15228 20412
rect 13988 18844 15228 20356
rect 13988 18788 14008 18844
rect 14064 18788 14112 18844
rect 14168 18788 14216 18844
rect 14272 18788 14320 18844
rect 14376 18788 14424 18844
rect 14480 18788 14528 18844
rect 14584 18788 14632 18844
rect 14688 18788 14736 18844
rect 14792 18788 14840 18844
rect 14896 18788 14944 18844
rect 15000 18788 15048 18844
rect 15104 18788 15152 18844
rect 15208 18788 15228 18844
rect 13988 17276 15228 18788
rect 13988 17220 14008 17276
rect 14064 17220 14112 17276
rect 14168 17220 14216 17276
rect 14272 17220 14320 17276
rect 14376 17220 14424 17276
rect 14480 17220 14528 17276
rect 14584 17220 14632 17276
rect 14688 17220 14736 17276
rect 14792 17220 14840 17276
rect 14896 17220 14944 17276
rect 15000 17220 15048 17276
rect 15104 17220 15152 17276
rect 15208 17220 15228 17276
rect 13988 15708 15228 17220
rect 13988 15652 14008 15708
rect 14064 15652 14112 15708
rect 14168 15652 14216 15708
rect 14272 15652 14320 15708
rect 14376 15652 14424 15708
rect 14480 15652 14528 15708
rect 14584 15652 14632 15708
rect 14688 15652 14736 15708
rect 14792 15652 14840 15708
rect 14896 15652 14944 15708
rect 15000 15652 15048 15708
rect 15104 15652 15152 15708
rect 15208 15652 15228 15708
rect 13988 14140 15228 15652
rect 13988 14084 14008 14140
rect 14064 14084 14112 14140
rect 14168 14084 14216 14140
rect 14272 14084 14320 14140
rect 14376 14084 14424 14140
rect 14480 14084 14528 14140
rect 14584 14084 14632 14140
rect 14688 14084 14736 14140
rect 14792 14084 14840 14140
rect 14896 14084 14944 14140
rect 15000 14084 15048 14140
rect 15104 14084 15152 14140
rect 15208 14084 15228 14140
rect 13988 12572 15228 14084
rect 13988 12516 14008 12572
rect 14064 12516 14112 12572
rect 14168 12516 14216 12572
rect 14272 12516 14320 12572
rect 14376 12516 14424 12572
rect 14480 12516 14528 12572
rect 14584 12516 14632 12572
rect 14688 12516 14736 12572
rect 14792 12516 14840 12572
rect 14896 12516 14944 12572
rect 15000 12516 15048 12572
rect 15104 12516 15152 12572
rect 15208 12516 15228 12572
rect 13988 11004 15228 12516
rect 13988 10948 14008 11004
rect 14064 10948 14112 11004
rect 14168 10948 14216 11004
rect 14272 10948 14320 11004
rect 14376 10948 14424 11004
rect 14480 10948 14528 11004
rect 14584 10948 14632 11004
rect 14688 10948 14736 11004
rect 14792 10948 14840 11004
rect 14896 10948 14944 11004
rect 15000 10948 15048 11004
rect 15104 10948 15152 11004
rect 15208 10948 15228 11004
rect 13988 9436 15228 10948
rect 13988 9380 14008 9436
rect 14064 9380 14112 9436
rect 14168 9380 14216 9436
rect 14272 9380 14320 9436
rect 14376 9380 14424 9436
rect 14480 9380 14528 9436
rect 14584 9380 14632 9436
rect 14688 9380 14736 9436
rect 14792 9380 14840 9436
rect 14896 9380 14944 9436
rect 15000 9380 15048 9436
rect 15104 9380 15152 9436
rect 15208 9380 15228 9436
rect 3988 8596 4008 8652
rect 4064 8596 4112 8652
rect 4168 8596 4216 8652
rect 4272 8596 4320 8652
rect 4376 8596 4424 8652
rect 4480 8596 4528 8652
rect 4584 8596 4632 8652
rect 4688 8596 4736 8652
rect 4792 8596 4840 8652
rect 4896 8596 4944 8652
rect 5000 8596 5048 8652
rect 5104 8596 5152 8652
rect 5208 8596 5228 8652
rect 3988 7084 5228 8596
rect 7420 8708 7476 8718
rect 3988 7028 4008 7084
rect 4064 7028 4112 7084
rect 4168 7028 4216 7084
rect 4272 7028 4320 7084
rect 4376 7028 4424 7084
rect 4480 7028 4528 7084
rect 4584 7028 4632 7084
rect 4688 7028 4736 7084
rect 4792 7028 4840 7084
rect 4896 7028 4944 7084
rect 5000 7028 5048 7084
rect 5104 7028 5152 7084
rect 5208 7028 5228 7084
rect 3988 5516 5228 7028
rect 3988 5460 4008 5516
rect 4064 5460 4112 5516
rect 4168 5460 4216 5516
rect 4272 5460 4320 5516
rect 4376 5460 4424 5516
rect 4480 5460 4528 5516
rect 4584 5460 4632 5516
rect 4688 5460 4736 5516
rect 4792 5460 4840 5516
rect 4896 5460 4944 5516
rect 5000 5460 5048 5516
rect 5104 5460 5152 5516
rect 5208 5460 5228 5516
rect 3988 3948 5228 5460
rect 5628 8260 5684 8270
rect 5628 5684 5684 8204
rect 6524 8036 6580 8046
rect 5740 7140 5796 7150
rect 5740 6020 5796 7084
rect 5740 5954 5796 5964
rect 6188 6244 6244 6254
rect 5628 5012 5684 5628
rect 5628 4946 5684 4956
rect 6188 4900 6244 6188
rect 6188 4834 6244 4844
rect 3988 3892 4008 3948
rect 4064 3892 4112 3948
rect 4168 3892 4216 3948
rect 4272 3892 4320 3948
rect 4376 3892 4424 3948
rect 4480 3892 4528 3948
rect 4584 3892 4632 3948
rect 4688 3892 4736 3948
rect 4792 3892 4840 3948
rect 4896 3892 4944 3948
rect 5000 3892 5048 3948
rect 5104 3892 5152 3948
rect 5208 3892 5228 3948
rect 3988 3076 5228 3892
rect 6524 3780 6580 7980
rect 6524 3714 6580 3724
rect 6972 8036 7028 8046
rect 6972 3332 7028 7980
rect 7084 7476 7140 7486
rect 7084 6244 7140 7420
rect 7420 6916 7476 8652
rect 7420 6356 7476 6860
rect 13988 7868 15228 9380
rect 13988 7812 14008 7868
rect 14064 7812 14112 7868
rect 14168 7812 14216 7868
rect 14272 7812 14320 7868
rect 14376 7812 14424 7868
rect 14480 7812 14528 7868
rect 14584 7812 14632 7868
rect 14688 7812 14736 7868
rect 14792 7812 14840 7868
rect 14896 7812 14944 7868
rect 15000 7812 15048 7868
rect 15104 7812 15152 7868
rect 15208 7812 15228 7868
rect 7420 6290 7476 6300
rect 7980 6692 8036 6702
rect 7084 6178 7140 6188
rect 7980 6244 8036 6636
rect 7980 6178 8036 6188
rect 13988 6300 15228 7812
rect 13988 6244 14008 6300
rect 14064 6244 14112 6300
rect 14168 6244 14216 6300
rect 14272 6244 14320 6300
rect 14376 6244 14424 6300
rect 14480 6244 14528 6300
rect 14584 6244 14632 6300
rect 14688 6244 14736 6300
rect 14792 6244 14840 6300
rect 14896 6244 14944 6300
rect 15000 6244 15048 6300
rect 15104 6244 15152 6300
rect 15208 6244 15228 6300
rect 6972 3266 7028 3276
rect 13988 4732 15228 6244
rect 23988 46284 25228 46316
rect 23988 46228 24008 46284
rect 24064 46228 24112 46284
rect 24168 46228 24216 46284
rect 24272 46228 24320 46284
rect 24376 46228 24424 46284
rect 24480 46228 24528 46284
rect 24584 46228 24632 46284
rect 24688 46228 24736 46284
rect 24792 46228 24840 46284
rect 24896 46228 24944 46284
rect 25000 46228 25048 46284
rect 25104 46228 25152 46284
rect 25208 46228 25228 46284
rect 23988 44716 25228 46228
rect 23988 44660 24008 44716
rect 24064 44660 24112 44716
rect 24168 44660 24216 44716
rect 24272 44660 24320 44716
rect 24376 44660 24424 44716
rect 24480 44660 24528 44716
rect 24584 44660 24632 44716
rect 24688 44660 24736 44716
rect 24792 44660 24840 44716
rect 24896 44660 24944 44716
rect 25000 44660 25048 44716
rect 25104 44660 25152 44716
rect 25208 44660 25228 44716
rect 23988 43148 25228 44660
rect 23988 43092 24008 43148
rect 24064 43092 24112 43148
rect 24168 43092 24216 43148
rect 24272 43092 24320 43148
rect 24376 43092 24424 43148
rect 24480 43092 24528 43148
rect 24584 43092 24632 43148
rect 24688 43092 24736 43148
rect 24792 43092 24840 43148
rect 24896 43092 24944 43148
rect 25000 43092 25048 43148
rect 25104 43092 25152 43148
rect 25208 43092 25228 43148
rect 23988 41580 25228 43092
rect 23988 41524 24008 41580
rect 24064 41524 24112 41580
rect 24168 41524 24216 41580
rect 24272 41524 24320 41580
rect 24376 41524 24424 41580
rect 24480 41524 24528 41580
rect 24584 41524 24632 41580
rect 24688 41524 24736 41580
rect 24792 41524 24840 41580
rect 24896 41524 24944 41580
rect 25000 41524 25048 41580
rect 25104 41524 25152 41580
rect 25208 41524 25228 41580
rect 23988 40012 25228 41524
rect 23988 39956 24008 40012
rect 24064 39956 24112 40012
rect 24168 39956 24216 40012
rect 24272 39956 24320 40012
rect 24376 39956 24424 40012
rect 24480 39956 24528 40012
rect 24584 39956 24632 40012
rect 24688 39956 24736 40012
rect 24792 39956 24840 40012
rect 24896 39956 24944 40012
rect 25000 39956 25048 40012
rect 25104 39956 25152 40012
rect 25208 39956 25228 40012
rect 23988 38444 25228 39956
rect 23988 38388 24008 38444
rect 24064 38388 24112 38444
rect 24168 38388 24216 38444
rect 24272 38388 24320 38444
rect 24376 38388 24424 38444
rect 24480 38388 24528 38444
rect 24584 38388 24632 38444
rect 24688 38388 24736 38444
rect 24792 38388 24840 38444
rect 24896 38388 24944 38444
rect 25000 38388 25048 38444
rect 25104 38388 25152 38444
rect 25208 38388 25228 38444
rect 23988 36876 25228 38388
rect 23988 36820 24008 36876
rect 24064 36820 24112 36876
rect 24168 36820 24216 36876
rect 24272 36820 24320 36876
rect 24376 36820 24424 36876
rect 24480 36820 24528 36876
rect 24584 36820 24632 36876
rect 24688 36820 24736 36876
rect 24792 36820 24840 36876
rect 24896 36820 24944 36876
rect 25000 36820 25048 36876
rect 25104 36820 25152 36876
rect 25208 36820 25228 36876
rect 23988 35308 25228 36820
rect 23988 35252 24008 35308
rect 24064 35252 24112 35308
rect 24168 35252 24216 35308
rect 24272 35252 24320 35308
rect 24376 35252 24424 35308
rect 24480 35252 24528 35308
rect 24584 35252 24632 35308
rect 24688 35252 24736 35308
rect 24792 35252 24840 35308
rect 24896 35252 24944 35308
rect 25000 35252 25048 35308
rect 25104 35252 25152 35308
rect 25208 35252 25228 35308
rect 23988 33740 25228 35252
rect 23988 33684 24008 33740
rect 24064 33684 24112 33740
rect 24168 33684 24216 33740
rect 24272 33684 24320 33740
rect 24376 33684 24424 33740
rect 24480 33684 24528 33740
rect 24584 33684 24632 33740
rect 24688 33684 24736 33740
rect 24792 33684 24840 33740
rect 24896 33684 24944 33740
rect 25000 33684 25048 33740
rect 25104 33684 25152 33740
rect 25208 33684 25228 33740
rect 23988 32172 25228 33684
rect 23988 32116 24008 32172
rect 24064 32116 24112 32172
rect 24168 32116 24216 32172
rect 24272 32116 24320 32172
rect 24376 32116 24424 32172
rect 24480 32116 24528 32172
rect 24584 32116 24632 32172
rect 24688 32116 24736 32172
rect 24792 32116 24840 32172
rect 24896 32116 24944 32172
rect 25000 32116 25048 32172
rect 25104 32116 25152 32172
rect 25208 32116 25228 32172
rect 23988 30604 25228 32116
rect 23988 30548 24008 30604
rect 24064 30548 24112 30604
rect 24168 30548 24216 30604
rect 24272 30548 24320 30604
rect 24376 30548 24424 30604
rect 24480 30548 24528 30604
rect 24584 30548 24632 30604
rect 24688 30548 24736 30604
rect 24792 30548 24840 30604
rect 24896 30548 24944 30604
rect 25000 30548 25048 30604
rect 25104 30548 25152 30604
rect 25208 30548 25228 30604
rect 23988 29036 25228 30548
rect 23988 28980 24008 29036
rect 24064 28980 24112 29036
rect 24168 28980 24216 29036
rect 24272 28980 24320 29036
rect 24376 28980 24424 29036
rect 24480 28980 24528 29036
rect 24584 28980 24632 29036
rect 24688 28980 24736 29036
rect 24792 28980 24840 29036
rect 24896 28980 24944 29036
rect 25000 28980 25048 29036
rect 25104 28980 25152 29036
rect 25208 28980 25228 29036
rect 23988 27468 25228 28980
rect 23988 27412 24008 27468
rect 24064 27412 24112 27468
rect 24168 27412 24216 27468
rect 24272 27412 24320 27468
rect 24376 27412 24424 27468
rect 24480 27412 24528 27468
rect 24584 27412 24632 27468
rect 24688 27412 24736 27468
rect 24792 27412 24840 27468
rect 24896 27412 24944 27468
rect 25000 27412 25048 27468
rect 25104 27412 25152 27468
rect 25208 27412 25228 27468
rect 23988 25900 25228 27412
rect 23988 25844 24008 25900
rect 24064 25844 24112 25900
rect 24168 25844 24216 25900
rect 24272 25844 24320 25900
rect 24376 25844 24424 25900
rect 24480 25844 24528 25900
rect 24584 25844 24632 25900
rect 24688 25844 24736 25900
rect 24792 25844 24840 25900
rect 24896 25844 24944 25900
rect 25000 25844 25048 25900
rect 25104 25844 25152 25900
rect 25208 25844 25228 25900
rect 23988 24332 25228 25844
rect 23988 24276 24008 24332
rect 24064 24276 24112 24332
rect 24168 24276 24216 24332
rect 24272 24276 24320 24332
rect 24376 24276 24424 24332
rect 24480 24276 24528 24332
rect 24584 24276 24632 24332
rect 24688 24276 24736 24332
rect 24792 24276 24840 24332
rect 24896 24276 24944 24332
rect 25000 24276 25048 24332
rect 25104 24276 25152 24332
rect 25208 24276 25228 24332
rect 23988 22764 25228 24276
rect 23988 22708 24008 22764
rect 24064 22708 24112 22764
rect 24168 22708 24216 22764
rect 24272 22708 24320 22764
rect 24376 22708 24424 22764
rect 24480 22708 24528 22764
rect 24584 22708 24632 22764
rect 24688 22708 24736 22764
rect 24792 22708 24840 22764
rect 24896 22708 24944 22764
rect 25000 22708 25048 22764
rect 25104 22708 25152 22764
rect 25208 22708 25228 22764
rect 23988 21196 25228 22708
rect 23988 21140 24008 21196
rect 24064 21140 24112 21196
rect 24168 21140 24216 21196
rect 24272 21140 24320 21196
rect 24376 21140 24424 21196
rect 24480 21140 24528 21196
rect 24584 21140 24632 21196
rect 24688 21140 24736 21196
rect 24792 21140 24840 21196
rect 24896 21140 24944 21196
rect 25000 21140 25048 21196
rect 25104 21140 25152 21196
rect 25208 21140 25228 21196
rect 23988 19628 25228 21140
rect 23988 19572 24008 19628
rect 24064 19572 24112 19628
rect 24168 19572 24216 19628
rect 24272 19572 24320 19628
rect 24376 19572 24424 19628
rect 24480 19572 24528 19628
rect 24584 19572 24632 19628
rect 24688 19572 24736 19628
rect 24792 19572 24840 19628
rect 24896 19572 24944 19628
rect 25000 19572 25048 19628
rect 25104 19572 25152 19628
rect 25208 19572 25228 19628
rect 23988 18060 25228 19572
rect 23988 18004 24008 18060
rect 24064 18004 24112 18060
rect 24168 18004 24216 18060
rect 24272 18004 24320 18060
rect 24376 18004 24424 18060
rect 24480 18004 24528 18060
rect 24584 18004 24632 18060
rect 24688 18004 24736 18060
rect 24792 18004 24840 18060
rect 24896 18004 24944 18060
rect 25000 18004 25048 18060
rect 25104 18004 25152 18060
rect 25208 18004 25228 18060
rect 23988 16492 25228 18004
rect 23988 16436 24008 16492
rect 24064 16436 24112 16492
rect 24168 16436 24216 16492
rect 24272 16436 24320 16492
rect 24376 16436 24424 16492
rect 24480 16436 24528 16492
rect 24584 16436 24632 16492
rect 24688 16436 24736 16492
rect 24792 16436 24840 16492
rect 24896 16436 24944 16492
rect 25000 16436 25048 16492
rect 25104 16436 25152 16492
rect 25208 16436 25228 16492
rect 23988 14924 25228 16436
rect 23988 14868 24008 14924
rect 24064 14868 24112 14924
rect 24168 14868 24216 14924
rect 24272 14868 24320 14924
rect 24376 14868 24424 14924
rect 24480 14868 24528 14924
rect 24584 14868 24632 14924
rect 24688 14868 24736 14924
rect 24792 14868 24840 14924
rect 24896 14868 24944 14924
rect 25000 14868 25048 14924
rect 25104 14868 25152 14924
rect 25208 14868 25228 14924
rect 23988 13356 25228 14868
rect 23988 13300 24008 13356
rect 24064 13300 24112 13356
rect 24168 13300 24216 13356
rect 24272 13300 24320 13356
rect 24376 13300 24424 13356
rect 24480 13300 24528 13356
rect 24584 13300 24632 13356
rect 24688 13300 24736 13356
rect 24792 13300 24840 13356
rect 24896 13300 24944 13356
rect 25000 13300 25048 13356
rect 25104 13300 25152 13356
rect 25208 13300 25228 13356
rect 23988 11788 25228 13300
rect 23988 11732 24008 11788
rect 24064 11732 24112 11788
rect 24168 11732 24216 11788
rect 24272 11732 24320 11788
rect 24376 11732 24424 11788
rect 24480 11732 24528 11788
rect 24584 11732 24632 11788
rect 24688 11732 24736 11788
rect 24792 11732 24840 11788
rect 24896 11732 24944 11788
rect 25000 11732 25048 11788
rect 25104 11732 25152 11788
rect 25208 11732 25228 11788
rect 23988 10220 25228 11732
rect 23988 10164 24008 10220
rect 24064 10164 24112 10220
rect 24168 10164 24216 10220
rect 24272 10164 24320 10220
rect 24376 10164 24424 10220
rect 24480 10164 24528 10220
rect 24584 10164 24632 10220
rect 24688 10164 24736 10220
rect 24792 10164 24840 10220
rect 24896 10164 24944 10220
rect 25000 10164 25048 10220
rect 25104 10164 25152 10220
rect 25208 10164 25228 10220
rect 23988 8652 25228 10164
rect 23988 8596 24008 8652
rect 24064 8596 24112 8652
rect 24168 8596 24216 8652
rect 24272 8596 24320 8652
rect 24376 8596 24424 8652
rect 24480 8596 24528 8652
rect 24584 8596 24632 8652
rect 24688 8596 24736 8652
rect 24792 8596 24840 8652
rect 24896 8596 24944 8652
rect 25000 8596 25048 8652
rect 25104 8596 25152 8652
rect 25208 8596 25228 8652
rect 23988 7084 25228 8596
rect 23988 7028 24008 7084
rect 24064 7028 24112 7084
rect 24168 7028 24216 7084
rect 24272 7028 24320 7084
rect 24376 7028 24424 7084
rect 24480 7028 24528 7084
rect 24584 7028 24632 7084
rect 24688 7028 24736 7084
rect 24792 7028 24840 7084
rect 24896 7028 24944 7084
rect 25000 7028 25048 7084
rect 25104 7028 25152 7084
rect 25208 7028 25228 7084
rect 23988 5516 25228 7028
rect 23988 5460 24008 5516
rect 24064 5460 24112 5516
rect 24168 5460 24216 5516
rect 24272 5460 24320 5516
rect 24376 5460 24424 5516
rect 24480 5460 24528 5516
rect 24584 5460 24632 5516
rect 24688 5460 24736 5516
rect 24792 5460 24840 5516
rect 24896 5460 24944 5516
rect 25000 5460 25048 5516
rect 25104 5460 25152 5516
rect 25208 5460 25228 5516
rect 13988 4676 14008 4732
rect 14064 4676 14112 4732
rect 14168 4676 14216 4732
rect 14272 4676 14320 4732
rect 14376 4676 14424 4732
rect 14480 4676 14528 4732
rect 14584 4676 14632 4732
rect 14688 4676 14736 4732
rect 14792 4676 14840 4732
rect 14896 4676 14944 4732
rect 15000 4676 15048 4732
rect 15104 4676 15152 4732
rect 15208 4676 15228 4732
rect 13988 3164 15228 4676
rect 15708 4788 15764 4798
rect 15708 4004 15764 4732
rect 15708 3938 15764 3948
rect 23988 3948 25228 5460
rect 13988 3108 14008 3164
rect 14064 3108 14112 3164
rect 14168 3108 14216 3164
rect 14272 3108 14320 3164
rect 14376 3108 14424 3164
rect 14480 3108 14528 3164
rect 14584 3108 14632 3164
rect 14688 3108 14736 3164
rect 14792 3108 14840 3164
rect 14896 3108 14944 3164
rect 15000 3108 15048 3164
rect 15104 3108 15152 3164
rect 15208 3108 15228 3164
rect 13988 3076 15228 3108
rect 23988 3892 24008 3948
rect 24064 3892 24112 3948
rect 24168 3892 24216 3948
rect 24272 3892 24320 3948
rect 24376 3892 24424 3948
rect 24480 3892 24528 3948
rect 24584 3892 24632 3948
rect 24688 3892 24736 3948
rect 24792 3892 24840 3948
rect 24896 3892 24944 3948
rect 25000 3892 25048 3948
rect 25104 3892 25152 3948
rect 25208 3892 25228 3948
rect 23988 3076 25228 3892
rect 33988 45500 35228 46316
rect 33988 45444 34008 45500
rect 34064 45444 34112 45500
rect 34168 45444 34216 45500
rect 34272 45444 34320 45500
rect 34376 45444 34424 45500
rect 34480 45444 34528 45500
rect 34584 45444 34632 45500
rect 34688 45444 34736 45500
rect 34792 45444 34840 45500
rect 34896 45444 34944 45500
rect 35000 45444 35048 45500
rect 35104 45444 35152 45500
rect 35208 45444 35228 45500
rect 33988 43932 35228 45444
rect 33988 43876 34008 43932
rect 34064 43876 34112 43932
rect 34168 43876 34216 43932
rect 34272 43876 34320 43932
rect 34376 43876 34424 43932
rect 34480 43876 34528 43932
rect 34584 43876 34632 43932
rect 34688 43876 34736 43932
rect 34792 43876 34840 43932
rect 34896 43876 34944 43932
rect 35000 43876 35048 43932
rect 35104 43876 35152 43932
rect 35208 43876 35228 43932
rect 33988 42364 35228 43876
rect 33988 42308 34008 42364
rect 34064 42308 34112 42364
rect 34168 42308 34216 42364
rect 34272 42308 34320 42364
rect 34376 42308 34424 42364
rect 34480 42308 34528 42364
rect 34584 42308 34632 42364
rect 34688 42308 34736 42364
rect 34792 42308 34840 42364
rect 34896 42308 34944 42364
rect 35000 42308 35048 42364
rect 35104 42308 35152 42364
rect 35208 42308 35228 42364
rect 33988 40796 35228 42308
rect 33988 40740 34008 40796
rect 34064 40740 34112 40796
rect 34168 40740 34216 40796
rect 34272 40740 34320 40796
rect 34376 40740 34424 40796
rect 34480 40740 34528 40796
rect 34584 40740 34632 40796
rect 34688 40740 34736 40796
rect 34792 40740 34840 40796
rect 34896 40740 34944 40796
rect 35000 40740 35048 40796
rect 35104 40740 35152 40796
rect 35208 40740 35228 40796
rect 33988 39228 35228 40740
rect 33988 39172 34008 39228
rect 34064 39172 34112 39228
rect 34168 39172 34216 39228
rect 34272 39172 34320 39228
rect 34376 39172 34424 39228
rect 34480 39172 34528 39228
rect 34584 39172 34632 39228
rect 34688 39172 34736 39228
rect 34792 39172 34840 39228
rect 34896 39172 34944 39228
rect 35000 39172 35048 39228
rect 35104 39172 35152 39228
rect 35208 39172 35228 39228
rect 33988 37660 35228 39172
rect 33988 37604 34008 37660
rect 34064 37604 34112 37660
rect 34168 37604 34216 37660
rect 34272 37604 34320 37660
rect 34376 37604 34424 37660
rect 34480 37604 34528 37660
rect 34584 37604 34632 37660
rect 34688 37604 34736 37660
rect 34792 37604 34840 37660
rect 34896 37604 34944 37660
rect 35000 37604 35048 37660
rect 35104 37604 35152 37660
rect 35208 37604 35228 37660
rect 33988 36092 35228 37604
rect 33988 36036 34008 36092
rect 34064 36036 34112 36092
rect 34168 36036 34216 36092
rect 34272 36036 34320 36092
rect 34376 36036 34424 36092
rect 34480 36036 34528 36092
rect 34584 36036 34632 36092
rect 34688 36036 34736 36092
rect 34792 36036 34840 36092
rect 34896 36036 34944 36092
rect 35000 36036 35048 36092
rect 35104 36036 35152 36092
rect 35208 36036 35228 36092
rect 33988 34524 35228 36036
rect 33988 34468 34008 34524
rect 34064 34468 34112 34524
rect 34168 34468 34216 34524
rect 34272 34468 34320 34524
rect 34376 34468 34424 34524
rect 34480 34468 34528 34524
rect 34584 34468 34632 34524
rect 34688 34468 34736 34524
rect 34792 34468 34840 34524
rect 34896 34468 34944 34524
rect 35000 34468 35048 34524
rect 35104 34468 35152 34524
rect 35208 34468 35228 34524
rect 33988 32956 35228 34468
rect 33988 32900 34008 32956
rect 34064 32900 34112 32956
rect 34168 32900 34216 32956
rect 34272 32900 34320 32956
rect 34376 32900 34424 32956
rect 34480 32900 34528 32956
rect 34584 32900 34632 32956
rect 34688 32900 34736 32956
rect 34792 32900 34840 32956
rect 34896 32900 34944 32956
rect 35000 32900 35048 32956
rect 35104 32900 35152 32956
rect 35208 32900 35228 32956
rect 33988 31388 35228 32900
rect 33988 31332 34008 31388
rect 34064 31332 34112 31388
rect 34168 31332 34216 31388
rect 34272 31332 34320 31388
rect 34376 31332 34424 31388
rect 34480 31332 34528 31388
rect 34584 31332 34632 31388
rect 34688 31332 34736 31388
rect 34792 31332 34840 31388
rect 34896 31332 34944 31388
rect 35000 31332 35048 31388
rect 35104 31332 35152 31388
rect 35208 31332 35228 31388
rect 33988 29820 35228 31332
rect 33988 29764 34008 29820
rect 34064 29764 34112 29820
rect 34168 29764 34216 29820
rect 34272 29764 34320 29820
rect 34376 29764 34424 29820
rect 34480 29764 34528 29820
rect 34584 29764 34632 29820
rect 34688 29764 34736 29820
rect 34792 29764 34840 29820
rect 34896 29764 34944 29820
rect 35000 29764 35048 29820
rect 35104 29764 35152 29820
rect 35208 29764 35228 29820
rect 33988 28252 35228 29764
rect 33988 28196 34008 28252
rect 34064 28196 34112 28252
rect 34168 28196 34216 28252
rect 34272 28196 34320 28252
rect 34376 28196 34424 28252
rect 34480 28196 34528 28252
rect 34584 28196 34632 28252
rect 34688 28196 34736 28252
rect 34792 28196 34840 28252
rect 34896 28196 34944 28252
rect 35000 28196 35048 28252
rect 35104 28196 35152 28252
rect 35208 28196 35228 28252
rect 33988 26684 35228 28196
rect 33988 26628 34008 26684
rect 34064 26628 34112 26684
rect 34168 26628 34216 26684
rect 34272 26628 34320 26684
rect 34376 26628 34424 26684
rect 34480 26628 34528 26684
rect 34584 26628 34632 26684
rect 34688 26628 34736 26684
rect 34792 26628 34840 26684
rect 34896 26628 34944 26684
rect 35000 26628 35048 26684
rect 35104 26628 35152 26684
rect 35208 26628 35228 26684
rect 33988 25116 35228 26628
rect 33988 25060 34008 25116
rect 34064 25060 34112 25116
rect 34168 25060 34216 25116
rect 34272 25060 34320 25116
rect 34376 25060 34424 25116
rect 34480 25060 34528 25116
rect 34584 25060 34632 25116
rect 34688 25060 34736 25116
rect 34792 25060 34840 25116
rect 34896 25060 34944 25116
rect 35000 25060 35048 25116
rect 35104 25060 35152 25116
rect 35208 25060 35228 25116
rect 33988 23548 35228 25060
rect 33988 23492 34008 23548
rect 34064 23492 34112 23548
rect 34168 23492 34216 23548
rect 34272 23492 34320 23548
rect 34376 23492 34424 23548
rect 34480 23492 34528 23548
rect 34584 23492 34632 23548
rect 34688 23492 34736 23548
rect 34792 23492 34840 23548
rect 34896 23492 34944 23548
rect 35000 23492 35048 23548
rect 35104 23492 35152 23548
rect 35208 23492 35228 23548
rect 33988 21980 35228 23492
rect 33988 21924 34008 21980
rect 34064 21924 34112 21980
rect 34168 21924 34216 21980
rect 34272 21924 34320 21980
rect 34376 21924 34424 21980
rect 34480 21924 34528 21980
rect 34584 21924 34632 21980
rect 34688 21924 34736 21980
rect 34792 21924 34840 21980
rect 34896 21924 34944 21980
rect 35000 21924 35048 21980
rect 35104 21924 35152 21980
rect 35208 21924 35228 21980
rect 33988 20412 35228 21924
rect 33988 20356 34008 20412
rect 34064 20356 34112 20412
rect 34168 20356 34216 20412
rect 34272 20356 34320 20412
rect 34376 20356 34424 20412
rect 34480 20356 34528 20412
rect 34584 20356 34632 20412
rect 34688 20356 34736 20412
rect 34792 20356 34840 20412
rect 34896 20356 34944 20412
rect 35000 20356 35048 20412
rect 35104 20356 35152 20412
rect 35208 20356 35228 20412
rect 33988 18844 35228 20356
rect 33988 18788 34008 18844
rect 34064 18788 34112 18844
rect 34168 18788 34216 18844
rect 34272 18788 34320 18844
rect 34376 18788 34424 18844
rect 34480 18788 34528 18844
rect 34584 18788 34632 18844
rect 34688 18788 34736 18844
rect 34792 18788 34840 18844
rect 34896 18788 34944 18844
rect 35000 18788 35048 18844
rect 35104 18788 35152 18844
rect 35208 18788 35228 18844
rect 33988 17276 35228 18788
rect 33988 17220 34008 17276
rect 34064 17220 34112 17276
rect 34168 17220 34216 17276
rect 34272 17220 34320 17276
rect 34376 17220 34424 17276
rect 34480 17220 34528 17276
rect 34584 17220 34632 17276
rect 34688 17220 34736 17276
rect 34792 17220 34840 17276
rect 34896 17220 34944 17276
rect 35000 17220 35048 17276
rect 35104 17220 35152 17276
rect 35208 17220 35228 17276
rect 33988 15708 35228 17220
rect 33988 15652 34008 15708
rect 34064 15652 34112 15708
rect 34168 15652 34216 15708
rect 34272 15652 34320 15708
rect 34376 15652 34424 15708
rect 34480 15652 34528 15708
rect 34584 15652 34632 15708
rect 34688 15652 34736 15708
rect 34792 15652 34840 15708
rect 34896 15652 34944 15708
rect 35000 15652 35048 15708
rect 35104 15652 35152 15708
rect 35208 15652 35228 15708
rect 33988 14140 35228 15652
rect 33988 14084 34008 14140
rect 34064 14084 34112 14140
rect 34168 14084 34216 14140
rect 34272 14084 34320 14140
rect 34376 14084 34424 14140
rect 34480 14084 34528 14140
rect 34584 14084 34632 14140
rect 34688 14084 34736 14140
rect 34792 14084 34840 14140
rect 34896 14084 34944 14140
rect 35000 14084 35048 14140
rect 35104 14084 35152 14140
rect 35208 14084 35228 14140
rect 33988 12572 35228 14084
rect 33988 12516 34008 12572
rect 34064 12516 34112 12572
rect 34168 12516 34216 12572
rect 34272 12516 34320 12572
rect 34376 12516 34424 12572
rect 34480 12516 34528 12572
rect 34584 12516 34632 12572
rect 34688 12516 34736 12572
rect 34792 12516 34840 12572
rect 34896 12516 34944 12572
rect 35000 12516 35048 12572
rect 35104 12516 35152 12572
rect 35208 12516 35228 12572
rect 33988 11004 35228 12516
rect 33988 10948 34008 11004
rect 34064 10948 34112 11004
rect 34168 10948 34216 11004
rect 34272 10948 34320 11004
rect 34376 10948 34424 11004
rect 34480 10948 34528 11004
rect 34584 10948 34632 11004
rect 34688 10948 34736 11004
rect 34792 10948 34840 11004
rect 34896 10948 34944 11004
rect 35000 10948 35048 11004
rect 35104 10948 35152 11004
rect 35208 10948 35228 11004
rect 33988 9436 35228 10948
rect 33988 9380 34008 9436
rect 34064 9380 34112 9436
rect 34168 9380 34216 9436
rect 34272 9380 34320 9436
rect 34376 9380 34424 9436
rect 34480 9380 34528 9436
rect 34584 9380 34632 9436
rect 34688 9380 34736 9436
rect 34792 9380 34840 9436
rect 34896 9380 34944 9436
rect 35000 9380 35048 9436
rect 35104 9380 35152 9436
rect 35208 9380 35228 9436
rect 33988 7868 35228 9380
rect 33988 7812 34008 7868
rect 34064 7812 34112 7868
rect 34168 7812 34216 7868
rect 34272 7812 34320 7868
rect 34376 7812 34424 7868
rect 34480 7812 34528 7868
rect 34584 7812 34632 7868
rect 34688 7812 34736 7868
rect 34792 7812 34840 7868
rect 34896 7812 34944 7868
rect 35000 7812 35048 7868
rect 35104 7812 35152 7868
rect 35208 7812 35228 7868
rect 33988 6300 35228 7812
rect 33988 6244 34008 6300
rect 34064 6244 34112 6300
rect 34168 6244 34216 6300
rect 34272 6244 34320 6300
rect 34376 6244 34424 6300
rect 34480 6244 34528 6300
rect 34584 6244 34632 6300
rect 34688 6244 34736 6300
rect 34792 6244 34840 6300
rect 34896 6244 34944 6300
rect 35000 6244 35048 6300
rect 35104 6244 35152 6300
rect 35208 6244 35228 6300
rect 33988 4732 35228 6244
rect 33988 4676 34008 4732
rect 34064 4676 34112 4732
rect 34168 4676 34216 4732
rect 34272 4676 34320 4732
rect 34376 4676 34424 4732
rect 34480 4676 34528 4732
rect 34584 4676 34632 4732
rect 34688 4676 34736 4732
rect 34792 4676 34840 4732
rect 34896 4676 34944 4732
rect 35000 4676 35048 4732
rect 35104 4676 35152 4732
rect 35208 4676 35228 4732
rect 33988 3164 35228 4676
rect 33988 3108 34008 3164
rect 34064 3108 34112 3164
rect 34168 3108 34216 3164
rect 34272 3108 34320 3164
rect 34376 3108 34424 3164
rect 34480 3108 34528 3164
rect 34584 3108 34632 3164
rect 34688 3108 34736 3164
rect 34792 3108 34840 3164
rect 34896 3108 34944 3164
rect 35000 3108 35048 3164
rect 35104 3108 35152 3164
rect 35208 3108 35228 3164
rect 33988 3076 35228 3108
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _042_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 7840 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _043_
timestamp 1698431365
transform -1 0 11424 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _044_
timestamp 1698431365
transform 1 0 9184 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _045_
timestamp 1698431365
transform -1 0 7952 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _046_
timestamp 1698431365
transform -1 0 7952 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _047_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 17920 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _048_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 22176 0 -1 4704
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _049_
timestamp 1698431365
transform -1 0 18368 0 1 4704
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _050_
timestamp 1698431365
transform 1 0 13328 0 1 6272
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  _051_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 15904 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _052_
timestamp 1698431365
transform -1 0 29232 0 -1 4704
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _053_
timestamp 1698431365
transform -1 0 26208 0 1 4704
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  _054_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 24304 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _055_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 34944 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _056_
timestamp 1698431365
transform -1 0 34160 0 1 4704
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _057_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 35616 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _058_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 9408 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _059_
timestamp 1698431365
transform 1 0 8512 0 1 6272
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _060_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 12768 0 1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _061_
timestamp 1698431365
transform 1 0 8960 0 1 7840
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _062_
timestamp 1698431365
transform 1 0 6048 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _063_
timestamp 1698431365
transform 1 0 9856 0 -1 7840
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _064_
timestamp 1698431365
transform 1 0 7840 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _065_
timestamp 1698431365
transform -1 0 6048 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _066_
timestamp 1698431365
transform -1 0 2464 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _067_
timestamp 1698431365
transform 1 0 5488 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _068_
timestamp 1698431365
transform -1 0 5264 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _069_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 7840 0 -1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _070_
timestamp 1698431365
transform -1 0 8512 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _071_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 12768 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _072_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 7616 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _073_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5824 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _074_
timestamp 1698431365
transform -1 0 7840 0 -1 6272
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _075_
timestamp 1698431365
transform -1 0 9184 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _076_
timestamp 1698431365
transform -1 0 7504 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _077_
timestamp 1698431365
transform -1 0 8288 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _078_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 6496 0 -1 4704
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _079_
timestamp 1698431365
transform 1 0 11424 0 -1 4704
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _080_
timestamp 1698431365
transform 1 0 11312 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _081_
timestamp 1698431365
transform -1 0 9184 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _082_
timestamp 1698431365
transform 1 0 11760 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _083_
timestamp 1698431365
transform 1 0 10080 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _084_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 4816 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _085_
timestamp 1698431365
transform -1 0 5712 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _086_
timestamp 1698431365
transform -1 0 7392 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _087_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13328 0 1 7840
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _088_
timestamp 1698431365
transform 1 0 9632 0 1 9408
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _089_
timestamp 1698431365
transform -1 0 20720 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _090_
timestamp 1698431365
transform -1 0 4928 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__045__I open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 7504 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__046__I
timestamp 1698431365
transform -1 0 8400 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__047__I
timestamp 1698431365
transform -1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__061__A3
timestamp 1698431365
transform -1 0 13776 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__063__A3
timestamp 1698431365
transform 1 0 14224 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__065__A2
timestamp 1698431365
transform 1 0 3920 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__070__A1
timestamp 1698431365
transform 1 0 8736 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__072__B
timestamp 1698431365
transform 1 0 7840 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__075__A1
timestamp 1698431365
transform 1 0 9632 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__076__B
timestamp 1698431365
transform 1 0 7392 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__079__A2
timestamp 1698431365
transform 1 0 15568 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__080__A1
timestamp 1698431365
transform 1 0 14672 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__080__B
timestamp 1698431365
transform 1 0 15120 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__082__A1
timestamp 1698431365
transform 1 0 12880 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__082__B
timestamp 1698431365
transform 1 0 13328 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__089__CLK
timestamp 1698431365
transform 1 0 21392 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__089__D
timestamp 1698431365
transform 1 0 20720 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__090__D
timestamp 1698431365
transform 1 0 3472 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I
timestamp 1698431365
transform -1 0 15456 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1698431365
transform -1 0 37744 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1698431365
transform -1 0 37744 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1698431365
transform -1 0 36624 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1698431365
transform -1 0 4704 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1698431365
transform 1 0 17472 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1698431365
transform -1 0 16912 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input7_I
timestamp 1698431365
transform 1 0 17920 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input8_I
timestamp 1698431365
transform -1 0 18816 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input9_I
timestamp 1698431365
transform -1 0 19600 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input10_I
timestamp 1698431365
transform -1 0 20608 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input11_I
timestamp 1698431365
transform -1 0 21616 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input12_I
timestamp 1698431365
transform -1 0 22064 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input13_I
timestamp 1698431365
transform 1 0 24528 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input14_I
timestamp 1698431365
transform -1 0 24416 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input15_I
timestamp 1698431365
transform -1 0 6496 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input16_I
timestamp 1698431365
transform 1 0 27664 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input17_I
timestamp 1698431365
transform 1 0 26432 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input18_I
timestamp 1698431365
transform 1 0 26880 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input19_I
timestamp 1698431365
transform -1 0 28224 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input20_I
timestamp 1698431365
transform 1 0 29456 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input21_I
timestamp 1698431365
transform 1 0 29904 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input22_I
timestamp 1698431365
transform -1 0 30576 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input23_I
timestamp 1698431365
transform 1 0 31808 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input24_I
timestamp 1698431365
transform 1 0 32480 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input25_I
timestamp 1698431365
transform 1 0 34384 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input26_I
timestamp 1698431365
transform 1 0 8736 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input27_I
timestamp 1698431365
transform -1 0 35056 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input28_I
timestamp 1698431365
transform -1 0 36064 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input29_I
timestamp 1698431365
transform -1 0 7056 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input30_I
timestamp 1698431365
transform -1 0 8512 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input31_I
timestamp 1698431365
transform -1 0 9856 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input32_I
timestamp 1698431365
transform -1 0 3136 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input33_I
timestamp 1698431365
transform -1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input34_I
timestamp 1698431365
transform 1 0 16128 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input35_I
timestamp 1698431365
transform -1 0 15904 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input36_I
timestamp 1698431365
transform -1 0 3136 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input37_I
timestamp 1698431365
transform -1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input38_I
timestamp 1698431365
transform -1 0 6608 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input39_I
timestamp 1698431365
transform 1 0 3360 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input40_I
timestamp 1698431365
transform -1 0 4032 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input41_I
timestamp 1698431365
transform -1 0 37520 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output42_I
timestamp 1698431365
transform -1 0 28000 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output43_I
timestamp 1698431365
transform -1 0 37296 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output47_I
timestamp 1698431365
transform 1 0 2688 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output48_I
timestamp 1698431365
transform 1 0 14784 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 15008 0 -1 6272
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1698431365
transform -1 0 11312 0 1 4704
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1698431365
transform 1 0 10976 0 -1 9408
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_12 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 2688 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_36
timestamp 1698431365
transform 1 0 5376 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_138 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 16800 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_145
timestamp 1698431365
transform 1 0 17584 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_153
timestamp 1698431365
transform 1 0 18480 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_161
timestamp 1698431365
transform 1 0 19376 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_169
timestamp 1698431365
transform 1 0 20272 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_178
timestamp 1698431365
transform 1 0 21280 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_185
timestamp 1698431365
transform 1 0 22064 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_193
timestamp 1698431365
transform 1 0 22960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_201
timestamp 1698431365
transform 1 0 23856 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_203
timestamp 1698431365
transform 1 0 24080 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_218
timestamp 1698431365
transform 1 0 25760 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_225
timestamp 1698431365
transform 1 0 26544 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_233
timestamp 1698431365
transform 1 0 27440 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_237
timestamp 1698431365
transform 1 0 27888 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_258
timestamp 1698431365
transform 1 0 30240 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_265
timestamp 1698431365
transform 1 0 31024 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_314
timestamp 1698431365
transform 1 0 36512 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_321
timestamp 1698431365
transform 1 0 37296 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_329
timestamp 1698431365
transform 1 0 38192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_31
timestamp 1698431365
transform 1 0 4816 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_46
timestamp 1698431365
transform 1 0 6496 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_127
timestamp 1698431365
transform 1 0 15568 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_129
timestamp 1698431365
transform 1 0 15792 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_136
timestamp 1698431365
transform 1 0 16576 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_148
timestamp 1698431365
transform 1 0 17920 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_186
timestamp 1698431365
transform 1 0 22176 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_188
timestamp 1698431365
transform 1 0 22400 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_205
timestamp 1698431365
transform 1 0 24304 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_209
timestamp 1698431365
transform 1 0 24752 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_249
timestamp 1698431365
transform 1 0 29232 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_253
timestamp 1698431365
transform 1 0 29680 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_257
timestamp 1698431365
transform 1 0 30128 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_261 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 30576 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_269
timestamp 1698431365
transform 1 0 31472 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_271
timestamp 1698431365
transform 1 0 31696 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_274 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 32032 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_306
timestamp 1698431365
transform 1 0 35616 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_310
timestamp 1698431365
transform 1 0 36064 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_312
timestamp 1698431365
transform 1 0 36288 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_315
timestamp 1698431365
transform 1 0 36624 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_319
timestamp 1698431365
transform 1 0 37072 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_323
timestamp 1698431365
transform 1 0 37520 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_16
timestamp 1698431365
transform 1 0 3136 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_37
timestamp 1698431365
transform 1 0 5488 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_102
timestamp 1698431365
transform 1 0 12768 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_104
timestamp 1698431365
transform 1 0 12992 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_107
timestamp 1698431365
transform 1 0 13328 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_152
timestamp 1698431365
transform 1 0 18368 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_156
timestamp 1698431365
transform 1 0 18816 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_160
timestamp 1698431365
transform 1 0 19264 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_163
timestamp 1698431365
transform 1 0 19600 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_167
timestamp 1698431365
transform 1 0 20048 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_169
timestamp 1698431365
transform 1 0 20272 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_172
timestamp 1698431365
transform 1 0 20608 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_174
timestamp 1698431365
transform 1 0 20832 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_177
timestamp 1698431365
transform 1 0 21168 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_181
timestamp 1698431365
transform 1 0 21616 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_222
timestamp 1698431365
transform 1 0 26208 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_226
timestamp 1698431365
transform 1 0 26656 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_230
timestamp 1698431365
transform 1 0 27104 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_240
timestamp 1698431365
transform 1 0 28224 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_244
timestamp 1698431365
transform 1 0 28672 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_247
timestamp 1698431365
transform 1 0 29008 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_255
timestamp 1698431365
transform 1 0 29904 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_293
timestamp 1698431365
transform 1 0 34160 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_297
timestamp 1698431365
transform 1 0 34608 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_301
timestamp 1698431365
transform 1 0 35056 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_309
timestamp 1698431365
transform 1 0 35952 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_313
timestamp 1698431365
transform 1 0 36400 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_317
timestamp 1698431365
transform 1 0 36848 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_325
timestamp 1698431365
transform 1 0 37744 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_329
timestamp 1698431365
transform 1 0 38192 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_2
timestamp 1698431365
transform 1 0 1568 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_39
timestamp 1698431365
transform 1 0 5712 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_122
timestamp 1698431365
transform 1 0 15008 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_126
timestamp 1698431365
transform 1 0 15456 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_130
timestamp 1698431365
transform 1 0 15904 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_134
timestamp 1698431365
transform 1 0 16352 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_136
timestamp 1698431365
transform 1 0 16576 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_139
timestamp 1698431365
transform 1 0 16912 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_142
timestamp 1698431365
transform 1 0 17248 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_146
timestamp 1698431365
transform 1 0 17696 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_150 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 18144 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_166
timestamp 1698431365
transform 1 0 19936 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_170
timestamp 1698431365
transform 1 0 20384 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_172
timestamp 1698431365
transform 1 0 20608 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_175
timestamp 1698431365
transform 1 0 20944 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_191
timestamp 1698431365
transform 1 0 22736 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_199
timestamp 1698431365
transform 1 0 23632 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_203
timestamp 1698431365
transform 1 0 24080 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_206
timestamp 1698431365
transform 1 0 24416 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_212 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25088 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_276
timestamp 1698431365
transform 1 0 32256 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_3_282 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 32928 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_314
timestamp 1698431365
transform 1 0 36512 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_330
timestamp 1698431365
transform 1 0 38304 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_2
timestamp 1698431365
transform 1 0 1568 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_32
timestamp 1698431365
transform 1 0 4928 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698431365
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_55
timestamp 1698431365
transform 1 0 7504 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_101
timestamp 1698431365
transform 1 0 12656 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_173
timestamp 1698431365
transform 1 0 20720 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_177
timestamp 1698431365
transform 1 0 21168 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_181
timestamp 1698431365
transform 1 0 21616 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_247
timestamp 1698431365
transform 1 0 29008 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698431365
transform 1 0 36176 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_317
timestamp 1698431365
transform 1 0 36848 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_321
timestamp 1698431365
transform 1 0 37296 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_16
timestamp 1698431365
transform 1 0 3136 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_18
timestamp 1698431365
transform 1 0 3360 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_21
timestamp 1698431365
transform 1 0 3696 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_62
timestamp 1698431365
transform 1 0 8288 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_64
timestamp 1698431365
transform 1 0 8512 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_72
timestamp 1698431365
transform 1 0 9408 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_113
timestamp 1698431365
transform 1 0 14000 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_117
timestamp 1698431365
transform 1 0 14448 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_121
timestamp 1698431365
transform 1 0 14896 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_125
timestamp 1698431365
transform 1 0 15344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_129
timestamp 1698431365
transform 1 0 15792 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_137
timestamp 1698431365
transform 1 0 16688 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_139
timestamp 1698431365
transform 1 0 16912 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_142
timestamp 1698431365
transform 1 0 17248 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_206
timestamp 1698431365
transform 1 0 24416 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_212
timestamp 1698431365
transform 1 0 25088 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_276
timestamp 1698431365
transform 1 0 32256 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_5_282
timestamp 1698431365
transform 1 0 32928 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_314
timestamp 1698431365
transform 1 0 36512 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_330
timestamp 1698431365
transform 1 0 38304 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_6
timestamp 1698431365
transform 1 0 2016 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_16
timestamp 1698431365
transform 1 0 3136 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_20
timestamp 1698431365
transform 1 0 3584 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_24
timestamp 1698431365
transform 1 0 4032 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_30
timestamp 1698431365
transform 1 0 4704 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_32
timestamp 1698431365
transform 1 0 4928 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_42
timestamp 1698431365
transform 1 0 6048 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_44
timestamp 1698431365
transform 1 0 6272 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_47
timestamp 1698431365
transform 1 0 6608 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_51
timestamp 1698431365
transform 1 0 7056 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_64
timestamp 1698431365
transform 1 0 8512 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_138
timestamp 1698431365
transform 1 0 16800 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_170
timestamp 1698431365
transform 1 0 20384 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_174
timestamp 1698431365
transform 1 0 20832 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_177
timestamp 1698431365
transform 1 0 21168 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_241
timestamp 1698431365
transform 1 0 28336 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_247
timestamp 1698431365
transform 1 0 29008 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_311
timestamp 1698431365
transform 1 0 36176 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_317
timestamp 1698431365
transform 1 0 36848 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_325
timestamp 1698431365
transform 1 0 37744 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_329
timestamp 1698431365
transform 1 0 38192 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_7_2
timestamp 1698431365
transform 1 0 1568 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_34
timestamp 1698431365
transform 1 0 5152 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_42
timestamp 1698431365
transform 1 0 6048 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_46
timestamp 1698431365
transform 1 0 6496 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_56
timestamp 1698431365
transform 1 0 7616 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_60
timestamp 1698431365
transform 1 0 8064 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_64
timestamp 1698431365
transform 1 0 8512 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_68
timestamp 1698431365
transform 1 0 8960 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_72
timestamp 1698431365
transform 1 0 9408 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_76
timestamp 1698431365
transform 1 0 9856 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_136
timestamp 1698431365
transform 1 0 16576 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_142
timestamp 1698431365
transform 1 0 17248 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_206
timestamp 1698431365
transform 1 0 24416 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_212
timestamp 1698431365
transform 1 0 25088 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_276
timestamp 1698431365
transform 1 0 32256 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_7_282
timestamp 1698431365
transform 1 0 32928 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_314
timestamp 1698431365
transform 1 0 36512 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_330
timestamp 1698431365
transform 1 0 38304 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_6
timestamp 1698431365
transform 1 0 2016 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_22
timestamp 1698431365
transform 1 0 3808 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_30
timestamp 1698431365
transform 1 0 4704 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698431365
transform 1 0 5152 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_37
timestamp 1698431365
transform 1 0 5488 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_53
timestamp 1698431365
transform 1 0 7280 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_59
timestamp 1698431365
transform 1 0 7952 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_63
timestamp 1698431365
transform 1 0 8400 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_71
timestamp 1698431365
transform 1 0 9296 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_73
timestamp 1698431365
transform 1 0 9520 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_107
timestamp 1698431365
transform 1 0 13328 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_111
timestamp 1698431365
transform 1 0 13776 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_177
timestamp 1698431365
transform 1 0 21168 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_241
timestamp 1698431365
transform 1 0 28336 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_247
timestamp 1698431365
transform 1 0 29008 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_311
timestamp 1698431365
transform 1 0 36176 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_317
timestamp 1698431365
transform 1 0 36848 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_325
timestamp 1698431365
transform 1 0 37744 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_329
timestamp 1698431365
transform 1 0 38192 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2
timestamp 1698431365
transform 1 0 1568 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698431365
transform 1 0 8736 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_72
timestamp 1698431365
transform 1 0 9408 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_88
timestamp 1698431365
transform 1 0 11200 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_92
timestamp 1698431365
transform 1 0 11648 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_101
timestamp 1698431365
transform 1 0 12656 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_105
timestamp 1698431365
transform 1 0 13104 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_109
timestamp 1698431365
transform 1 0 13552 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_125
timestamp 1698431365
transform 1 0 15344 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_133
timestamp 1698431365
transform 1 0 16240 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_137
timestamp 1698431365
transform 1 0 16688 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_139
timestamp 1698431365
transform 1 0 16912 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_142
timestamp 1698431365
transform 1 0 17248 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_206
timestamp 1698431365
transform 1 0 24416 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_212
timestamp 1698431365
transform 1 0 25088 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_276
timestamp 1698431365
transform 1 0 32256 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_9_282
timestamp 1698431365
transform 1 0 32928 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_314
timestamp 1698431365
transform 1 0 36512 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_330
timestamp 1698431365
transform 1 0 38304 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_6
timestamp 1698431365
transform 1 0 2016 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_22
timestamp 1698431365
transform 1 0 3808 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_30
timestamp 1698431365
transform 1 0 4704 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698431365
transform 1 0 5152 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_37
timestamp 1698431365
transform 1 0 5488 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698431365
transform 1 0 12656 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_107
timestamp 1698431365
transform 1 0 13328 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_171
timestamp 1698431365
transform 1 0 20496 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_177
timestamp 1698431365
transform 1 0 21168 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_241
timestamp 1698431365
transform 1 0 28336 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_247
timestamp 1698431365
transform 1 0 29008 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_311
timestamp 1698431365
transform 1 0 36176 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_317
timestamp 1698431365
transform 1 0 36848 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_325
timestamp 1698431365
transform 1 0 37744 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_329
timestamp 1698431365
transform 1 0 38192 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2
timestamp 1698431365
transform 1 0 1568 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_66
timestamp 1698431365
transform 1 0 8736 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_72
timestamp 1698431365
transform 1 0 9408 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_136
timestamp 1698431365
transform 1 0 16576 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_142
timestamp 1698431365
transform 1 0 17248 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_206
timestamp 1698431365
transform 1 0 24416 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_212
timestamp 1698431365
transform 1 0 25088 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_276
timestamp 1698431365
transform 1 0 32256 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_11_282
timestamp 1698431365
transform 1 0 32928 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_314
timestamp 1698431365
transform 1 0 36512 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_330
timestamp 1698431365
transform 1 0 38304 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_6
timestamp 1698431365
transform 1 0 2016 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_22
timestamp 1698431365
transform 1 0 3808 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_30
timestamp 1698431365
transform 1 0 4704 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698431365
transform 1 0 5152 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_37
timestamp 1698431365
transform 1 0 5488 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_101
timestamp 1698431365
transform 1 0 12656 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_107
timestamp 1698431365
transform 1 0 13328 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_171
timestamp 1698431365
transform 1 0 20496 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_177
timestamp 1698431365
transform 1 0 21168 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_241
timestamp 1698431365
transform 1 0 28336 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_247
timestamp 1698431365
transform 1 0 29008 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_311
timestamp 1698431365
transform 1 0 36176 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_317
timestamp 1698431365
transform 1 0 36848 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_325
timestamp 1698431365
transform 1 0 37744 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_329
timestamp 1698431365
transform 1 0 38192 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_6
timestamp 1698431365
transform 1 0 2016 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_72
timestamp 1698431365
transform 1 0 9408 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_136
timestamp 1698431365
transform 1 0 16576 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_142
timestamp 1698431365
transform 1 0 17248 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_206
timestamp 1698431365
transform 1 0 24416 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_212
timestamp 1698431365
transform 1 0 25088 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_276
timestamp 1698431365
transform 1 0 32256 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_282
timestamp 1698431365
transform 1 0 32928 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_314
timestamp 1698431365
transform 1 0 36512 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_330
timestamp 1698431365
transform 1 0 38304 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_2
timestamp 1698431365
transform 1 0 1568 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698431365
transform 1 0 5152 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_37
timestamp 1698431365
transform 1 0 5488 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_101
timestamp 1698431365
transform 1 0 12656 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_107
timestamp 1698431365
transform 1 0 13328 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_171
timestamp 1698431365
transform 1 0 20496 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_177
timestamp 1698431365
transform 1 0 21168 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_241
timestamp 1698431365
transform 1 0 28336 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_247
timestamp 1698431365
transform 1 0 29008 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_311
timestamp 1698431365
transform 1 0 36176 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_317
timestamp 1698431365
transform 1 0 36848 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_325
timestamp 1698431365
transform 1 0 37744 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_329
timestamp 1698431365
transform 1 0 38192 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_6
timestamp 1698431365
transform 1 0 2016 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_72
timestamp 1698431365
transform 1 0 9408 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_136
timestamp 1698431365
transform 1 0 16576 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_142
timestamp 1698431365
transform 1 0 17248 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_206
timestamp 1698431365
transform 1 0 24416 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_212
timestamp 1698431365
transform 1 0 25088 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_276
timestamp 1698431365
transform 1 0 32256 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_282
timestamp 1698431365
transform 1 0 32928 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_314
timestamp 1698431365
transform 1 0 36512 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_330
timestamp 1698431365
transform 1 0 38304 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_2
timestamp 1698431365
transform 1 0 1568 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698431365
transform 1 0 5152 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_37
timestamp 1698431365
transform 1 0 5488 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_101
timestamp 1698431365
transform 1 0 12656 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_107
timestamp 1698431365
transform 1 0 13328 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_171
timestamp 1698431365
transform 1 0 20496 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_177
timestamp 1698431365
transform 1 0 21168 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_241
timestamp 1698431365
transform 1 0 28336 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_247
timestamp 1698431365
transform 1 0 29008 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_311
timestamp 1698431365
transform 1 0 36176 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_317
timestamp 1698431365
transform 1 0 36848 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_325
timestamp 1698431365
transform 1 0 37744 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_329
timestamp 1698431365
transform 1 0 38192 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_6
timestamp 1698431365
transform 1 0 2016 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_72
timestamp 1698431365
transform 1 0 9408 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_136
timestamp 1698431365
transform 1 0 16576 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_142
timestamp 1698431365
transform 1 0 17248 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_206
timestamp 1698431365
transform 1 0 24416 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_212
timestamp 1698431365
transform 1 0 25088 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_276
timestamp 1698431365
transform 1 0 32256 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_282
timestamp 1698431365
transform 1 0 32928 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_314
timestamp 1698431365
transform 1 0 36512 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_330
timestamp 1698431365
transform 1 0 38304 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_6
timestamp 1698431365
transform 1 0 2016 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_22
timestamp 1698431365
transform 1 0 3808 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_30
timestamp 1698431365
transform 1 0 4704 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698431365
transform 1 0 5152 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_37
timestamp 1698431365
transform 1 0 5488 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_101
timestamp 1698431365
transform 1 0 12656 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_107
timestamp 1698431365
transform 1 0 13328 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_171
timestamp 1698431365
transform 1 0 20496 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_177
timestamp 1698431365
transform 1 0 21168 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_241
timestamp 1698431365
transform 1 0 28336 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_247
timestamp 1698431365
transform 1 0 29008 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_311
timestamp 1698431365
transform 1 0 36176 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_317
timestamp 1698431365
transform 1 0 36848 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_325
timestamp 1698431365
transform 1 0 37744 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_329
timestamp 1698431365
transform 1 0 38192 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_2
timestamp 1698431365
transform 1 0 1568 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_66
timestamp 1698431365
transform 1 0 8736 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_72
timestamp 1698431365
transform 1 0 9408 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_136
timestamp 1698431365
transform 1 0 16576 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_142
timestamp 1698431365
transform 1 0 17248 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_206
timestamp 1698431365
transform 1 0 24416 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_212
timestamp 1698431365
transform 1 0 25088 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_276
timestamp 1698431365
transform 1 0 32256 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_282
timestamp 1698431365
transform 1 0 32928 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_314
timestamp 1698431365
transform 1 0 36512 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_330
timestamp 1698431365
transform 1 0 38304 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_6
timestamp 1698431365
transform 1 0 2016 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_22
timestamp 1698431365
transform 1 0 3808 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_30
timestamp 1698431365
transform 1 0 4704 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698431365
transform 1 0 5152 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_37
timestamp 1698431365
transform 1 0 5488 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_101
timestamp 1698431365
transform 1 0 12656 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_107
timestamp 1698431365
transform 1 0 13328 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_171
timestamp 1698431365
transform 1 0 20496 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_177
timestamp 1698431365
transform 1 0 21168 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_241
timestamp 1698431365
transform 1 0 28336 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_247
timestamp 1698431365
transform 1 0 29008 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_311
timestamp 1698431365
transform 1 0 36176 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_317
timestamp 1698431365
transform 1 0 36848 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_325
timestamp 1698431365
transform 1 0 37744 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_2
timestamp 1698431365
transform 1 0 1568 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_66
timestamp 1698431365
transform 1 0 8736 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_72
timestamp 1698431365
transform 1 0 9408 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_136
timestamp 1698431365
transform 1 0 16576 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_142
timestamp 1698431365
transform 1 0 17248 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_206
timestamp 1698431365
transform 1 0 24416 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_212
timestamp 1698431365
transform 1 0 25088 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_276
timestamp 1698431365
transform 1 0 32256 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_282
timestamp 1698431365
transform 1 0 32928 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_314
timestamp 1698431365
transform 1 0 36512 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_330
timestamp 1698431365
transform 1 0 38304 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_6
timestamp 1698431365
transform 1 0 2016 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_22
timestamp 1698431365
transform 1 0 3808 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_30
timestamp 1698431365
transform 1 0 4704 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698431365
transform 1 0 5152 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_37
timestamp 1698431365
transform 1 0 5488 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_101
timestamp 1698431365
transform 1 0 12656 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_107
timestamp 1698431365
transform 1 0 13328 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_171
timestamp 1698431365
transform 1 0 20496 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_177
timestamp 1698431365
transform 1 0 21168 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_241
timestamp 1698431365
transform 1 0 28336 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_247
timestamp 1698431365
transform 1 0 29008 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_311
timestamp 1698431365
transform 1 0 36176 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_317
timestamp 1698431365
transform 1 0 36848 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_325
timestamp 1698431365
transform 1 0 37744 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_329
timestamp 1698431365
transform 1 0 38192 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_2
timestamp 1698431365
transform 1 0 1568 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_66
timestamp 1698431365
transform 1 0 8736 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_72
timestamp 1698431365
transform 1 0 9408 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_136
timestamp 1698431365
transform 1 0 16576 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_142
timestamp 1698431365
transform 1 0 17248 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_206
timestamp 1698431365
transform 1 0 24416 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_212
timestamp 1698431365
transform 1 0 25088 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_276
timestamp 1698431365
transform 1 0 32256 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_282
timestamp 1698431365
transform 1 0 32928 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_314
timestamp 1698431365
transform 1 0 36512 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_330
timestamp 1698431365
transform 1 0 38304 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_6
timestamp 1698431365
transform 1 0 2016 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_22
timestamp 1698431365
transform 1 0 3808 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_30
timestamp 1698431365
transform 1 0 4704 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698431365
transform 1 0 5152 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_37
timestamp 1698431365
transform 1 0 5488 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_101
timestamp 1698431365
transform 1 0 12656 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_107
timestamp 1698431365
transform 1 0 13328 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_171
timestamp 1698431365
transform 1 0 20496 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_177
timestamp 1698431365
transform 1 0 21168 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_241
timestamp 1698431365
transform 1 0 28336 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_247
timestamp 1698431365
transform 1 0 29008 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_311
timestamp 1698431365
transform 1 0 36176 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_317
timestamp 1698431365
transform 1 0 36848 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_325
timestamp 1698431365
transform 1 0 37744 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_329
timestamp 1698431365
transform 1 0 38192 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_6
timestamp 1698431365
transform 1 0 2016 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_72
timestamp 1698431365
transform 1 0 9408 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_136
timestamp 1698431365
transform 1 0 16576 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_142
timestamp 1698431365
transform 1 0 17248 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_206
timestamp 1698431365
transform 1 0 24416 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_212
timestamp 1698431365
transform 1 0 25088 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_276
timestamp 1698431365
transform 1 0 32256 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_282
timestamp 1698431365
transform 1 0 32928 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_314
timestamp 1698431365
transform 1 0 36512 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_330
timestamp 1698431365
transform 1 0 38304 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_2
timestamp 1698431365
transform 1 0 1568 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698431365
transform 1 0 5152 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_37
timestamp 1698431365
transform 1 0 5488 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_101
timestamp 1698431365
transform 1 0 12656 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_107
timestamp 1698431365
transform 1 0 13328 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_171
timestamp 1698431365
transform 1 0 20496 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_177
timestamp 1698431365
transform 1 0 21168 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_241
timestamp 1698431365
transform 1 0 28336 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_247
timestamp 1698431365
transform 1 0 29008 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_311
timestamp 1698431365
transform 1 0 36176 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_317
timestamp 1698431365
transform 1 0 36848 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_325
timestamp 1698431365
transform 1 0 37744 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_329
timestamp 1698431365
transform 1 0 38192 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_6
timestamp 1698431365
transform 1 0 2016 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_72
timestamp 1698431365
transform 1 0 9408 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_136
timestamp 1698431365
transform 1 0 16576 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_142
timestamp 1698431365
transform 1 0 17248 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_206
timestamp 1698431365
transform 1 0 24416 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_212
timestamp 1698431365
transform 1 0 25088 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_276
timestamp 1698431365
transform 1 0 32256 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_282
timestamp 1698431365
transform 1 0 32928 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_314
timestamp 1698431365
transform 1 0 36512 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_330
timestamp 1698431365
transform 1 0 38304 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_2
timestamp 1698431365
transform 1 0 1568 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698431365
transform 1 0 5152 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_37
timestamp 1698431365
transform 1 0 5488 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_101
timestamp 1698431365
transform 1 0 12656 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_107
timestamp 1698431365
transform 1 0 13328 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_171
timestamp 1698431365
transform 1 0 20496 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_177
timestamp 1698431365
transform 1 0 21168 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_241
timestamp 1698431365
transform 1 0 28336 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_247
timestamp 1698431365
transform 1 0 29008 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_311
timestamp 1698431365
transform 1 0 36176 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_317
timestamp 1698431365
transform 1 0 36848 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_325
timestamp 1698431365
transform 1 0 37744 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_329
timestamp 1698431365
transform 1 0 38192 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_6
timestamp 1698431365
transform 1 0 2016 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_72
timestamp 1698431365
transform 1 0 9408 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_136
timestamp 1698431365
transform 1 0 16576 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_142
timestamp 1698431365
transform 1 0 17248 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_206
timestamp 1698431365
transform 1 0 24416 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_212
timestamp 1698431365
transform 1 0 25088 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_276
timestamp 1698431365
transform 1 0 32256 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_282
timestamp 1698431365
transform 1 0 32928 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_314
timestamp 1698431365
transform 1 0 36512 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_330
timestamp 1698431365
transform 1 0 38304 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_6
timestamp 1698431365
transform 1 0 2016 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_22
timestamp 1698431365
transform 1 0 3808 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_30
timestamp 1698431365
transform 1 0 4704 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698431365
transform 1 0 5152 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_37
timestamp 1698431365
transform 1 0 5488 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_101
timestamp 1698431365
transform 1 0 12656 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_107
timestamp 1698431365
transform 1 0 13328 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_171
timestamp 1698431365
transform 1 0 20496 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_177
timestamp 1698431365
transform 1 0 21168 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_241
timestamp 1698431365
transform 1 0 28336 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_247
timestamp 1698431365
transform 1 0 29008 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_311
timestamp 1698431365
transform 1 0 36176 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_317
timestamp 1698431365
transform 1 0 36848 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_325
timestamp 1698431365
transform 1 0 37744 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_329
timestamp 1698431365
transform 1 0 38192 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_2
timestamp 1698431365
transform 1 0 1568 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_66
timestamp 1698431365
transform 1 0 8736 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_72
timestamp 1698431365
transform 1 0 9408 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_136
timestamp 1698431365
transform 1 0 16576 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_142
timestamp 1698431365
transform 1 0 17248 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_206
timestamp 1698431365
transform 1 0 24416 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_212
timestamp 1698431365
transform 1 0 25088 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_276
timestamp 1698431365
transform 1 0 32256 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_282
timestamp 1698431365
transform 1 0 32928 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_314
timestamp 1698431365
transform 1 0 36512 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_330
timestamp 1698431365
transform 1 0 38304 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_6
timestamp 1698431365
transform 1 0 2016 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_22
timestamp 1698431365
transform 1 0 3808 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_30
timestamp 1698431365
transform 1 0 4704 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698431365
transform 1 0 5152 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_37
timestamp 1698431365
transform 1 0 5488 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_101
timestamp 1698431365
transform 1 0 12656 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_107
timestamp 1698431365
transform 1 0 13328 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_171
timestamp 1698431365
transform 1 0 20496 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_177
timestamp 1698431365
transform 1 0 21168 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_241
timestamp 1698431365
transform 1 0 28336 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_247
timestamp 1698431365
transform 1 0 29008 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_311
timestamp 1698431365
transform 1 0 36176 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_317
timestamp 1698431365
transform 1 0 36848 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_325
timestamp 1698431365
transform 1 0 37744 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_329
timestamp 1698431365
transform 1 0 38192 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_2
timestamp 1698431365
transform 1 0 1568 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_66
timestamp 1698431365
transform 1 0 8736 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_72
timestamp 1698431365
transform 1 0 9408 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_136
timestamp 1698431365
transform 1 0 16576 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_142
timestamp 1698431365
transform 1 0 17248 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_206
timestamp 1698431365
transform 1 0 24416 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_212
timestamp 1698431365
transform 1 0 25088 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_276
timestamp 1698431365
transform 1 0 32256 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_33_282
timestamp 1698431365
transform 1 0 32928 0 -1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_314
timestamp 1698431365
transform 1 0 36512 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_330
timestamp 1698431365
transform 1 0 38304 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_6
timestamp 1698431365
transform 1 0 2016 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_22
timestamp 1698431365
transform 1 0 3808 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_30
timestamp 1698431365
transform 1 0 4704 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698431365
transform 1 0 5152 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_37
timestamp 1698431365
transform 1 0 5488 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_101
timestamp 1698431365
transform 1 0 12656 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_107
timestamp 1698431365
transform 1 0 13328 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_171
timestamp 1698431365
transform 1 0 20496 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_177
timestamp 1698431365
transform 1 0 21168 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_241
timestamp 1698431365
transform 1 0 28336 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_247
timestamp 1698431365
transform 1 0 29008 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_311
timestamp 1698431365
transform 1 0 36176 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_317
timestamp 1698431365
transform 1 0 36848 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_325
timestamp 1698431365
transform 1 0 37744 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_329
timestamp 1698431365
transform 1 0 38192 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_2
timestamp 1698431365
transform 1 0 1568 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_66
timestamp 1698431365
transform 1 0 8736 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_72
timestamp 1698431365
transform 1 0 9408 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_136
timestamp 1698431365
transform 1 0 16576 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_142
timestamp 1698431365
transform 1 0 17248 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_206
timestamp 1698431365
transform 1 0 24416 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_212
timestamp 1698431365
transform 1 0 25088 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_276
timestamp 1698431365
transform 1 0 32256 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_35_282
timestamp 1698431365
transform 1 0 32928 0 -1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_314
timestamp 1698431365
transform 1 0 36512 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_330
timestamp 1698431365
transform 1 0 38304 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_6
timestamp 1698431365
transform 1 0 2016 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_22
timestamp 1698431365
transform 1 0 3808 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_30
timestamp 1698431365
transform 1 0 4704 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698431365
transform 1 0 5152 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_37
timestamp 1698431365
transform 1 0 5488 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_101
timestamp 1698431365
transform 1 0 12656 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_107
timestamp 1698431365
transform 1 0 13328 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_171
timestamp 1698431365
transform 1 0 20496 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_177
timestamp 1698431365
transform 1 0 21168 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_241
timestamp 1698431365
transform 1 0 28336 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_247
timestamp 1698431365
transform 1 0 29008 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_311
timestamp 1698431365
transform 1 0 36176 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_317
timestamp 1698431365
transform 1 0 36848 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_321
timestamp 1698431365
transform 1 0 37296 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_6
timestamp 1698431365
transform 1 0 2016 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_72
timestamp 1698431365
transform 1 0 9408 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_136
timestamp 1698431365
transform 1 0 16576 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_142
timestamp 1698431365
transform 1 0 17248 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_206
timestamp 1698431365
transform 1 0 24416 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_212
timestamp 1698431365
transform 1 0 25088 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_276
timestamp 1698431365
transform 1 0 32256 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_37_282
timestamp 1698431365
transform 1 0 32928 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_314
timestamp 1698431365
transform 1 0 36512 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_330
timestamp 1698431365
transform 1 0 38304 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_2
timestamp 1698431365
transform 1 0 1568 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698431365
transform 1 0 5152 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_37
timestamp 1698431365
transform 1 0 5488 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_101
timestamp 1698431365
transform 1 0 12656 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_107
timestamp 1698431365
transform 1 0 13328 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_171
timestamp 1698431365
transform 1 0 20496 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_177
timestamp 1698431365
transform 1 0 21168 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_241
timestamp 1698431365
transform 1 0 28336 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_247
timestamp 1698431365
transform 1 0 29008 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_311
timestamp 1698431365
transform 1 0 36176 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_317
timestamp 1698431365
transform 1 0 36848 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_325
timestamp 1698431365
transform 1 0 37744 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_329
timestamp 1698431365
transform 1 0 38192 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_6
timestamp 1698431365
transform 1 0 2016 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_72
timestamp 1698431365
transform 1 0 9408 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_136
timestamp 1698431365
transform 1 0 16576 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_142
timestamp 1698431365
transform 1 0 17248 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_206
timestamp 1698431365
transform 1 0 24416 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_212
timestamp 1698431365
transform 1 0 25088 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_276
timestamp 1698431365
transform 1 0 32256 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_39_282
timestamp 1698431365
transform 1 0 32928 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_314
timestamp 1698431365
transform 1 0 36512 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_330
timestamp 1698431365
transform 1 0 38304 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_2
timestamp 1698431365
transform 1 0 1568 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698431365
transform 1 0 5152 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_37
timestamp 1698431365
transform 1 0 5488 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_101
timestamp 1698431365
transform 1 0 12656 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_107
timestamp 1698431365
transform 1 0 13328 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_171
timestamp 1698431365
transform 1 0 20496 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_177
timestamp 1698431365
transform 1 0 21168 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_241
timestamp 1698431365
transform 1 0 28336 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_247
timestamp 1698431365
transform 1 0 29008 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_311
timestamp 1698431365
transform 1 0 36176 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_317
timestamp 1698431365
transform 1 0 36848 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_325
timestamp 1698431365
transform 1 0 37744 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_329
timestamp 1698431365
transform 1 0 38192 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_6
timestamp 1698431365
transform 1 0 2016 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_72
timestamp 1698431365
transform 1 0 9408 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_136
timestamp 1698431365
transform 1 0 16576 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_142
timestamp 1698431365
transform 1 0 17248 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_206
timestamp 1698431365
transform 1 0 24416 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_212
timestamp 1698431365
transform 1 0 25088 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_276
timestamp 1698431365
transform 1 0 32256 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_41_282
timestamp 1698431365
transform 1 0 32928 0 -1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_314
timestamp 1698431365
transform 1 0 36512 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_330
timestamp 1698431365
transform 1 0 38304 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_6
timestamp 1698431365
transform 1 0 2016 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_22
timestamp 1698431365
transform 1 0 3808 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_30
timestamp 1698431365
transform 1 0 4704 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698431365
transform 1 0 5152 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_37
timestamp 1698431365
transform 1 0 5488 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_101
timestamp 1698431365
transform 1 0 12656 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_107
timestamp 1698431365
transform 1 0 13328 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_171
timestamp 1698431365
transform 1 0 20496 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_177
timestamp 1698431365
transform 1 0 21168 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_241
timestamp 1698431365
transform 1 0 28336 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_247
timestamp 1698431365
transform 1 0 29008 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_311
timestamp 1698431365
transform 1 0 36176 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_317
timestamp 1698431365
transform 1 0 36848 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_325
timestamp 1698431365
transform 1 0 37744 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_329
timestamp 1698431365
transform 1 0 38192 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_2
timestamp 1698431365
transform 1 0 1568 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_66
timestamp 1698431365
transform 1 0 8736 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_72
timestamp 1698431365
transform 1 0 9408 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_136
timestamp 1698431365
transform 1 0 16576 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_142
timestamp 1698431365
transform 1 0 17248 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_206
timestamp 1698431365
transform 1 0 24416 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_212
timestamp 1698431365
transform 1 0 25088 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_276
timestamp 1698431365
transform 1 0 32256 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_282
timestamp 1698431365
transform 1 0 32928 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_314
timestamp 1698431365
transform 1 0 36512 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_330
timestamp 1698431365
transform 1 0 38304 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_6
timestamp 1698431365
transform 1 0 2016 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_22
timestamp 1698431365
transform 1 0 3808 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_30
timestamp 1698431365
transform 1 0 4704 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_34
timestamp 1698431365
transform 1 0 5152 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_37
timestamp 1698431365
transform 1 0 5488 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_101
timestamp 1698431365
transform 1 0 12656 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_107
timestamp 1698431365
transform 1 0 13328 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_171
timestamp 1698431365
transform 1 0 20496 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_177
timestamp 1698431365
transform 1 0 21168 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_241
timestamp 1698431365
transform 1 0 28336 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_247
timestamp 1698431365
transform 1 0 29008 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_311
timestamp 1698431365
transform 1 0 36176 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_317
timestamp 1698431365
transform 1 0 36848 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_325
timestamp 1698431365
transform 1 0 37744 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_329
timestamp 1698431365
transform 1 0 38192 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_2
timestamp 1698431365
transform 1 0 1568 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_66
timestamp 1698431365
transform 1 0 8736 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_72
timestamp 1698431365
transform 1 0 9408 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_136
timestamp 1698431365
transform 1 0 16576 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_142
timestamp 1698431365
transform 1 0 17248 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_206
timestamp 1698431365
transform 1 0 24416 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_212
timestamp 1698431365
transform 1 0 25088 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_276
timestamp 1698431365
transform 1 0 32256 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_45_282
timestamp 1698431365
transform 1 0 32928 0 -1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_314
timestamp 1698431365
transform 1 0 36512 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_330
timestamp 1698431365
transform 1 0 38304 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_6
timestamp 1698431365
transform 1 0 2016 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_22
timestamp 1698431365
transform 1 0 3808 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_30
timestamp 1698431365
transform 1 0 4704 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_34
timestamp 1698431365
transform 1 0 5152 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_37
timestamp 1698431365
transform 1 0 5488 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_101
timestamp 1698431365
transform 1 0 12656 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_107
timestamp 1698431365
transform 1 0 13328 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_171
timestamp 1698431365
transform 1 0 20496 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_177
timestamp 1698431365
transform 1 0 21168 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_241
timestamp 1698431365
transform 1 0 28336 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_247
timestamp 1698431365
transform 1 0 29008 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_311
timestamp 1698431365
transform 1 0 36176 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_317
timestamp 1698431365
transform 1 0 36848 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_325
timestamp 1698431365
transform 1 0 37744 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_329
timestamp 1698431365
transform 1 0 38192 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_2
timestamp 1698431365
transform 1 0 1568 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_66
timestamp 1698431365
transform 1 0 8736 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_72
timestamp 1698431365
transform 1 0 9408 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_136
timestamp 1698431365
transform 1 0 16576 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_142
timestamp 1698431365
transform 1 0 17248 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_206
timestamp 1698431365
transform 1 0 24416 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_212
timestamp 1698431365
transform 1 0 25088 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_276
timestamp 1698431365
transform 1 0 32256 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_47_282
timestamp 1698431365
transform 1 0 32928 0 -1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_314
timestamp 1698431365
transform 1 0 36512 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_330
timestamp 1698431365
transform 1 0 38304 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_48_6
timestamp 1698431365
transform 1 0 2016 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_22
timestamp 1698431365
transform 1 0 3808 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_30
timestamp 1698431365
transform 1 0 4704 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_34
timestamp 1698431365
transform 1 0 5152 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_37
timestamp 1698431365
transform 1 0 5488 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_101
timestamp 1698431365
transform 1 0 12656 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_107
timestamp 1698431365
transform 1 0 13328 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_171
timestamp 1698431365
transform 1 0 20496 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_177
timestamp 1698431365
transform 1 0 21168 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_241
timestamp 1698431365
transform 1 0 28336 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_247
timestamp 1698431365
transform 1 0 29008 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_311
timestamp 1698431365
transform 1 0 36176 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_317
timestamp 1698431365
transform 1 0 36848 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_325
timestamp 1698431365
transform 1 0 37744 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_329
timestamp 1698431365
transform 1 0 38192 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_6
timestamp 1698431365
transform 1 0 2016 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_72
timestamp 1698431365
transform 1 0 9408 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_136
timestamp 1698431365
transform 1 0 16576 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_142
timestamp 1698431365
transform 1 0 17248 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_206
timestamp 1698431365
transform 1 0 24416 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_212
timestamp 1698431365
transform 1 0 25088 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_276
timestamp 1698431365
transform 1 0 32256 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_49_282
timestamp 1698431365
transform 1 0 32928 0 -1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_314
timestamp 1698431365
transform 1 0 36512 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_330
timestamp 1698431365
transform 1 0 38304 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_50_2
timestamp 1698431365
transform 1 0 1568 0 1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_34
timestamp 1698431365
transform 1 0 5152 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_37
timestamp 1698431365
transform 1 0 5488 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_101
timestamp 1698431365
transform 1 0 12656 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_107
timestamp 1698431365
transform 1 0 13328 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_171
timestamp 1698431365
transform 1 0 20496 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_177
timestamp 1698431365
transform 1 0 21168 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_241
timestamp 1698431365
transform 1 0 28336 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_247
timestamp 1698431365
transform 1 0 29008 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_311
timestamp 1698431365
transform 1 0 36176 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_317
timestamp 1698431365
transform 1 0 36848 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_325
timestamp 1698431365
transform 1 0 37744 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_329
timestamp 1698431365
transform 1 0 38192 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_6
timestamp 1698431365
transform 1 0 2016 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_72
timestamp 1698431365
transform 1 0 9408 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_136
timestamp 1698431365
transform 1 0 16576 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_142
timestamp 1698431365
transform 1 0 17248 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_206
timestamp 1698431365
transform 1 0 24416 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_212
timestamp 1698431365
transform 1 0 25088 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_276
timestamp 1698431365
transform 1 0 32256 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_51_282
timestamp 1698431365
transform 1 0 32928 0 -1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_314
timestamp 1698431365
transform 1 0 36512 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_322
timestamp 1698431365
transform 1 0 37408 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_326
timestamp 1698431365
transform 1 0 37856 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_52_2
timestamp 1698431365
transform 1 0 1568 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_34
timestamp 1698431365
transform 1 0 5152 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_37
timestamp 1698431365
transform 1 0 5488 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_101
timestamp 1698431365
transform 1 0 12656 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_107
timestamp 1698431365
transform 1 0 13328 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_171
timestamp 1698431365
transform 1 0 20496 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_177
timestamp 1698431365
transform 1 0 21168 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_241
timestamp 1698431365
transform 1 0 28336 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_247
timestamp 1698431365
transform 1 0 29008 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_311
timestamp 1698431365
transform 1 0 36176 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_317
timestamp 1698431365
transform 1 0 36848 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_325
timestamp 1698431365
transform 1 0 37744 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_329
timestamp 1698431365
transform 1 0 38192 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_10
timestamp 1698431365
transform 1 0 2464 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_53_14
timestamp 1698431365
transform 1 0 2912 0 -1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_53_46
timestamp 1698431365
transform 1 0 6496 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_62
timestamp 1698431365
transform 1 0 8288 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_72
timestamp 1698431365
transform 1 0 9408 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_136
timestamp 1698431365
transform 1 0 16576 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_142
timestamp 1698431365
transform 1 0 17248 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_206
timestamp 1698431365
transform 1 0 24416 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_212
timestamp 1698431365
transform 1 0 25088 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_276
timestamp 1698431365
transform 1 0 32256 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_53_282
timestamp 1698431365
transform 1 0 32928 0 -1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_53_314
timestamp 1698431365
transform 1 0 36512 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_330
timestamp 1698431365
transform 1 0 38304 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_2
timestamp 1698431365
transform 1 0 1568 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_4
timestamp 1698431365
transform 1 0 1792 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_23
timestamp 1698431365
transform 1 0 3920 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_31
timestamp 1698431365
transform 1 0 4816 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_33
timestamp 1698431365
transform 1 0 5040 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_36
timestamp 1698431365
transform 1 0 5376 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_52
timestamp 1698431365
transform 1 0 7168 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_56
timestamp 1698431365
transform 1 0 7616 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_61
timestamp 1698431365
transform 1 0 8176 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_65
timestamp 1698431365
transform 1 0 8624 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_67
timestamp 1698431365
transform 1 0 8848 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_54_70
timestamp 1698431365
transform 1 0 9184 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_118
timestamp 1698431365
transform 1 0 14560 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_122
timestamp 1698431365
transform 1 0 15008 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_130
timestamp 1698431365
transform 1 0 15904 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_134
timestamp 1698431365
transform 1 0 16352 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_138
timestamp 1698431365
transform 1 0 16800 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_142
timestamp 1698431365
transform 1 0 17248 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_144
timestamp 1698431365
transform 1 0 17472 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_149
timestamp 1698431365
transform 1 0 18032 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_165
timestamp 1698431365
transform 1 0 19824 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_169
timestamp 1698431365
transform 1 0 20272 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_172
timestamp 1698431365
transform 1 0 20608 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_188
timestamp 1698431365
transform 1 0 22400 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_193
timestamp 1698431365
transform 1 0 22960 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_201
timestamp 1698431365
transform 1 0 23856 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_203
timestamp 1698431365
transform 1 0 24080 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_206
timestamp 1698431365
transform 1 0 24416 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_222
timestamp 1698431365
transform 1 0 26208 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_230
timestamp 1698431365
transform 1 0 27104 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_234
timestamp 1698431365
transform 1 0 27552 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_250
timestamp 1698431365
transform 1 0 29344 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_266
timestamp 1698431365
transform 1 0 31136 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_270
timestamp 1698431365
transform 1 0 31584 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_274
timestamp 1698431365
transform 1 0 32032 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_276
timestamp 1698431365
transform 1 0 32256 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_281
timestamp 1698431365
transform 1 0 32816 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_297
timestamp 1698431365
transform 1 0 34608 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_305
timestamp 1698431365
transform 1 0 35504 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_308
timestamp 1698431365
transform 1 0 35840 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_316
timestamp 1698431365
transform 1 0 36736 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_318
timestamp 1698431365
transform 1 0 36960 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input1 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 38416 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input2 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 38416 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input3
timestamp 1698431365
transform -1 0 37296 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input4
timestamp 1698431365
transform 1 0 3808 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input5
timestamp 1698431365
transform 1 0 15904 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input6
timestamp 1698431365
transform -1 0 17584 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input7
timestamp 1698431365
transform 1 0 17808 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input8
timestamp 1698431365
transform 1 0 18704 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input9
timestamp 1698431365
transform 1 0 19600 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input10
timestamp 1698431365
transform 1 0 20608 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input11
timestamp 1698431365
transform 1 0 21392 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input12
timestamp 1698431365
transform 1 0 22288 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input13
timestamp 1698431365
transform 1 0 23184 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input14
timestamp 1698431365
transform -1 0 25088 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input15
timestamp 1698431365
transform 1 0 5600 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input16
timestamp 1698431365
transform 1 0 25088 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input17
timestamp 1698431365
transform -1 0 26544 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input18
timestamp 1698431365
transform -1 0 27440 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input19
timestamp 1698431365
transform -1 0 28896 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input20
timestamp 1698431365
transform 1 0 28896 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input21
timestamp 1698431365
transform 1 0 29568 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input22
timestamp 1698431365
transform 1 0 30352 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input23
timestamp 1698431365
transform 1 0 31136 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input24
timestamp 1698431365
transform -1 0 33600 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input25
timestamp 1698431365
transform -1 0 34272 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input26
timestamp 1698431365
transform 1 0 8512 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input27
timestamp 1698431365
transform -1 0 35616 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input28
timestamp 1698431365
transform -1 0 36512 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input29
timestamp 1698431365
transform 1 0 6944 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input30
timestamp 1698431365
transform 1 0 7616 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input31
timestamp 1698431365
transform 1 0 9632 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input32
timestamp 1698431365
transform 1 0 8288 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input33
timestamp 1698431365
transform 1 0 10304 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input34
timestamp 1698431365
transform 1 0 13552 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input35
timestamp 1698431365
transform 1 0 15904 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input36
timestamp 1698431365
transform 1 0 3920 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input37
timestamp 1698431365
transform 1 0 4480 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input38
timestamp 1698431365
transform 1 0 6272 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input39
timestamp 1698431365
transform 1 0 3248 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input40
timestamp 1698431365
transform 1 0 3136 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input41
timestamp 1698431365
transform -1 0 38192 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output42 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 28224 0 1 45472
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output43
timestamp 1698431365
transform 1 0 37296 0 1 45472
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output44
timestamp 1698431365
transform 1 0 1568 0 1 3136
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output45
timestamp 1698431365
transform -1 0 3136 0 1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output46 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 3136 0 -1 7840
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output47
timestamp 1698431365
transform -1 0 3920 0 1 45472
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output48
timestamp 1698431365
transform -1 0 14560 0 1 45472
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_55 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698431365
transform -1 0 38640 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_56
timestamp 1698431365
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698431365
transform -1 0 38640 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_57
timestamp 1698431365
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698431365
transform -1 0 38640 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_58
timestamp 1698431365
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698431365
transform -1 0 38640 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_59
timestamp 1698431365
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698431365
transform -1 0 38640 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_60
timestamp 1698431365
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698431365
transform -1 0 38640 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_61
timestamp 1698431365
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698431365
transform -1 0 38640 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_62
timestamp 1698431365
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698431365
transform -1 0 38640 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_63
timestamp 1698431365
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698431365
transform -1 0 38640 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_64
timestamp 1698431365
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698431365
transform -1 0 38640 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_65
timestamp 1698431365
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698431365
transform -1 0 38640 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_66
timestamp 1698431365
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698431365
transform -1 0 38640 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_67
timestamp 1698431365
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698431365
transform -1 0 38640 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_68
timestamp 1698431365
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698431365
transform -1 0 38640 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_69
timestamp 1698431365
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698431365
transform -1 0 38640 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_70
timestamp 1698431365
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698431365
transform -1 0 38640 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_71
timestamp 1698431365
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698431365
transform -1 0 38640 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_72
timestamp 1698431365
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698431365
transform -1 0 38640 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_73
timestamp 1698431365
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698431365
transform -1 0 38640 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_74
timestamp 1698431365
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698431365
transform -1 0 38640 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_75
timestamp 1698431365
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698431365
transform -1 0 38640 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_76
timestamp 1698431365
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698431365
transform -1 0 38640 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_77
timestamp 1698431365
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698431365
transform -1 0 38640 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_78
timestamp 1698431365
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698431365
transform -1 0 38640 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_79
timestamp 1698431365
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698431365
transform -1 0 38640 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_80
timestamp 1698431365
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698431365
transform -1 0 38640 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_81
timestamp 1698431365
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698431365
transform -1 0 38640 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_82
timestamp 1698431365
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698431365
transform -1 0 38640 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_83
timestamp 1698431365
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698431365
transform -1 0 38640 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_84
timestamp 1698431365
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698431365
transform -1 0 38640 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_85
timestamp 1698431365
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698431365
transform -1 0 38640 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_86
timestamp 1698431365
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698431365
transform -1 0 38640 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_87
timestamp 1698431365
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698431365
transform -1 0 38640 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_88
timestamp 1698431365
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698431365
transform -1 0 38640 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_89
timestamp 1698431365
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698431365
transform -1 0 38640 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_90
timestamp 1698431365
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698431365
transform -1 0 38640 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_91
timestamp 1698431365
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698431365
transform -1 0 38640 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_92
timestamp 1698431365
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698431365
transform -1 0 38640 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_93
timestamp 1698431365
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698431365
transform -1 0 38640 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_94
timestamp 1698431365
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698431365
transform -1 0 38640 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_95
timestamp 1698431365
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698431365
transform -1 0 38640 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_96
timestamp 1698431365
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698431365
transform -1 0 38640 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_97
timestamp 1698431365
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698431365
transform -1 0 38640 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_98
timestamp 1698431365
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698431365
transform -1 0 38640 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_99
timestamp 1698431365
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698431365
transform -1 0 38640 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Left_100
timestamp 1698431365
transform 1 0 1344 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Right_45
timestamp 1698431365
transform -1 0 38640 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Left_101
timestamp 1698431365
transform 1 0 1344 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Right_46
timestamp 1698431365
transform -1 0 38640 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Left_102
timestamp 1698431365
transform 1 0 1344 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Right_47
timestamp 1698431365
transform -1 0 38640 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Left_103
timestamp 1698431365
transform 1 0 1344 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Right_48
timestamp 1698431365
transform -1 0 38640 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Left_104
timestamp 1698431365
transform 1 0 1344 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Right_49
timestamp 1698431365
transform -1 0 38640 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Left_105
timestamp 1698431365
transform 1 0 1344 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Right_50
timestamp 1698431365
transform -1 0 38640 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Left_106
timestamp 1698431365
transform 1 0 1344 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Right_51
timestamp 1698431365
transform -1 0 38640 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Left_107
timestamp 1698431365
transform 1 0 1344 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Right_52
timestamp 1698431365
transform -1 0 38640 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Left_108
timestamp 1698431365
transform 1 0 1344 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Right_53
timestamp 1698431365
transform -1 0 38640 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Left_109
timestamp 1698431365
transform 1 0 1344 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Right_54
timestamp 1698431365
transform -1 0 38640 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_110 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_111
timestamp 1698431365
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_112
timestamp 1698431365
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_113
timestamp 1698431365
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_114
timestamp 1698431365
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_115
timestamp 1698431365
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_116
timestamp 1698431365
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_117
timestamp 1698431365
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_118
timestamp 1698431365
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_119
timestamp 1698431365
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_120
timestamp 1698431365
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_121
timestamp 1698431365
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_122
timestamp 1698431365
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_123
timestamp 1698431365
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_124
timestamp 1698431365
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_125
timestamp 1698431365
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_126
timestamp 1698431365
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_127
timestamp 1698431365
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_128
timestamp 1698431365
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_129
timestamp 1698431365
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_130
timestamp 1698431365
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_131
timestamp 1698431365
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_132
timestamp 1698431365
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_133
timestamp 1698431365
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_134
timestamp 1698431365
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_135
timestamp 1698431365
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_136
timestamp 1698431365
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_137
timestamp 1698431365
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_138
timestamp 1698431365
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_139
timestamp 1698431365
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_140
timestamp 1698431365
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_141
timestamp 1698431365
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_142
timestamp 1698431365
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_143
timestamp 1698431365
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_144
timestamp 1698431365
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_145
timestamp 1698431365
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_146
timestamp 1698431365
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_147
timestamp 1698431365
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_148
timestamp 1698431365
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_149
timestamp 1698431365
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_150
timestamp 1698431365
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_151
timestamp 1698431365
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_152
timestamp 1698431365
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_153
timestamp 1698431365
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_154
timestamp 1698431365
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_155
timestamp 1698431365
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_156
timestamp 1698431365
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_157
timestamp 1698431365
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_158
timestamp 1698431365
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_159
timestamp 1698431365
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_160
timestamp 1698431365
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_161
timestamp 1698431365
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_162
timestamp 1698431365
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_163
timestamp 1698431365
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_164
timestamp 1698431365
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_165
timestamp 1698431365
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_166
timestamp 1698431365
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_167
timestamp 1698431365
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_168
timestamp 1698431365
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_169
timestamp 1698431365
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_170
timestamp 1698431365
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_171
timestamp 1698431365
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_172
timestamp 1698431365
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_173
timestamp 1698431365
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_174
timestamp 1698431365
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_175
timestamp 1698431365
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_176
timestamp 1698431365
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_177
timestamp 1698431365
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_178
timestamp 1698431365
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_179
timestamp 1698431365
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_180
timestamp 1698431365
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_181
timestamp 1698431365
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_182
timestamp 1698431365
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_183
timestamp 1698431365
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_184
timestamp 1698431365
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_185
timestamp 1698431365
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_186
timestamp 1698431365
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_187
timestamp 1698431365
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_188
timestamp 1698431365
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_189
timestamp 1698431365
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_190
timestamp 1698431365
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_191
timestamp 1698431365
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_192
timestamp 1698431365
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_193
timestamp 1698431365
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_194
timestamp 1698431365
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_195
timestamp 1698431365
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_196
timestamp 1698431365
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_197
timestamp 1698431365
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_198
timestamp 1698431365
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_199
timestamp 1698431365
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_200
timestamp 1698431365
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_201
timestamp 1698431365
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_202
timestamp 1698431365
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_203
timestamp 1698431365
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_204
timestamp 1698431365
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_205
timestamp 1698431365
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_206
timestamp 1698431365
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_207
timestamp 1698431365
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_208
timestamp 1698431365
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_209
timestamp 1698431365
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_210
timestamp 1698431365
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_211
timestamp 1698431365
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_212
timestamp 1698431365
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_213
timestamp 1698431365
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_214
timestamp 1698431365
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_215
timestamp 1698431365
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_216
timestamp 1698431365
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_217
timestamp 1698431365
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_218
timestamp 1698431365
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_219
timestamp 1698431365
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_220
timestamp 1698431365
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_221
timestamp 1698431365
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_222
timestamp 1698431365
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_223
timestamp 1698431365
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_224
timestamp 1698431365
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_225
timestamp 1698431365
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_226
timestamp 1698431365
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_227
timestamp 1698431365
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_228
timestamp 1698431365
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_229
timestamp 1698431365
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_230
timestamp 1698431365
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_231
timestamp 1698431365
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_232
timestamp 1698431365
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_233
timestamp 1698431365
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_234
timestamp 1698431365
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_235
timestamp 1698431365
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_236
timestamp 1698431365
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_237
timestamp 1698431365
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_238
timestamp 1698431365
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_239
timestamp 1698431365
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_240
timestamp 1698431365
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_241
timestamp 1698431365
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_242
timestamp 1698431365
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_243
timestamp 1698431365
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_244
timestamp 1698431365
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_245
timestamp 1698431365
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_246
timestamp 1698431365
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_247
timestamp 1698431365
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_248
timestamp 1698431365
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_249
timestamp 1698431365
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_250
timestamp 1698431365
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_251
timestamp 1698431365
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_252
timestamp 1698431365
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_253
timestamp 1698431365
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_254
timestamp 1698431365
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_255
timestamp 1698431365
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_256
timestamp 1698431365
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_257
timestamp 1698431365
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_258
timestamp 1698431365
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_259
timestamp 1698431365
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_260
timestamp 1698431365
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_261
timestamp 1698431365
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_262
timestamp 1698431365
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_263
timestamp 1698431365
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_264
timestamp 1698431365
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_265
timestamp 1698431365
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_266
timestamp 1698431365
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_267
timestamp 1698431365
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_268
timestamp 1698431365
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_269
timestamp 1698431365
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_270
timestamp 1698431365
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_271
timestamp 1698431365
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_272
timestamp 1698431365
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_273
timestamp 1698431365
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_274
timestamp 1698431365
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_275
timestamp 1698431365
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_276
timestamp 1698431365
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_277
timestamp 1698431365
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_278
timestamp 1698431365
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_279
timestamp 1698431365
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_280
timestamp 1698431365
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_281
timestamp 1698431365
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_282
timestamp 1698431365
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_283
timestamp 1698431365
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_284
timestamp 1698431365
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_285
timestamp 1698431365
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_286
timestamp 1698431365
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_287
timestamp 1698431365
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_288
timestamp 1698431365
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_289
timestamp 1698431365
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_290
timestamp 1698431365
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_291
timestamp 1698431365
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_292
timestamp 1698431365
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_293
timestamp 1698431365
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_294
timestamp 1698431365
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_295
timestamp 1698431365
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_296
timestamp 1698431365
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_297
timestamp 1698431365
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_298
timestamp 1698431365
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_299
timestamp 1698431365
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_300
timestamp 1698431365
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_301
timestamp 1698431365
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_302
timestamp 1698431365
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_303
timestamp 1698431365
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_304
timestamp 1698431365
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_305
timestamp 1698431365
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_306
timestamp 1698431365
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_307
timestamp 1698431365
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_308
timestamp 1698431365
transform 1 0 9184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_309
timestamp 1698431365
transform 1 0 17024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_310
timestamp 1698431365
transform 1 0 24864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_311
timestamp 1698431365
transform 1 0 32704 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_312
timestamp 1698431365
transform 1 0 5264 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_313
timestamp 1698431365
transform 1 0 13104 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_314
timestamp 1698431365
transform 1 0 20944 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_315
timestamp 1698431365
transform 1 0 28784 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_316
timestamp 1698431365
transform 1 0 36624 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_317
timestamp 1698431365
transform 1 0 9184 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_318
timestamp 1698431365
transform 1 0 17024 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_319
timestamp 1698431365
transform 1 0 24864 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_320
timestamp 1698431365
transform 1 0 32704 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_321
timestamp 1698431365
transform 1 0 5264 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_322
timestamp 1698431365
transform 1 0 13104 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_323
timestamp 1698431365
transform 1 0 20944 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_324
timestamp 1698431365
transform 1 0 28784 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_325
timestamp 1698431365
transform 1 0 36624 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_326
timestamp 1698431365
transform 1 0 9184 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_327
timestamp 1698431365
transform 1 0 17024 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_328
timestamp 1698431365
transform 1 0 24864 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_329
timestamp 1698431365
transform 1 0 32704 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_330
timestamp 1698431365
transform 1 0 5264 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_331
timestamp 1698431365
transform 1 0 13104 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_332
timestamp 1698431365
transform 1 0 20944 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_333
timestamp 1698431365
transform 1 0 28784 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_334
timestamp 1698431365
transform 1 0 36624 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_335
timestamp 1698431365
transform 1 0 9184 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_336
timestamp 1698431365
transform 1 0 17024 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_337
timestamp 1698431365
transform 1 0 24864 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_338
timestamp 1698431365
transform 1 0 32704 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_339
timestamp 1698431365
transform 1 0 5264 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_340
timestamp 1698431365
transform 1 0 13104 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_341
timestamp 1698431365
transform 1 0 20944 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_342
timestamp 1698431365
transform 1 0 28784 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_343
timestamp 1698431365
transform 1 0 36624 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_344
timestamp 1698431365
transform 1 0 9184 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_345
timestamp 1698431365
transform 1 0 17024 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_346
timestamp 1698431365
transform 1 0 24864 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_347
timestamp 1698431365
transform 1 0 32704 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_348
timestamp 1698431365
transform 1 0 5264 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_349
timestamp 1698431365
transform 1 0 13104 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_350
timestamp 1698431365
transform 1 0 20944 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_351
timestamp 1698431365
transform 1 0 28784 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_352
timestamp 1698431365
transform 1 0 36624 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_353
timestamp 1698431365
transform 1 0 9184 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_354
timestamp 1698431365
transform 1 0 17024 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_355
timestamp 1698431365
transform 1 0 24864 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_356
timestamp 1698431365
transform 1 0 32704 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_357
timestamp 1698431365
transform 1 0 5152 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_358
timestamp 1698431365
transform 1 0 8960 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_359
timestamp 1698431365
transform 1 0 12768 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_360
timestamp 1698431365
transform 1 0 16576 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_361
timestamp 1698431365
transform 1 0 20384 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_362
timestamp 1698431365
transform 1 0 24192 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_363
timestamp 1698431365
transform 1 0 28000 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_364
timestamp 1698431365
transform 1 0 31808 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_365
timestamp 1698431365
transform 1 0 35616 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_49 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 37968 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_50
timestamp 1698431365
transform -1 0 22960 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_51
timestamp 1698431365
transform -1 0 32816 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_52
timestamp 1698431365
transform -1 0 2016 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_53
timestamp 1698431365
transform -1 0 2016 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_54
timestamp 1698431365
transform -1 0 2016 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_55
timestamp 1698431365
transform -1 0 2016 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_56
timestamp 1698431365
transform -1 0 2016 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_57
timestamp 1698431365
transform -1 0 2016 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_58
timestamp 1698431365
transform -1 0 2016 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_59
timestamp 1698431365
transform -1 0 2016 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_60
timestamp 1698431365
transform -1 0 2016 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_61
timestamp 1698431365
transform -1 0 2016 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_62
timestamp 1698431365
transform -1 0 2016 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_63
timestamp 1698431365
transform -1 0 2016 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_64
timestamp 1698431365
transform -1 0 2016 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_65
timestamp 1698431365
transform -1 0 2016 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_66
timestamp 1698431365
transform -1 0 2016 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_67
timestamp 1698431365
transform -1 0 2016 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_68
timestamp 1698431365
transform -1 0 2016 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_69
timestamp 1698431365
transform -1 0 2016 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_70
timestamp 1698431365
transform -1 0 2016 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_71
timestamp 1698431365
transform -1 0 2016 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_72
timestamp 1698431365
transform -1 0 2016 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_73
timestamp 1698431365
transform -1 0 2016 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_74
timestamp 1698431365
transform -1 0 2016 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_75
timestamp 1698431365
transform -1 0 2016 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_76
timestamp 1698431365
transform -1 0 2016 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_77
timestamp 1698431365
transform -1 0 2016 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_78
timestamp 1698431365
transform -1 0 2016 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_79
timestamp 1698431365
transform -1 0 2016 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_80
timestamp 1698431365
transform -1 0 2464 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_81
timestamp 1698431365
transform -1 0 2352 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_82
timestamp 1698431365
transform -1 0 2016 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_83
timestamp 1698431365
transform -1 0 8176 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_84
timestamp 1698431365
transform -1 0 18032 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  wb_buttons_leds_85 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 37968 0 -1 43904
box -86 -86 534 870
<< labels >>
flabel metal3 s 39200 6272 40000 6384 0 FreeSans 448 0 0 0 buttons[0]
port 0 nsew signal input
flabel metal3 s 39200 30912 40000 31024 0 FreeSans 448 0 0 0 buttons[1]
port 1 nsew signal input
flabel metal3 s 39200 43232 40000 43344 0 FreeSans 448 0 0 0 buttons_enb[0]
port 2 nsew signal tristate
flabel metal3 s 39200 18592 40000 18704 0 FreeSans 448 0 0 0 buttons_enb[1]
port 3 nsew signal tristate
flabel metal2 s 35616 0 35728 800 0 FreeSans 448 90 0 0 clk
port 4 nsew signal input
flabel metal2 s 36512 0 36624 800 0 FreeSans 448 90 0 0 clk2
port 5 nsew signal input
flabel metal2 s 5152 0 5264 800 0 FreeSans 448 90 0 0 i_wb_addr[0]
port 6 nsew signal input
flabel metal2 s 15904 0 16016 800 0 FreeSans 448 90 0 0 i_wb_addr[10]
port 7 nsew signal input
flabel metal2 s 16800 0 16912 800 0 FreeSans 448 90 0 0 i_wb_addr[11]
port 8 nsew signal input
flabel metal2 s 17696 0 17808 800 0 FreeSans 448 90 0 0 i_wb_addr[12]
port 9 nsew signal input
flabel metal2 s 18592 0 18704 800 0 FreeSans 448 90 0 0 i_wb_addr[13]
port 10 nsew signal input
flabel metal2 s 19488 0 19600 800 0 FreeSans 448 90 0 0 i_wb_addr[14]
port 11 nsew signal input
flabel metal2 s 20384 0 20496 800 0 FreeSans 448 90 0 0 i_wb_addr[15]
port 12 nsew signal input
flabel metal2 s 21280 0 21392 800 0 FreeSans 448 90 0 0 i_wb_addr[16]
port 13 nsew signal input
flabel metal2 s 22176 0 22288 800 0 FreeSans 448 90 0 0 i_wb_addr[17]
port 14 nsew signal input
flabel metal2 s 23072 0 23184 800 0 FreeSans 448 90 0 0 i_wb_addr[18]
port 15 nsew signal input
flabel metal2 s 23968 0 24080 800 0 FreeSans 448 90 0 0 i_wb_addr[19]
port 16 nsew signal input
flabel metal2 s 6944 0 7056 800 0 FreeSans 448 90 0 0 i_wb_addr[1]
port 17 nsew signal input
flabel metal2 s 24864 0 24976 800 0 FreeSans 448 90 0 0 i_wb_addr[20]
port 18 nsew signal input
flabel metal2 s 25760 0 25872 800 0 FreeSans 448 90 0 0 i_wb_addr[21]
port 19 nsew signal input
flabel metal2 s 26656 0 26768 800 0 FreeSans 448 90 0 0 i_wb_addr[22]
port 20 nsew signal input
flabel metal2 s 27552 0 27664 800 0 FreeSans 448 90 0 0 i_wb_addr[23]
port 21 nsew signal input
flabel metal2 s 28448 0 28560 800 0 FreeSans 448 90 0 0 i_wb_addr[24]
port 22 nsew signal input
flabel metal2 s 29344 0 29456 800 0 FreeSans 448 90 0 0 i_wb_addr[25]
port 23 nsew signal input
flabel metal2 s 30240 0 30352 800 0 FreeSans 448 90 0 0 i_wb_addr[26]
port 24 nsew signal input
flabel metal2 s 31136 0 31248 800 0 FreeSans 448 90 0 0 i_wb_addr[27]
port 25 nsew signal input
flabel metal2 s 32032 0 32144 800 0 FreeSans 448 90 0 0 i_wb_addr[28]
port 26 nsew signal input
flabel metal2 s 32928 0 33040 800 0 FreeSans 448 90 0 0 i_wb_addr[29]
port 27 nsew signal input
flabel metal2 s 8736 0 8848 800 0 FreeSans 448 90 0 0 i_wb_addr[2]
port 28 nsew signal input
flabel metal2 s 33824 0 33936 800 0 FreeSans 448 90 0 0 i_wb_addr[30]
port 29 nsew signal input
flabel metal2 s 34720 0 34832 800 0 FreeSans 448 90 0 0 i_wb_addr[31]
port 30 nsew signal input
flabel metal2 s 9632 0 9744 800 0 FreeSans 448 90 0 0 i_wb_addr[3]
port 31 nsew signal input
flabel metal2 s 10528 0 10640 800 0 FreeSans 448 90 0 0 i_wb_addr[4]
port 32 nsew signal input
flabel metal2 s 11424 0 11536 800 0 FreeSans 448 90 0 0 i_wb_addr[5]
port 33 nsew signal input
flabel metal2 s 12320 0 12432 800 0 FreeSans 448 90 0 0 i_wb_addr[6]
port 34 nsew signal input
flabel metal2 s 13216 0 13328 800 0 FreeSans 448 90 0 0 i_wb_addr[7]
port 35 nsew signal input
flabel metal2 s 14112 0 14224 800 0 FreeSans 448 90 0 0 i_wb_addr[8]
port 36 nsew signal input
flabel metal2 s 15008 0 15120 800 0 FreeSans 448 90 0 0 i_wb_addr[9]
port 37 nsew signal input
flabel metal2 s 2464 0 2576 800 0 FreeSans 448 90 0 0 i_wb_cyc
port 38 nsew signal input
flabel metal2 s 6048 0 6160 800 0 FreeSans 448 90 0 0 i_wb_data[0]
port 39 nsew signal input
flabel metal2 s 7840 0 7952 800 0 FreeSans 448 90 0 0 i_wb_data[1]
port 40 nsew signal input
flabel metal2 s 3360 0 3472 800 0 FreeSans 448 90 0 0 i_wb_stb
port 41 nsew signal input
flabel metal2 s 4256 0 4368 800 0 FreeSans 448 90 0 0 i_wb_we
port 42 nsew signal input
flabel metal2 s 22400 49200 22512 50000 0 FreeSans 448 90 0 0 led_enb[0]
port 43 nsew signal tristate
flabel metal2 s 32256 49200 32368 50000 0 FreeSans 448 90 0 0 led_enb[1]
port 44 nsew signal tristate
flabel metal2 s 27328 49200 27440 50000 0 FreeSans 448 90 0 0 leds[0]
port 45 nsew signal tristate
flabel metal2 s 37184 49200 37296 50000 0 FreeSans 448 90 0 0 leds[1]
port 46 nsew signal tristate
flabel metal3 s 0 2688 800 2800 0 FreeSans 448 0 0 0 o_wb_ack
port 47 nsew signal tristate
flabel metal3 s 0 5376 800 5488 0 FreeSans 448 0 0 0 o_wb_data[0]
port 48 nsew signal tristate
flabel metal3 s 0 18816 800 18928 0 FreeSans 448 0 0 0 o_wb_data[10]
port 49 nsew signal tristate
flabel metal3 s 0 20160 800 20272 0 FreeSans 448 0 0 0 o_wb_data[11]
port 50 nsew signal tristate
flabel metal3 s 0 21504 800 21616 0 FreeSans 448 0 0 0 o_wb_data[12]
port 51 nsew signal tristate
flabel metal3 s 0 22848 800 22960 0 FreeSans 448 0 0 0 o_wb_data[13]
port 52 nsew signal tristate
flabel metal3 s 0 24192 800 24304 0 FreeSans 448 0 0 0 o_wb_data[14]
port 53 nsew signal tristate
flabel metal3 s 0 25536 800 25648 0 FreeSans 448 0 0 0 o_wb_data[15]
port 54 nsew signal tristate
flabel metal3 s 0 26880 800 26992 0 FreeSans 448 0 0 0 o_wb_data[16]
port 55 nsew signal tristate
flabel metal3 s 0 28224 800 28336 0 FreeSans 448 0 0 0 o_wb_data[17]
port 56 nsew signal tristate
flabel metal3 s 0 29568 800 29680 0 FreeSans 448 0 0 0 o_wb_data[18]
port 57 nsew signal tristate
flabel metal3 s 0 30912 800 31024 0 FreeSans 448 0 0 0 o_wb_data[19]
port 58 nsew signal tristate
flabel metal3 s 0 6720 800 6832 0 FreeSans 448 0 0 0 o_wb_data[1]
port 59 nsew signal tristate
flabel metal3 s 0 32256 800 32368 0 FreeSans 448 0 0 0 o_wb_data[20]
port 60 nsew signal tristate
flabel metal3 s 0 33600 800 33712 0 FreeSans 448 0 0 0 o_wb_data[21]
port 61 nsew signal tristate
flabel metal3 s 0 34944 800 35056 0 FreeSans 448 0 0 0 o_wb_data[22]
port 62 nsew signal tristate
flabel metal3 s 0 36288 800 36400 0 FreeSans 448 0 0 0 o_wb_data[23]
port 63 nsew signal tristate
flabel metal3 s 0 37632 800 37744 0 FreeSans 448 0 0 0 o_wb_data[24]
port 64 nsew signal tristate
flabel metal3 s 0 38976 800 39088 0 FreeSans 448 0 0 0 o_wb_data[25]
port 65 nsew signal tristate
flabel metal3 s 0 40320 800 40432 0 FreeSans 448 0 0 0 o_wb_data[26]
port 66 nsew signal tristate
flabel metal3 s 0 41664 800 41776 0 FreeSans 448 0 0 0 o_wb_data[27]
port 67 nsew signal tristate
flabel metal3 s 0 43008 800 43120 0 FreeSans 448 0 0 0 o_wb_data[28]
port 68 nsew signal tristate
flabel metal3 s 0 44352 800 44464 0 FreeSans 448 0 0 0 o_wb_data[29]
port 69 nsew signal tristate
flabel metal3 s 0 8064 800 8176 0 FreeSans 448 0 0 0 o_wb_data[2]
port 70 nsew signal tristate
flabel metal3 s 0 45696 800 45808 0 FreeSans 448 0 0 0 o_wb_data[30]
port 71 nsew signal tristate
flabel metal3 s 0 47040 800 47152 0 FreeSans 448 0 0 0 o_wb_data[31]
port 72 nsew signal tristate
flabel metal3 s 0 9408 800 9520 0 FreeSans 448 0 0 0 o_wb_data[3]
port 73 nsew signal tristate
flabel metal3 s 0 10752 800 10864 0 FreeSans 448 0 0 0 o_wb_data[4]
port 74 nsew signal tristate
flabel metal3 s 0 12096 800 12208 0 FreeSans 448 0 0 0 o_wb_data[5]
port 75 nsew signal tristate
flabel metal3 s 0 13440 800 13552 0 FreeSans 448 0 0 0 o_wb_data[6]
port 76 nsew signal tristate
flabel metal3 s 0 14784 800 14896 0 FreeSans 448 0 0 0 o_wb_data[7]
port 77 nsew signal tristate
flabel metal3 s 0 16128 800 16240 0 FreeSans 448 0 0 0 o_wb_data[8]
port 78 nsew signal tristate
flabel metal3 s 0 17472 800 17584 0 FreeSans 448 0 0 0 o_wb_data[9]
port 79 nsew signal tristate
flabel metal3 s 0 4032 800 4144 0 FreeSans 448 0 0 0 o_wb_stall
port 80 nsew signal tristate
flabel metal2 s 37408 0 37520 800 0 FreeSans 448 90 0 0 reset
port 81 nsew signal input
flabel metal4 s 3988 3076 5228 46316 0 FreeSans 5120 90 0 0 vdd
port 82 nsew power bidirectional
flabel metal4 s 23988 3076 25228 46316 0 FreeSans 5120 90 0 0 vdd
port 82 nsew power bidirectional
flabel metal4 s 13988 3076 15228 46316 0 FreeSans 5120 90 0 0 vss
port 83 nsew ground bidirectional
flabel metal4 s 33988 3076 35228 46316 0 FreeSans 5120 90 0 0 vss
port 83 nsew ground bidirectional
flabel metal2 s 7616 49200 7728 50000 0 FreeSans 448 90 0 0 xtal_clk[0]
port 84 nsew signal tristate
flabel metal2 s 17472 49200 17584 50000 0 FreeSans 448 90 0 0 xtal_clk[1]
port 85 nsew signal tristate
flabel metal2 s 2688 49200 2800 50000 0 FreeSans 448 90 0 0 xtal_clk_enb[0]
port 86 nsew signal tristate
flabel metal2 s 12544 49200 12656 50000 0 FreeSans 448 90 0 0 xtal_clk_enb[1]
port 87 nsew signal tristate
rlabel metal1 19992 46256 19992 46256 0 vdd
rlabel metal1 19992 45472 19992 45472 0 vss
rlabel metal2 15176 6944 15176 6944 0 _000_
rlabel metal2 2072 5096 2072 5096 0 _001_
rlabel metal3 5432 5768 5432 5768 0 _002_
rlabel metal3 7224 7336 7224 7336 0 _003_
rlabel metal2 8904 5712 8904 5712 0 _004_
rlabel metal2 10472 9464 10472 9464 0 _005_
rlabel metal2 8176 5992 8176 5992 0 _006_
rlabel metal2 11200 4536 11200 4536 0 _007_
rlabel metal2 9464 4312 9464 4312 0 _008_
rlabel metal2 7504 4424 7504 4424 0 _009_
rlabel metal2 7448 6272 7448 6272 0 _010_
rlabel metal2 18648 3976 18648 3976 0 _011_
rlabel metal2 15288 3976 15288 3976 0 _012_
rlabel metal2 15512 5488 15512 5488 0 _013_
rlabel metal2 13160 6944 13160 6944 0 _014_
rlabel metal2 24136 4424 24136 4424 0 _015_
rlabel metal2 23800 4648 23800 4648 0 _016_
rlabel metal2 14728 4256 14728 4256 0 _017_
rlabel metal2 34440 3808 34440 3808 0 _018_
rlabel metal3 34216 3416 34216 3416 0 _019_
rlabel metal3 31920 4368 31920 4368 0 _020_
rlabel metal2 9912 4648 9912 4648 0 _021_
rlabel metal2 11088 3528 11088 3528 0 _022_
rlabel metal2 12264 5208 12264 5208 0 _023_
rlabel metal2 9016 7784 9016 7784 0 _024_
rlabel metal2 6552 7112 6552 7112 0 _025_
rlabel metal3 9744 5992 9744 5992 0 _026_
rlabel metal2 8120 4480 8120 4480 0 _027_
rlabel metal2 2296 6216 2296 6216 0 _028_
rlabel metal2 5096 4928 5096 4928 0 _029_
rlabel metal2 7784 6328 7784 6328 0 _030_
rlabel metal2 6328 5208 6328 5208 0 _031_
rlabel metal2 5992 6832 5992 6832 0 _032_
rlabel metal2 11480 4032 11480 4032 0 _033_
rlabel metal2 6608 5992 6608 5992 0 _034_
rlabel metal2 6888 6160 6888 6160 0 _035_
rlabel metal3 8456 7448 8456 7448 0 _036_
rlabel metal2 7280 6776 7280 6776 0 _037_
rlabel metal2 12152 4368 12152 4368 0 _038_
rlabel metal2 11480 4704 11480 4704 0 _039_
rlabel metal2 11592 5544 11592 5544 0 _040_
rlabel metal2 10808 9800 10808 9800 0 _041_
rlabel metal2 38248 6440 38248 6440 0 buttons[0]
rlabel metal2 38248 31248 38248 31248 0 buttons[1]
rlabel metal2 35672 2478 35672 2478 0 clk
rlabel metal2 36960 3528 36960 3528 0 clk2
rlabel metal2 11368 7504 11368 7504 0 clknet_0_clk
rlabel metal2 5544 5544 5544 5544 0 clknet_1_0__leaf_clk
rlabel metal2 9800 9184 9800 9184 0 clknet_1_1__leaf_clk
rlabel metal2 3864 3528 3864 3528 0 i_wb_addr[0]
rlabel metal2 15960 2058 15960 2058 0 i_wb_addr[10]
rlabel metal2 17080 3080 17080 3080 0 i_wb_addr[11]
rlabel metal2 17752 2058 17752 2058 0 i_wb_addr[12]
rlabel metal2 18648 2058 18648 2058 0 i_wb_addr[13]
rlabel metal2 19656 3528 19656 3528 0 i_wb_addr[14]
rlabel metal2 20440 2058 20440 2058 0 i_wb_addr[15]
rlabel metal2 21336 2058 21336 2058 0 i_wb_addr[16]
rlabel metal2 22120 4872 22120 4872 0 i_wb_addr[17]
rlabel metal2 23128 2058 23128 2058 0 i_wb_addr[18]
rlabel metal2 24528 728 24528 728 0 i_wb_addr[19]
rlabel metal2 5768 4256 5768 4256 0 i_wb_addr[1]
rlabel metal2 25032 2184 25032 2184 0 i_wb_addr[20]
rlabel metal2 26040 2744 26040 2744 0 i_wb_addr[21]
rlabel metal2 27160 3472 27160 3472 0 i_wb_addr[22]
rlabel metal3 28112 3528 28112 3528 0 i_wb_addr[23]
rlabel metal3 28784 3416 28784 3416 0 i_wb_addr[24]
rlabel metal2 29736 2968 29736 2968 0 i_wb_addr[25]
rlabel metal2 30520 2968 30520 2968 0 i_wb_addr[26]
rlabel metal2 31248 3416 31248 3416 0 i_wb_addr[27]
rlabel metal2 32536 3976 32536 3976 0 i_wb_addr[28]
rlabel metal3 33600 4312 33600 4312 0 i_wb_addr[29]
rlabel metal2 8792 1246 8792 1246 0 i_wb_addr[2]
rlabel metal2 35336 3976 35336 3976 0 i_wb_addr[30]
rlabel metal2 36232 3472 36232 3472 0 i_wb_addr[31]
rlabel metal2 7112 3136 7112 3136 0 i_wb_addr[3]
rlabel metal2 10584 1974 10584 1974 0 i_wb_addr[4]
rlabel metal2 9800 5432 9800 5432 0 i_wb_addr[5]
rlabel metal2 3080 3864 3080 3864 0 i_wb_addr[6]
rlabel metal2 13272 2058 13272 2058 0 i_wb_addr[7]
rlabel metal2 14168 854 14168 854 0 i_wb_addr[8]
rlabel metal2 16072 4480 16072 4480 0 i_wb_addr[9]
rlabel metal2 2520 2926 2520 2926 0 i_wb_cyc
rlabel metal2 6104 1246 6104 1246 0 i_wb_data[0]
rlabel metal2 6552 3640 6552 3640 0 i_wb_data[1]
rlabel metal2 3192 3528 3192 3528 0 i_wb_stb
rlabel metal2 3304 3584 3304 3584 0 i_wb_we
rlabel metal2 28840 46032 28840 46032 0 leds[0]
rlabel metal2 37912 46256 37912 46256 0 leds[1]
rlabel metal2 37912 7448 37912 7448 0 net1
rlabel metal2 21112 3640 21112 3640 0 net10
rlabel metal2 21896 4256 21896 4256 0 net11
rlabel metal2 22848 3416 22848 3416 0 net12
rlabel metal2 23688 4200 23688 4200 0 net13
rlabel metal3 25200 3416 25200 3416 0 net14
rlabel metal2 10136 4648 10136 4648 0 net15
rlabel metal2 25368 3864 25368 3864 0 net16
rlabel metal2 26040 3920 26040 3920 0 net17
rlabel metal2 26936 3976 26936 3976 0 net18
rlabel metal2 28392 3640 28392 3640 0 net19
rlabel metal2 37912 20608 37912 20608 0 net2
rlabel metal2 29400 3752 29400 3752 0 net20
rlabel metal2 30184 3416 30184 3416 0 net21
rlabel metal2 30856 4200 30856 4200 0 net22
rlabel metal2 31640 3360 31640 3360 0 net23
rlabel metal2 33096 3976 33096 3976 0 net24
rlabel metal2 33768 3920 33768 3920 0 net25
rlabel metal3 7504 6552 7504 6552 0 net26
rlabel metal2 34944 4424 34944 4424 0 net27
rlabel metal2 36008 3360 36008 3360 0 net28
rlabel metal2 10024 5432 10024 5432 0 net29
rlabel metal2 36792 3360 36792 3360 0 net3
rlabel metal4 15736 4368 15736 4368 0 net30
rlabel metal2 16072 5712 16072 5712 0 net31
rlabel metal2 8848 3416 8848 3416 0 net32
rlabel metal2 10808 5040 10808 5040 0 net33
rlabel metal2 14056 5040 14056 5040 0 net34
rlabel metal2 15624 4760 15624 4760 0 net35
rlabel metal2 6160 4424 6160 4424 0 net36
rlabel metal3 8120 3416 8120 3416 0 net37
rlabel metal2 6776 4144 6776 4144 0 net38
rlabel metal2 5712 6552 5712 6552 0 net39
rlabel metal2 9912 4200 9912 4200 0 net4
rlabel metal2 5320 4256 5320 4256 0 net40
rlabel metal2 37688 3360 37688 3360 0 net41
rlabel metal2 28168 45640 28168 45640 0 net42
rlabel metal2 37352 45640 37352 45640 0 net43
rlabel metal2 1736 3864 1736 3864 0 net44
rlabel metal2 2632 5936 2632 5936 0 net45
rlabel metal2 4312 7280 4312 7280 0 net46
rlabel metal3 2296 44968 2296 44968 0 net47
rlabel metal2 14000 45864 14000 45864 0 net48
rlabel metal2 38248 18816 38248 18816 0 net49
rlabel metal2 16464 3416 16464 3416 0 net5
rlabel metal2 22568 45752 22568 45752 0 net50
rlabel metal2 32424 45752 32424 45752 0 net51
rlabel metal3 1246 8120 1246 8120 0 net52
rlabel metal3 1246 9464 1246 9464 0 net53
rlabel metal3 1246 10808 1246 10808 0 net54
rlabel metal3 1246 12152 1246 12152 0 net55
rlabel metal3 1246 13496 1246 13496 0 net56
rlabel metal3 1246 14840 1246 14840 0 net57
rlabel metal3 1246 16184 1246 16184 0 net58
rlabel metal3 1246 17528 1246 17528 0 net59
rlabel metal2 16968 3416 16968 3416 0 net6
rlabel metal3 1246 18872 1246 18872 0 net60
rlabel metal3 1246 20216 1246 20216 0 net61
rlabel metal3 1246 21560 1246 21560 0 net62
rlabel metal3 1246 22904 1246 22904 0 net63
rlabel metal3 1246 24248 1246 24248 0 net64
rlabel metal3 1246 25592 1246 25592 0 net65
rlabel metal2 1736 26880 1736 26880 0 net66
rlabel metal3 1246 28280 1246 28280 0 net67
rlabel metal3 1246 29624 1246 29624 0 net68
rlabel metal3 1246 30968 1246 30968 0 net69
rlabel metal2 18312 3864 18312 3864 0 net7
rlabel metal3 1246 32312 1246 32312 0 net70
rlabel metal3 1246 33656 1246 33656 0 net71
rlabel metal3 1246 35000 1246 35000 0 net72
rlabel metal3 1246 36344 1246 36344 0 net73
rlabel metal3 1246 37688 1246 37688 0 net74
rlabel metal3 1246 39032 1246 39032 0 net75
rlabel metal3 1246 40376 1246 40376 0 net76
rlabel metal3 1246 41720 1246 41720 0 net77
rlabel metal3 1246 43064 1246 43064 0 net78
rlabel metal3 1246 44408 1246 44408 0 net79
rlabel metal2 19208 3920 19208 3920 0 net8
rlabel metal2 2184 45528 2184 45528 0 net80
rlabel metal2 2072 46368 2072 46368 0 net81
rlabel metal3 1246 4088 1246 4088 0 net82
rlabel metal2 7784 45752 7784 45752 0 net83
rlabel metal2 17640 45752 17640 45752 0 net84
rlabel metal3 38738 43288 38738 43288 0 net85
rlabel metal2 20104 3920 20104 3920 0 net9
rlabel metal3 1470 2744 1470 2744 0 o_wb_ack
rlabel metal3 1470 5432 1470 5432 0 o_wb_data[0]
rlabel metal3 1358 6776 1358 6776 0 o_wb_data[1]
rlabel metal2 37912 3024 37912 3024 0 reset
rlabel metal2 2744 47642 2744 47642 0 xtal_clk_enb[0]
rlabel metal3 13104 45976 13104 45976 0 xtal_clk_enb[1]
<< properties >>
string FIXED_BBOX 0 0 40000 50000
<< end >>
