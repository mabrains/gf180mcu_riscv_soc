module mabrains_logo ();
endmodule
