VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO pinmux_top
  CLASS BLOCK ;
  FOREIGN pinmux_top ;
  ORIGIN 0.000 0.000 ;
  SIZE 900.000 BY 1000.000 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 15.380 331.040 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 483.040 15.380 484.640 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 636.640 15.380 638.240 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 790.240 15.380 791.840 984.220 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 406.240 15.380 407.840 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 559.840 15.380 561.440 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 713.440 15.380 715.040 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 867.040 15.380 868.640 984.220 ;
    END
  END VSS
  PIN digital_io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 31.360 900.000 31.920 ;
    END
  END digital_io_in[0]
  PIN digital_io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 669.760 900.000 670.320 ;
    END
  END digital_io_in[10]
  PIN digital_io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 733.600 900.000 734.160 ;
    END
  END digital_io_in[11]
  PIN digital_io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 797.440 900.000 798.000 ;
    END
  END digital_io_in[12]
  PIN digital_io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 861.280 900.000 861.840 ;
    END
  END digital_io_in[13]
  PIN digital_io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 925.120 900.000 925.680 ;
    END
  END digital_io_in[14]
  PIN digital_io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 863.520 996.000 864.080 1000.000 ;
    END
  END digital_io_in[15]
  PIN digital_io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 846.720 996.000 847.280 1000.000 ;
    END
  END digital_io_in[16]
  PIN digital_io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 829.920 996.000 830.480 1000.000 ;
    END
  END digital_io_in[17]
  PIN digital_io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 813.120 996.000 813.680 1000.000 ;
    END
  END digital_io_in[18]
  PIN digital_io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 796.320 996.000 796.880 1000.000 ;
    END
  END digital_io_in[19]
  PIN digital_io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 95.200 900.000 95.760 ;
    END
  END digital_io_in[1]
  PIN digital_io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 779.520 996.000 780.080 1000.000 ;
    END
  END digital_io_in[20]
  PIN digital_io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 762.720 996.000 763.280 1000.000 ;
    END
  END digital_io_in[21]
  PIN digital_io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 745.920 996.000 746.480 1000.000 ;
    END
  END digital_io_in[22]
  PIN digital_io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 729.120 996.000 729.680 1000.000 ;
    END
  END digital_io_in[23]
  PIN digital_io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 253.120 996.000 253.680 1000.000 ;
    END
  END digital_io_in[24]
  PIN digital_io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 236.320 996.000 236.880 1000.000 ;
    END
  END digital_io_in[25]
  PIN digital_io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 219.520 996.000 220.080 1000.000 ;
    END
  END digital_io_in[26]
  PIN digital_io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 202.720 996.000 203.280 1000.000 ;
    END
  END digital_io_in[27]
  PIN digital_io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 185.920 996.000 186.480 1000.000 ;
    END
  END digital_io_in[28]
  PIN digital_io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 169.120 996.000 169.680 1000.000 ;
    END
  END digital_io_in[29]
  PIN digital_io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 159.040 900.000 159.600 ;
    END
  END digital_io_in[2]
  PIN digital_io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 152.320 996.000 152.880 1000.000 ;
    END
  END digital_io_in[30]
  PIN digital_io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 135.520 996.000 136.080 1000.000 ;
    END
  END digital_io_in[31]
  PIN digital_io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 118.720 996.000 119.280 1000.000 ;
    END
  END digital_io_in[32]
  PIN digital_io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 101.920 996.000 102.480 1000.000 ;
    END
  END digital_io_in[33]
  PIN digital_io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 85.120 996.000 85.680 1000.000 ;
    END
  END digital_io_in[34]
  PIN digital_io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 68.320 996.000 68.880 1000.000 ;
    END
  END digital_io_in[35]
  PIN digital_io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 51.520 996.000 52.080 1000.000 ;
    END
  END digital_io_in[36]
  PIN digital_io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 34.720 996.000 35.280 1000.000 ;
    END
  END digital_io_in[37]
  PIN digital_io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 222.880 900.000 223.440 ;
    END
  END digital_io_in[3]
  PIN digital_io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 286.720 900.000 287.280 ;
    END
  END digital_io_in[4]
  PIN digital_io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 350.560 900.000 351.120 ;
    END
  END digital_io_in[5]
  PIN digital_io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 414.400 900.000 414.960 ;
    END
  END digital_io_in[6]
  PIN digital_io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 478.240 900.000 478.800 ;
    END
  END digital_io_in[7]
  PIN digital_io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 542.080 900.000 542.640 ;
    END
  END digital_io_in[8]
  PIN digital_io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 605.920 900.000 606.480 ;
    END
  END digital_io_in[9]
  PIN digital_io_oen[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 73.920 900.000 74.480 ;
    END
  END digital_io_oen[0]
  PIN digital_io_oen[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 712.320 900.000 712.880 ;
    END
  END digital_io_oen[10]
  PIN digital_io_oen[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 776.160 900.000 776.720 ;
    END
  END digital_io_oen[11]
  PIN digital_io_oen[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 840.000 900.000 840.560 ;
    END
  END digital_io_oen[12]
  PIN digital_io_oen[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 903.840 900.000 904.400 ;
    END
  END digital_io_oen[13]
  PIN digital_io_oen[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 967.680 900.000 968.240 ;
    END
  END digital_io_oen[14]
  PIN digital_io_oen[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 874.720 996.000 875.280 1000.000 ;
    END
  END digital_io_oen[15]
  PIN digital_io_oen[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 857.920 996.000 858.480 1000.000 ;
    END
  END digital_io_oen[16]
  PIN digital_io_oen[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 841.120 996.000 841.680 1000.000 ;
    END
  END digital_io_oen[17]
  PIN digital_io_oen[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 824.320 996.000 824.880 1000.000 ;
    END
  END digital_io_oen[18]
  PIN digital_io_oen[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 807.520 996.000 808.080 1000.000 ;
    END
  END digital_io_oen[19]
  PIN digital_io_oen[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 137.760 900.000 138.320 ;
    END
  END digital_io_oen[1]
  PIN digital_io_oen[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 790.720 996.000 791.280 1000.000 ;
    END
  END digital_io_oen[20]
  PIN digital_io_oen[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 773.920 996.000 774.480 1000.000 ;
    END
  END digital_io_oen[21]
  PIN digital_io_oen[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 757.120 996.000 757.680 1000.000 ;
    END
  END digital_io_oen[22]
  PIN digital_io_oen[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 740.320 996.000 740.880 1000.000 ;
    END
  END digital_io_oen[23]
  PIN digital_io_oen[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 241.920 996.000 242.480 1000.000 ;
    END
  END digital_io_oen[24]
  PIN digital_io_oen[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 225.120 996.000 225.680 1000.000 ;
    END
  END digital_io_oen[25]
  PIN digital_io_oen[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 208.320 996.000 208.880 1000.000 ;
    END
  END digital_io_oen[26]
  PIN digital_io_oen[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 191.520 996.000 192.080 1000.000 ;
    END
  END digital_io_oen[27]
  PIN digital_io_oen[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 174.720 996.000 175.280 1000.000 ;
    END
  END digital_io_oen[28]
  PIN digital_io_oen[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 157.920 996.000 158.480 1000.000 ;
    END
  END digital_io_oen[29]
  PIN digital_io_oen[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 201.600 900.000 202.160 ;
    END
  END digital_io_oen[2]
  PIN digital_io_oen[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 141.120 996.000 141.680 1000.000 ;
    END
  END digital_io_oen[30]
  PIN digital_io_oen[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 124.320 996.000 124.880 1000.000 ;
    END
  END digital_io_oen[31]
  PIN digital_io_oen[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 107.520 996.000 108.080 1000.000 ;
    END
  END digital_io_oen[32]
  PIN digital_io_oen[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 90.720 996.000 91.280 1000.000 ;
    END
  END digital_io_oen[33]
  PIN digital_io_oen[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 73.920 996.000 74.480 1000.000 ;
    END
  END digital_io_oen[34]
  PIN digital_io_oen[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 57.120 996.000 57.680 1000.000 ;
    END
  END digital_io_oen[35]
  PIN digital_io_oen[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 40.320 996.000 40.880 1000.000 ;
    END
  END digital_io_oen[36]
  PIN digital_io_oen[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 23.520 996.000 24.080 1000.000 ;
    END
  END digital_io_oen[37]
  PIN digital_io_oen[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 265.440 900.000 266.000 ;
    END
  END digital_io_oen[3]
  PIN digital_io_oen[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 329.280 900.000 329.840 ;
    END
  END digital_io_oen[4]
  PIN digital_io_oen[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 393.120 900.000 393.680 ;
    END
  END digital_io_oen[5]
  PIN digital_io_oen[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 456.960 900.000 457.520 ;
    END
  END digital_io_oen[6]
  PIN digital_io_oen[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 520.800 900.000 521.360 ;
    END
  END digital_io_oen[7]
  PIN digital_io_oen[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 584.640 900.000 585.200 ;
    END
  END digital_io_oen[8]
  PIN digital_io_oen[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 648.480 900.000 649.040 ;
    END
  END digital_io_oen[9]
  PIN digital_io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 52.640 900.000 53.200 ;
    END
  END digital_io_out[0]
  PIN digital_io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 691.040 900.000 691.600 ;
    END
  END digital_io_out[10]
  PIN digital_io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 754.880 900.000 755.440 ;
    END
  END digital_io_out[11]
  PIN digital_io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 818.720 900.000 819.280 ;
    END
  END digital_io_out[12]
  PIN digital_io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 882.560 900.000 883.120 ;
    END
  END digital_io_out[13]
  PIN digital_io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 946.400 900.000 946.960 ;
    END
  END digital_io_out[14]
  PIN digital_io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 869.120 996.000 869.680 1000.000 ;
    END
  END digital_io_out[15]
  PIN digital_io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 852.320 996.000 852.880 1000.000 ;
    END
  END digital_io_out[16]
  PIN digital_io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 835.520 996.000 836.080 1000.000 ;
    END
  END digital_io_out[17]
  PIN digital_io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 818.720 996.000 819.280 1000.000 ;
    END
  END digital_io_out[18]
  PIN digital_io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 801.920 996.000 802.480 1000.000 ;
    END
  END digital_io_out[19]
  PIN digital_io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 116.480 900.000 117.040 ;
    END
  END digital_io_out[1]
  PIN digital_io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 785.120 996.000 785.680 1000.000 ;
    END
  END digital_io_out[20]
  PIN digital_io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 768.320 996.000 768.880 1000.000 ;
    END
  END digital_io_out[21]
  PIN digital_io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 751.520 996.000 752.080 1000.000 ;
    END
  END digital_io_out[22]
  PIN digital_io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 734.720 996.000 735.280 1000.000 ;
    END
  END digital_io_out[23]
  PIN digital_io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 247.520 996.000 248.080 1000.000 ;
    END
  END digital_io_out[24]
  PIN digital_io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 230.720 996.000 231.280 1000.000 ;
    END
  END digital_io_out[25]
  PIN digital_io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 213.920 996.000 214.480 1000.000 ;
    END
  END digital_io_out[26]
  PIN digital_io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 197.120 996.000 197.680 1000.000 ;
    END
  END digital_io_out[27]
  PIN digital_io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 180.320 996.000 180.880 1000.000 ;
    END
  END digital_io_out[28]
  PIN digital_io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 163.520 996.000 164.080 1000.000 ;
    END
  END digital_io_out[29]
  PIN digital_io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 180.320 900.000 180.880 ;
    END
  END digital_io_out[2]
  PIN digital_io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 146.720 996.000 147.280 1000.000 ;
    END
  END digital_io_out[30]
  PIN digital_io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 129.920 996.000 130.480 1000.000 ;
    END
  END digital_io_out[31]
  PIN digital_io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 113.120 996.000 113.680 1000.000 ;
    END
  END digital_io_out[32]
  PIN digital_io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 96.320 996.000 96.880 1000.000 ;
    END
  END digital_io_out[33]
  PIN digital_io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 79.520 996.000 80.080 1000.000 ;
    END
  END digital_io_out[34]
  PIN digital_io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 62.720 996.000 63.280 1000.000 ;
    END
  END digital_io_out[35]
  PIN digital_io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 45.920 996.000 46.480 1000.000 ;
    END
  END digital_io_out[36]
  PIN digital_io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 29.120 996.000 29.680 1000.000 ;
    END
  END digital_io_out[37]
  PIN digital_io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 244.160 900.000 244.720 ;
    END
  END digital_io_out[3]
  PIN digital_io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 308.000 900.000 308.560 ;
    END
  END digital_io_out[4]
  PIN digital_io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 371.840 900.000 372.400 ;
    END
  END digital_io_out[5]
  PIN digital_io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 435.680 900.000 436.240 ;
    END
  END digital_io_out[6]
  PIN digital_io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 499.520 900.000 500.080 ;
    END
  END digital_io_out[7]
  PIN digital_io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 563.360 900.000 563.920 ;
    END
  END digital_io_out[8]
  PIN digital_io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 627.200 900.000 627.760 ;
    END
  END digital_io_out[9]
  PIN e_reset_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 40.320 4.000 40.880 ;
    END
  END e_reset_n
  PIN i2cm_clk_i
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 437.920 0.000 438.480 4.000 ;
    END
  END i2cm_clk_i
  PIN i2cm_clk_o
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 414.400 0.000 414.960 4.000 ;
    END
  END i2cm_clk_o
  PIN i2cm_clk_oen
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 461.440 0.000 462.000 4.000 ;
    END
  END i2cm_clk_oen
  PIN i2cm_data_i
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 532.000 0.000 532.560 4.000 ;
    END
  END i2cm_data_i
  PIN i2cm_data_o
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 508.480 0.000 509.040 4.000 ;
    END
  END i2cm_data_o
  PIN i2cm_data_oen
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 484.960 0.000 485.520 4.000 ;
    END
  END i2cm_data_oen
  PIN i2cm_intr
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 743.680 0.000 744.240 4.000 ;
    END
  END i2cm_intr
  PIN i2cm_rst_n
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 85.120 0.000 85.680 4.000 ;
    END
  END i2cm_rst_n
  PIN mclk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 51.520 4.000 52.080 ;
    END
  END mclk
  PIN p_reset_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 29.120 4.000 29.680 ;
    END
  END p_reset_n
  PIN pulse1m_mclk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 720.160 0.000 720.720 4.000 ;
    END
  END pulse1m_mclk
  PIN reg_ack
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 969.920 4.000 970.480 ;
    END
  END reg_ack
  PIN reg_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 197.120 4.000 197.680 ;
    END
  END reg_addr[0]
  PIN reg_addr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.408000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 85.120 4.000 85.680 ;
    END
  END reg_addr[10]
  PIN reg_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 185.920 4.000 186.480 ;
    END
  END reg_addr[1]
  PIN reg_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 174.720 4.000 175.280 ;
    END
  END reg_addr[2]
  PIN reg_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 163.520 4.000 164.080 ;
    END
  END reg_addr[3]
  PIN reg_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 152.320 4.000 152.880 ;
    END
  END reg_addr[4]
  PIN reg_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 141.120 4.000 141.680 ;
    END
  END reg_addr[5]
  PIN reg_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 129.920 4.000 130.480 ;
    END
  END reg_addr[6]
  PIN reg_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 118.720 4.000 119.280 ;
    END
  END reg_addr[7]
  PIN reg_addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 107.520 4.000 108.080 ;
    END
  END reg_addr[8]
  PIN reg_addr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.408000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 96.320 4.000 96.880 ;
    END
  END reg_addr[9]
  PIN reg_be[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.408000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 241.920 4.000 242.480 ;
    END
  END reg_be[0]
  PIN reg_be[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 230.720 4.000 231.280 ;
    END
  END reg_be[1]
  PIN reg_be[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 219.520 4.000 220.080 ;
    END
  END reg_be[2]
  PIN reg_be[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 208.320 4.000 208.880 ;
    END
  END reg_be[3]
  PIN reg_cs
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 62.720 4.000 63.280 ;
    END
  END reg_cs
  PIN reg_peri_ack
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 723.520 996.000 724.080 1000.000 ;
    END
  END reg_peri_ack
  PIN reg_peri_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 337.120 996.000 337.680 1000.000 ;
    END
  END reg_peri_addr[0]
  PIN reg_peri_addr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 281.120 996.000 281.680 1000.000 ;
    END
  END reg_peri_addr[10]
  PIN reg_peri_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 331.520 996.000 332.080 1000.000 ;
    END
  END reg_peri_addr[1]
  PIN reg_peri_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 325.920 996.000 326.480 1000.000 ;
    END
  END reg_peri_addr[2]
  PIN reg_peri_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 320.320 996.000 320.880 1000.000 ;
    END
  END reg_peri_addr[3]
  PIN reg_peri_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 314.720 996.000 315.280 1000.000 ;
    END
  END reg_peri_addr[4]
  PIN reg_peri_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 309.120 996.000 309.680 1000.000 ;
    END
  END reg_peri_addr[5]
  PIN reg_peri_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 303.520 996.000 304.080 1000.000 ;
    END
  END reg_peri_addr[6]
  PIN reg_peri_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 297.920 996.000 298.480 1000.000 ;
    END
  END reg_peri_addr[7]
  PIN reg_peri_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 292.320 996.000 292.880 1000.000 ;
    END
  END reg_peri_addr[8]
  PIN reg_peri_addr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 286.720 996.000 287.280 1000.000 ;
    END
  END reg_peri_addr[9]
  PIN reg_peri_be[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 359.520 996.000 360.080 1000.000 ;
    END
  END reg_peri_be[0]
  PIN reg_peri_be[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 353.920 996.000 354.480 1000.000 ;
    END
  END reg_peri_be[1]
  PIN reg_peri_be[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 348.320 996.000 348.880 1000.000 ;
    END
  END reg_peri_be[2]
  PIN reg_peri_be[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 342.720 996.000 343.280 1000.000 ;
    END
  END reg_peri_be[3]
  PIN reg_peri_cs
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 269.920 996.000 270.480 1000.000 ;
    END
  END reg_peri_cs
  PIN reg_peri_rdata[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 717.920 996.000 718.480 1000.000 ;
    END
  END reg_peri_rdata[0]
  PIN reg_peri_rdata[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 661.920 996.000 662.480 1000.000 ;
    END
  END reg_peri_rdata[10]
  PIN reg_peri_rdata[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 656.320 996.000 656.880 1000.000 ;
    END
  END reg_peri_rdata[11]
  PIN reg_peri_rdata[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 650.720 996.000 651.280 1000.000 ;
    END
  END reg_peri_rdata[12]
  PIN reg_peri_rdata[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 645.120 996.000 645.680 1000.000 ;
    END
  END reg_peri_rdata[13]
  PIN reg_peri_rdata[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 639.520 996.000 640.080 1000.000 ;
    END
  END reg_peri_rdata[14]
  PIN reg_peri_rdata[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 633.920 996.000 634.480 1000.000 ;
    END
  END reg_peri_rdata[15]
  PIN reg_peri_rdata[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 628.320 996.000 628.880 1000.000 ;
    END
  END reg_peri_rdata[16]
  PIN reg_peri_rdata[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 622.720 996.000 623.280 1000.000 ;
    END
  END reg_peri_rdata[17]
  PIN reg_peri_rdata[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 617.120 996.000 617.680 1000.000 ;
    END
  END reg_peri_rdata[18]
  PIN reg_peri_rdata[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 611.520 996.000 612.080 1000.000 ;
    END
  END reg_peri_rdata[19]
  PIN reg_peri_rdata[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 712.320 996.000 712.880 1000.000 ;
    END
  END reg_peri_rdata[1]
  PIN reg_peri_rdata[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 605.920 996.000 606.480 1000.000 ;
    END
  END reg_peri_rdata[20]
  PIN reg_peri_rdata[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 600.320 996.000 600.880 1000.000 ;
    END
  END reg_peri_rdata[21]
  PIN reg_peri_rdata[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 594.720 996.000 595.280 1000.000 ;
    END
  END reg_peri_rdata[22]
  PIN reg_peri_rdata[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 589.120 996.000 589.680 1000.000 ;
    END
  END reg_peri_rdata[23]
  PIN reg_peri_rdata[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 583.520 996.000 584.080 1000.000 ;
    END
  END reg_peri_rdata[24]
  PIN reg_peri_rdata[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 577.920 996.000 578.480 1000.000 ;
    END
  END reg_peri_rdata[25]
  PIN reg_peri_rdata[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 572.320 996.000 572.880 1000.000 ;
    END
  END reg_peri_rdata[26]
  PIN reg_peri_rdata[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 566.720 996.000 567.280 1000.000 ;
    END
  END reg_peri_rdata[27]
  PIN reg_peri_rdata[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 561.120 996.000 561.680 1000.000 ;
    END
  END reg_peri_rdata[28]
  PIN reg_peri_rdata[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 555.520 996.000 556.080 1000.000 ;
    END
  END reg_peri_rdata[29]
  PIN reg_peri_rdata[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 706.720 996.000 707.280 1000.000 ;
    END
  END reg_peri_rdata[2]
  PIN reg_peri_rdata[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 549.920 996.000 550.480 1000.000 ;
    END
  END reg_peri_rdata[30]
  PIN reg_peri_rdata[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 544.320 996.000 544.880 1000.000 ;
    END
  END reg_peri_rdata[31]
  PIN reg_peri_rdata[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 701.120 996.000 701.680 1000.000 ;
    END
  END reg_peri_rdata[3]
  PIN reg_peri_rdata[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 695.520 996.000 696.080 1000.000 ;
    END
  END reg_peri_rdata[4]
  PIN reg_peri_rdata[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 689.920 996.000 690.480 1000.000 ;
    END
  END reg_peri_rdata[5]
  PIN reg_peri_rdata[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 684.320 996.000 684.880 1000.000 ;
    END
  END reg_peri_rdata[6]
  PIN reg_peri_rdata[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 678.720 996.000 679.280 1000.000 ;
    END
  END reg_peri_rdata[7]
  PIN reg_peri_rdata[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 673.120 996.000 673.680 1000.000 ;
    END
  END reg_peri_rdata[8]
  PIN reg_peri_rdata[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 667.520 996.000 668.080 1000.000 ;
    END
  END reg_peri_rdata[9]
  PIN reg_peri_wdata[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 538.720 996.000 539.280 1000.000 ;
    END
  END reg_peri_wdata[0]
  PIN reg_peri_wdata[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 482.720 996.000 483.280 1000.000 ;
    END
  END reg_peri_wdata[10]
  PIN reg_peri_wdata[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 477.120 996.000 477.680 1000.000 ;
    END
  END reg_peri_wdata[11]
  PIN reg_peri_wdata[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 471.520 996.000 472.080 1000.000 ;
    END
  END reg_peri_wdata[12]
  PIN reg_peri_wdata[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 465.920 996.000 466.480 1000.000 ;
    END
  END reg_peri_wdata[13]
  PIN reg_peri_wdata[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 460.320 996.000 460.880 1000.000 ;
    END
  END reg_peri_wdata[14]
  PIN reg_peri_wdata[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 454.720 996.000 455.280 1000.000 ;
    END
  END reg_peri_wdata[15]
  PIN reg_peri_wdata[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal2 ;
        RECT 449.120 996.000 449.680 1000.000 ;
    END
  END reg_peri_wdata[16]
  PIN reg_peri_wdata[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 443.520 996.000 444.080 1000.000 ;
    END
  END reg_peri_wdata[17]
  PIN reg_peri_wdata[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 437.920 996.000 438.480 1000.000 ;
    END
  END reg_peri_wdata[18]
  PIN reg_peri_wdata[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 432.320 996.000 432.880 1000.000 ;
    END
  END reg_peri_wdata[19]
  PIN reg_peri_wdata[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 533.120 996.000 533.680 1000.000 ;
    END
  END reg_peri_wdata[1]
  PIN reg_peri_wdata[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 426.720 996.000 427.280 1000.000 ;
    END
  END reg_peri_wdata[20]
  PIN reg_peri_wdata[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 421.120 996.000 421.680 1000.000 ;
    END
  END reg_peri_wdata[21]
  PIN reg_peri_wdata[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal2 ;
        RECT 415.520 996.000 416.080 1000.000 ;
    END
  END reg_peri_wdata[22]
  PIN reg_peri_wdata[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 409.920 996.000 410.480 1000.000 ;
    END
  END reg_peri_wdata[23]
  PIN reg_peri_wdata[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 404.320 996.000 404.880 1000.000 ;
    END
  END reg_peri_wdata[24]
  PIN reg_peri_wdata[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 398.720 996.000 399.280 1000.000 ;
    END
  END reg_peri_wdata[25]
  PIN reg_peri_wdata[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 393.120 996.000 393.680 1000.000 ;
    END
  END reg_peri_wdata[26]
  PIN reg_peri_wdata[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 387.520 996.000 388.080 1000.000 ;
    END
  END reg_peri_wdata[27]
  PIN reg_peri_wdata[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 381.920 996.000 382.480 1000.000 ;
    END
  END reg_peri_wdata[28]
  PIN reg_peri_wdata[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 376.320 996.000 376.880 1000.000 ;
    END
  END reg_peri_wdata[29]
  PIN reg_peri_wdata[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 527.520 996.000 528.080 1000.000 ;
    END
  END reg_peri_wdata[2]
  PIN reg_peri_wdata[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 370.720 996.000 371.280 1000.000 ;
    END
  END reg_peri_wdata[30]
  PIN reg_peri_wdata[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 365.120 996.000 365.680 1000.000 ;
    END
  END reg_peri_wdata[31]
  PIN reg_peri_wdata[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 521.920 996.000 522.480 1000.000 ;
    END
  END reg_peri_wdata[3]
  PIN reg_peri_wdata[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 516.320 996.000 516.880 1000.000 ;
    END
  END reg_peri_wdata[4]
  PIN reg_peri_wdata[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 510.720 996.000 511.280 1000.000 ;
    END
  END reg_peri_wdata[5]
  PIN reg_peri_wdata[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 505.120 996.000 505.680 1000.000 ;
    END
  END reg_peri_wdata[6]
  PIN reg_peri_wdata[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 499.520 996.000 500.080 1000.000 ;
    END
  END reg_peri_wdata[7]
  PIN reg_peri_wdata[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 493.920 996.000 494.480 1000.000 ;
    END
  END reg_peri_wdata[8]
  PIN reg_peri_wdata[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 488.320 996.000 488.880 1000.000 ;
    END
  END reg_peri_wdata[9]
  PIN reg_peri_wr
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 275.520 996.000 276.080 1000.000 ;
    END
  END reg_peri_wr
  PIN reg_rdata[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 958.720 4.000 959.280 ;
    END
  END reg_rdata[0]
  PIN reg_rdata[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 846.720 4.000 847.280 ;
    END
  END reg_rdata[10]
  PIN reg_rdata[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 835.520 4.000 836.080 ;
    END
  END reg_rdata[11]
  PIN reg_rdata[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 824.320 4.000 824.880 ;
    END
  END reg_rdata[12]
  PIN reg_rdata[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 813.120 4.000 813.680 ;
    END
  END reg_rdata[13]
  PIN reg_rdata[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 801.920 4.000 802.480 ;
    END
  END reg_rdata[14]
  PIN reg_rdata[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 790.720 4.000 791.280 ;
    END
  END reg_rdata[15]
  PIN reg_rdata[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 779.520 4.000 780.080 ;
    END
  END reg_rdata[16]
  PIN reg_rdata[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 768.320 4.000 768.880 ;
    END
  END reg_rdata[17]
  PIN reg_rdata[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 757.120 4.000 757.680 ;
    END
  END reg_rdata[18]
  PIN reg_rdata[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 745.920 4.000 746.480 ;
    END
  END reg_rdata[19]
  PIN reg_rdata[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 947.520 4.000 948.080 ;
    END
  END reg_rdata[1]
  PIN reg_rdata[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 734.720 4.000 735.280 ;
    END
  END reg_rdata[20]
  PIN reg_rdata[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 723.520 4.000 724.080 ;
    END
  END reg_rdata[21]
  PIN reg_rdata[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 712.320 4.000 712.880 ;
    END
  END reg_rdata[22]
  PIN reg_rdata[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 701.120 4.000 701.680 ;
    END
  END reg_rdata[23]
  PIN reg_rdata[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 689.920 4.000 690.480 ;
    END
  END reg_rdata[24]
  PIN reg_rdata[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 678.720 4.000 679.280 ;
    END
  END reg_rdata[25]
  PIN reg_rdata[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 667.520 4.000 668.080 ;
    END
  END reg_rdata[26]
  PIN reg_rdata[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 656.320 4.000 656.880 ;
    END
  END reg_rdata[27]
  PIN reg_rdata[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 645.120 4.000 645.680 ;
    END
  END reg_rdata[28]
  PIN reg_rdata[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 633.920 4.000 634.480 ;
    END
  END reg_rdata[29]
  PIN reg_rdata[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 936.320 4.000 936.880 ;
    END
  END reg_rdata[2]
  PIN reg_rdata[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 622.720 4.000 623.280 ;
    END
  END reg_rdata[30]
  PIN reg_rdata[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 611.520 4.000 612.080 ;
    END
  END reg_rdata[31]
  PIN reg_rdata[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 925.120 4.000 925.680 ;
    END
  END reg_rdata[3]
  PIN reg_rdata[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 913.920 4.000 914.480 ;
    END
  END reg_rdata[4]
  PIN reg_rdata[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 902.720 4.000 903.280 ;
    END
  END reg_rdata[5]
  PIN reg_rdata[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 891.520 4.000 892.080 ;
    END
  END reg_rdata[6]
  PIN reg_rdata[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 880.320 4.000 880.880 ;
    END
  END reg_rdata[7]
  PIN reg_rdata[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 869.120 4.000 869.680 ;
    END
  END reg_rdata[8]
  PIN reg_rdata[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 857.920 4.000 858.480 ;
    END
  END reg_rdata[9]
  PIN reg_wdata[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 600.320 4.000 600.880 ;
    END
  END reg_wdata[0]
  PIN reg_wdata[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 488.320 4.000 488.880 ;
    END
  END reg_wdata[10]
  PIN reg_wdata[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 477.120 4.000 477.680 ;
    END
  END reg_wdata[11]
  PIN reg_wdata[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 465.920 4.000 466.480 ;
    END
  END reg_wdata[12]
  PIN reg_wdata[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 454.720 4.000 455.280 ;
    END
  END reg_wdata[13]
  PIN reg_wdata[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 443.520 4.000 444.080 ;
    END
  END reg_wdata[14]
  PIN reg_wdata[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 432.320 4.000 432.880 ;
    END
  END reg_wdata[15]
  PIN reg_wdata[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 421.120 4.000 421.680 ;
    END
  END reg_wdata[16]
  PIN reg_wdata[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 409.920 4.000 410.480 ;
    END
  END reg_wdata[17]
  PIN reg_wdata[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 398.720 4.000 399.280 ;
    END
  END reg_wdata[18]
  PIN reg_wdata[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 387.520 4.000 388.080 ;
    END
  END reg_wdata[19]
  PIN reg_wdata[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 589.120 4.000 589.680 ;
    END
  END reg_wdata[1]
  PIN reg_wdata[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 376.320 4.000 376.880 ;
    END
  END reg_wdata[20]
  PIN reg_wdata[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 365.120 4.000 365.680 ;
    END
  END reg_wdata[21]
  PIN reg_wdata[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 353.920 4.000 354.480 ;
    END
  END reg_wdata[22]
  PIN reg_wdata[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 342.720 4.000 343.280 ;
    END
  END reg_wdata[23]
  PIN reg_wdata[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 331.520 4.000 332.080 ;
    END
  END reg_wdata[24]
  PIN reg_wdata[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 320.320 4.000 320.880 ;
    END
  END reg_wdata[25]
  PIN reg_wdata[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 309.120 4.000 309.680 ;
    END
  END reg_wdata[26]
  PIN reg_wdata[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 297.920 4.000 298.480 ;
    END
  END reg_wdata[27]
  PIN reg_wdata[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 286.720 4.000 287.280 ;
    END
  END reg_wdata[28]
  PIN reg_wdata[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 275.520 4.000 276.080 ;
    END
  END reg_wdata[29]
  PIN reg_wdata[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 577.920 4.000 578.480 ;
    END
  END reg_wdata[2]
  PIN reg_wdata[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 264.320 4.000 264.880 ;
    END
  END reg_wdata[30]
  PIN reg_wdata[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 253.120 4.000 253.680 ;
    END
  END reg_wdata[31]
  PIN reg_wdata[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 566.720 4.000 567.280 ;
    END
  END reg_wdata[3]
  PIN reg_wdata[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 555.520 4.000 556.080 ;
    END
  END reg_wdata[4]
  PIN reg_wdata[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 544.320 4.000 544.880 ;
    END
  END reg_wdata[5]
  PIN reg_wdata[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 533.120 4.000 533.680 ;
    END
  END reg_wdata[6]
  PIN reg_wdata[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 521.920 4.000 522.480 ;
    END
  END reg_wdata[7]
  PIN reg_wdata[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 510.720 4.000 511.280 ;
    END
  END reg_wdata[8]
  PIN reg_wdata[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 499.520 4.000 500.080 ;
    END
  END reg_wdata[9]
  PIN reg_wr
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 73.920 4.000 74.480 ;
    END
  END reg_wr
  PIN rtc_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 258.720 996.000 259.280 1000.000 ;
    END
  END rtc_clk
  PIN rtc_intr
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 264.320 996.000 264.880 1000.000 ;
    END
  END rtc_intr
  PIN s_reset_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 861.280 0.000 861.840 4.000 ;
    END
  END s_reset_n
  PIN spim_miso
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 673.120 0.000 673.680 4.000 ;
    END
  END spim_miso
  PIN spim_mosi
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 696.640 0.000 697.200 4.000 ;
    END
  END spim_mosi
  PIN spim_sck
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 555.520 0.000 556.080 4.000 ;
    END
  END spim_sck
  PIN spim_ssn[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 649.600 0.000 650.160 4.000 ;
    END
  END spim_ssn[0]
  PIN spim_ssn[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 626.080 0.000 626.640 4.000 ;
    END
  END spim_ssn[1]
  PIN spim_ssn[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 602.560 0.000 603.120 4.000 ;
    END
  END spim_ssn[2]
  PIN spim_ssn[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 579.040 0.000 579.600 4.000 ;
    END
  END spim_ssn[3]
  PIN sspim_rst_n
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 14.560 0.000 15.120 4.000 ;
    END
  END sspim_rst_n
  PIN uart_rst_n[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 61.600 0.000 62.160 4.000 ;
    END
  END uart_rst_n[0]
  PIN uart_rst_n[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 38.080 0.000 38.640 4.000 ;
    END
  END uart_rst_n[1]
  PIN uart_rxd[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 390.880 0.000 391.440 4.000 ;
    END
  END uart_rxd[0]
  PIN uart_rxd[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 343.840 0.000 344.400 4.000 ;
    END
  END uart_rxd[1]
  PIN uart_txd[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 367.360 0.000 367.920 4.000 ;
    END
  END uart_txd[0]
  PIN uart_txd[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 320.320 0.000 320.880 4.000 ;
    END
  END uart_txd[1]
  PIN usb_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 884.800 0.000 885.360 4.000 ;
    END
  END usb_clk
  PIN usb_dn_i
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 296.800 0.000 297.360 4.000 ;
    END
  END usb_dn_i
  PIN usb_dn_o
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 226.240 0.000 226.800 4.000 ;
    END
  END usb_dn_o
  PIN usb_dp_i
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 273.280 0.000 273.840 4.000 ;
    END
  END usb_dp_i
  PIN usb_dp_o
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 202.720 0.000 203.280 4.000 ;
    END
  END usb_dp_o
  PIN usb_intr
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 767.200 0.000 767.760 4.000 ;
    END
  END usb_intr
  PIN usb_oen
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 249.760 0.000 250.320 4.000 ;
    END
  END usb_oen
  PIN usb_rst_n
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 108.640 0.000 109.200 4.000 ;
    END
  END usb_rst_n
  PIN user_clock1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 790.720 0.000 791.280 4.000 ;
    END
  END user_clock1
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 814.240 0.000 814.800 4.000 ;
    END
  END user_clock2
  PIN user_irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 132.160 0.000 132.720 4.000 ;
    END
  END user_irq[0]
  PIN user_irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 155.680 0.000 156.240 4.000 ;
    END
  END user_irq[1]
  PIN user_irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 179.200 0.000 179.760 4.000 ;
    END
  END user_irq[2]
  PIN xtal_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 837.760 0.000 838.320 4.000 ;
    END
  END xtal_clk
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 893.200 989.370 ;
      LAYER Metal2 ;
        RECT 7.980 995.700 23.220 996.660 ;
        RECT 24.380 995.700 28.820 996.660 ;
        RECT 29.980 995.700 34.420 996.660 ;
        RECT 35.580 995.700 40.020 996.660 ;
        RECT 41.180 995.700 45.620 996.660 ;
        RECT 46.780 995.700 51.220 996.660 ;
        RECT 52.380 995.700 56.820 996.660 ;
        RECT 57.980 995.700 62.420 996.660 ;
        RECT 63.580 995.700 68.020 996.660 ;
        RECT 69.180 995.700 73.620 996.660 ;
        RECT 74.780 995.700 79.220 996.660 ;
        RECT 80.380 995.700 84.820 996.660 ;
        RECT 85.980 995.700 90.420 996.660 ;
        RECT 91.580 995.700 96.020 996.660 ;
        RECT 97.180 995.700 101.620 996.660 ;
        RECT 102.780 995.700 107.220 996.660 ;
        RECT 108.380 995.700 112.820 996.660 ;
        RECT 113.980 995.700 118.420 996.660 ;
        RECT 119.580 995.700 124.020 996.660 ;
        RECT 125.180 995.700 129.620 996.660 ;
        RECT 130.780 995.700 135.220 996.660 ;
        RECT 136.380 995.700 140.820 996.660 ;
        RECT 141.980 995.700 146.420 996.660 ;
        RECT 147.580 995.700 152.020 996.660 ;
        RECT 153.180 995.700 157.620 996.660 ;
        RECT 158.780 995.700 163.220 996.660 ;
        RECT 164.380 995.700 168.820 996.660 ;
        RECT 169.980 995.700 174.420 996.660 ;
        RECT 175.580 995.700 180.020 996.660 ;
        RECT 181.180 995.700 185.620 996.660 ;
        RECT 186.780 995.700 191.220 996.660 ;
        RECT 192.380 995.700 196.820 996.660 ;
        RECT 197.980 995.700 202.420 996.660 ;
        RECT 203.580 995.700 208.020 996.660 ;
        RECT 209.180 995.700 213.620 996.660 ;
        RECT 214.780 995.700 219.220 996.660 ;
        RECT 220.380 995.700 224.820 996.660 ;
        RECT 225.980 995.700 230.420 996.660 ;
        RECT 231.580 995.700 236.020 996.660 ;
        RECT 237.180 995.700 241.620 996.660 ;
        RECT 242.780 995.700 247.220 996.660 ;
        RECT 248.380 995.700 252.820 996.660 ;
        RECT 253.980 995.700 258.420 996.660 ;
        RECT 259.580 995.700 264.020 996.660 ;
        RECT 265.180 995.700 269.620 996.660 ;
        RECT 270.780 995.700 275.220 996.660 ;
        RECT 276.380 995.700 280.820 996.660 ;
        RECT 281.980 995.700 286.420 996.660 ;
        RECT 287.580 995.700 292.020 996.660 ;
        RECT 293.180 995.700 297.620 996.660 ;
        RECT 298.780 995.700 303.220 996.660 ;
        RECT 304.380 995.700 308.820 996.660 ;
        RECT 309.980 995.700 314.420 996.660 ;
        RECT 315.580 995.700 320.020 996.660 ;
        RECT 321.180 995.700 325.620 996.660 ;
        RECT 326.780 995.700 331.220 996.660 ;
        RECT 332.380 995.700 336.820 996.660 ;
        RECT 337.980 995.700 342.420 996.660 ;
        RECT 343.580 995.700 348.020 996.660 ;
        RECT 349.180 995.700 353.620 996.660 ;
        RECT 354.780 995.700 359.220 996.660 ;
        RECT 360.380 995.700 364.820 996.660 ;
        RECT 365.980 995.700 370.420 996.660 ;
        RECT 371.580 995.700 376.020 996.660 ;
        RECT 377.180 995.700 381.620 996.660 ;
        RECT 382.780 995.700 387.220 996.660 ;
        RECT 388.380 995.700 392.820 996.660 ;
        RECT 393.980 995.700 398.420 996.660 ;
        RECT 399.580 995.700 404.020 996.660 ;
        RECT 405.180 995.700 409.620 996.660 ;
        RECT 410.780 995.700 415.220 996.660 ;
        RECT 416.380 995.700 420.820 996.660 ;
        RECT 421.980 995.700 426.420 996.660 ;
        RECT 427.580 995.700 432.020 996.660 ;
        RECT 433.180 995.700 437.620 996.660 ;
        RECT 438.780 995.700 443.220 996.660 ;
        RECT 444.380 995.700 448.820 996.660 ;
        RECT 449.980 995.700 454.420 996.660 ;
        RECT 455.580 995.700 460.020 996.660 ;
        RECT 461.180 995.700 465.620 996.660 ;
        RECT 466.780 995.700 471.220 996.660 ;
        RECT 472.380 995.700 476.820 996.660 ;
        RECT 477.980 995.700 482.420 996.660 ;
        RECT 483.580 995.700 488.020 996.660 ;
        RECT 489.180 995.700 493.620 996.660 ;
        RECT 494.780 995.700 499.220 996.660 ;
        RECT 500.380 995.700 504.820 996.660 ;
        RECT 505.980 995.700 510.420 996.660 ;
        RECT 511.580 995.700 516.020 996.660 ;
        RECT 517.180 995.700 521.620 996.660 ;
        RECT 522.780 995.700 527.220 996.660 ;
        RECT 528.380 995.700 532.820 996.660 ;
        RECT 533.980 995.700 538.420 996.660 ;
        RECT 539.580 995.700 544.020 996.660 ;
        RECT 545.180 995.700 549.620 996.660 ;
        RECT 550.780 995.700 555.220 996.660 ;
        RECT 556.380 995.700 560.820 996.660 ;
        RECT 561.980 995.700 566.420 996.660 ;
        RECT 567.580 995.700 572.020 996.660 ;
        RECT 573.180 995.700 577.620 996.660 ;
        RECT 578.780 995.700 583.220 996.660 ;
        RECT 584.380 995.700 588.820 996.660 ;
        RECT 589.980 995.700 594.420 996.660 ;
        RECT 595.580 995.700 600.020 996.660 ;
        RECT 601.180 995.700 605.620 996.660 ;
        RECT 606.780 995.700 611.220 996.660 ;
        RECT 612.380 995.700 616.820 996.660 ;
        RECT 617.980 995.700 622.420 996.660 ;
        RECT 623.580 995.700 628.020 996.660 ;
        RECT 629.180 995.700 633.620 996.660 ;
        RECT 634.780 995.700 639.220 996.660 ;
        RECT 640.380 995.700 644.820 996.660 ;
        RECT 645.980 995.700 650.420 996.660 ;
        RECT 651.580 995.700 656.020 996.660 ;
        RECT 657.180 995.700 661.620 996.660 ;
        RECT 662.780 995.700 667.220 996.660 ;
        RECT 668.380 995.700 672.820 996.660 ;
        RECT 673.980 995.700 678.420 996.660 ;
        RECT 679.580 995.700 684.020 996.660 ;
        RECT 685.180 995.700 689.620 996.660 ;
        RECT 690.780 995.700 695.220 996.660 ;
        RECT 696.380 995.700 700.820 996.660 ;
        RECT 701.980 995.700 706.420 996.660 ;
        RECT 707.580 995.700 712.020 996.660 ;
        RECT 713.180 995.700 717.620 996.660 ;
        RECT 718.780 995.700 723.220 996.660 ;
        RECT 724.380 995.700 728.820 996.660 ;
        RECT 729.980 995.700 734.420 996.660 ;
        RECT 735.580 995.700 740.020 996.660 ;
        RECT 741.180 995.700 745.620 996.660 ;
        RECT 746.780 995.700 751.220 996.660 ;
        RECT 752.380 995.700 756.820 996.660 ;
        RECT 757.980 995.700 762.420 996.660 ;
        RECT 763.580 995.700 768.020 996.660 ;
        RECT 769.180 995.700 773.620 996.660 ;
        RECT 774.780 995.700 779.220 996.660 ;
        RECT 780.380 995.700 784.820 996.660 ;
        RECT 785.980 995.700 790.420 996.660 ;
        RECT 791.580 995.700 796.020 996.660 ;
        RECT 797.180 995.700 801.620 996.660 ;
        RECT 802.780 995.700 807.220 996.660 ;
        RECT 808.380 995.700 812.820 996.660 ;
        RECT 813.980 995.700 818.420 996.660 ;
        RECT 819.580 995.700 824.020 996.660 ;
        RECT 825.180 995.700 829.620 996.660 ;
        RECT 830.780 995.700 835.220 996.660 ;
        RECT 836.380 995.700 840.820 996.660 ;
        RECT 841.980 995.700 846.420 996.660 ;
        RECT 847.580 995.700 852.020 996.660 ;
        RECT 853.180 995.700 857.620 996.660 ;
        RECT 858.780 995.700 863.220 996.660 ;
        RECT 864.380 995.700 868.820 996.660 ;
        RECT 869.980 995.700 874.420 996.660 ;
        RECT 875.580 995.700 892.500 996.660 ;
        RECT 7.980 4.300 892.500 995.700 ;
        RECT 7.980 3.500 14.260 4.300 ;
        RECT 15.420 3.500 37.780 4.300 ;
        RECT 38.940 3.500 61.300 4.300 ;
        RECT 62.460 3.500 84.820 4.300 ;
        RECT 85.980 3.500 108.340 4.300 ;
        RECT 109.500 3.500 131.860 4.300 ;
        RECT 133.020 3.500 155.380 4.300 ;
        RECT 156.540 3.500 178.900 4.300 ;
        RECT 180.060 3.500 202.420 4.300 ;
        RECT 203.580 3.500 225.940 4.300 ;
        RECT 227.100 3.500 249.460 4.300 ;
        RECT 250.620 3.500 272.980 4.300 ;
        RECT 274.140 3.500 296.500 4.300 ;
        RECT 297.660 3.500 320.020 4.300 ;
        RECT 321.180 3.500 343.540 4.300 ;
        RECT 344.700 3.500 367.060 4.300 ;
        RECT 368.220 3.500 390.580 4.300 ;
        RECT 391.740 3.500 414.100 4.300 ;
        RECT 415.260 3.500 437.620 4.300 ;
        RECT 438.780 3.500 461.140 4.300 ;
        RECT 462.300 3.500 484.660 4.300 ;
        RECT 485.820 3.500 508.180 4.300 ;
        RECT 509.340 3.500 531.700 4.300 ;
        RECT 532.860 3.500 555.220 4.300 ;
        RECT 556.380 3.500 578.740 4.300 ;
        RECT 579.900 3.500 602.260 4.300 ;
        RECT 603.420 3.500 625.780 4.300 ;
        RECT 626.940 3.500 649.300 4.300 ;
        RECT 650.460 3.500 672.820 4.300 ;
        RECT 673.980 3.500 696.340 4.300 ;
        RECT 697.500 3.500 719.860 4.300 ;
        RECT 721.020 3.500 743.380 4.300 ;
        RECT 744.540 3.500 766.900 4.300 ;
        RECT 768.060 3.500 790.420 4.300 ;
        RECT 791.580 3.500 813.940 4.300 ;
        RECT 815.100 3.500 837.460 4.300 ;
        RECT 838.620 3.500 860.980 4.300 ;
        RECT 862.140 3.500 884.500 4.300 ;
        RECT 885.660 3.500 892.500 4.300 ;
      LAYER Metal3 ;
        RECT 4.000 970.780 896.000 984.060 ;
        RECT 4.300 969.620 896.000 970.780 ;
        RECT 4.000 968.540 896.000 969.620 ;
        RECT 4.000 967.380 895.700 968.540 ;
        RECT 4.000 959.580 896.000 967.380 ;
        RECT 4.300 958.420 896.000 959.580 ;
        RECT 4.000 948.380 896.000 958.420 ;
        RECT 4.300 947.260 896.000 948.380 ;
        RECT 4.300 947.220 895.700 947.260 ;
        RECT 4.000 946.100 895.700 947.220 ;
        RECT 4.000 937.180 896.000 946.100 ;
        RECT 4.300 936.020 896.000 937.180 ;
        RECT 4.000 925.980 896.000 936.020 ;
        RECT 4.300 924.820 895.700 925.980 ;
        RECT 4.000 914.780 896.000 924.820 ;
        RECT 4.300 913.620 896.000 914.780 ;
        RECT 4.000 904.700 896.000 913.620 ;
        RECT 4.000 903.580 895.700 904.700 ;
        RECT 4.300 903.540 895.700 903.580 ;
        RECT 4.300 902.420 896.000 903.540 ;
        RECT 4.000 892.380 896.000 902.420 ;
        RECT 4.300 891.220 896.000 892.380 ;
        RECT 4.000 883.420 896.000 891.220 ;
        RECT 4.000 882.260 895.700 883.420 ;
        RECT 4.000 881.180 896.000 882.260 ;
        RECT 4.300 880.020 896.000 881.180 ;
        RECT 4.000 869.980 896.000 880.020 ;
        RECT 4.300 868.820 896.000 869.980 ;
        RECT 4.000 862.140 896.000 868.820 ;
        RECT 4.000 860.980 895.700 862.140 ;
        RECT 4.000 858.780 896.000 860.980 ;
        RECT 4.300 857.620 896.000 858.780 ;
        RECT 4.000 847.580 896.000 857.620 ;
        RECT 4.300 846.420 896.000 847.580 ;
        RECT 4.000 840.860 896.000 846.420 ;
        RECT 4.000 839.700 895.700 840.860 ;
        RECT 4.000 836.380 896.000 839.700 ;
        RECT 4.300 835.220 896.000 836.380 ;
        RECT 4.000 825.180 896.000 835.220 ;
        RECT 4.300 824.020 896.000 825.180 ;
        RECT 4.000 819.580 896.000 824.020 ;
        RECT 4.000 818.420 895.700 819.580 ;
        RECT 4.000 813.980 896.000 818.420 ;
        RECT 4.300 812.820 896.000 813.980 ;
        RECT 4.000 802.780 896.000 812.820 ;
        RECT 4.300 801.620 896.000 802.780 ;
        RECT 4.000 798.300 896.000 801.620 ;
        RECT 4.000 797.140 895.700 798.300 ;
        RECT 4.000 791.580 896.000 797.140 ;
        RECT 4.300 790.420 896.000 791.580 ;
        RECT 4.000 780.380 896.000 790.420 ;
        RECT 4.300 779.220 896.000 780.380 ;
        RECT 4.000 777.020 896.000 779.220 ;
        RECT 4.000 775.860 895.700 777.020 ;
        RECT 4.000 769.180 896.000 775.860 ;
        RECT 4.300 768.020 896.000 769.180 ;
        RECT 4.000 757.980 896.000 768.020 ;
        RECT 4.300 756.820 896.000 757.980 ;
        RECT 4.000 755.740 896.000 756.820 ;
        RECT 4.000 754.580 895.700 755.740 ;
        RECT 4.000 746.780 896.000 754.580 ;
        RECT 4.300 745.620 896.000 746.780 ;
        RECT 4.000 735.580 896.000 745.620 ;
        RECT 4.300 734.460 896.000 735.580 ;
        RECT 4.300 734.420 895.700 734.460 ;
        RECT 4.000 733.300 895.700 734.420 ;
        RECT 4.000 724.380 896.000 733.300 ;
        RECT 4.300 723.220 896.000 724.380 ;
        RECT 4.000 713.180 896.000 723.220 ;
        RECT 4.300 712.020 895.700 713.180 ;
        RECT 4.000 701.980 896.000 712.020 ;
        RECT 4.300 700.820 896.000 701.980 ;
        RECT 4.000 691.900 896.000 700.820 ;
        RECT 4.000 690.780 895.700 691.900 ;
        RECT 4.300 690.740 895.700 690.780 ;
        RECT 4.300 689.620 896.000 690.740 ;
        RECT 4.000 679.580 896.000 689.620 ;
        RECT 4.300 678.420 896.000 679.580 ;
        RECT 4.000 670.620 896.000 678.420 ;
        RECT 4.000 669.460 895.700 670.620 ;
        RECT 4.000 668.380 896.000 669.460 ;
        RECT 4.300 667.220 896.000 668.380 ;
        RECT 4.000 657.180 896.000 667.220 ;
        RECT 4.300 656.020 896.000 657.180 ;
        RECT 4.000 649.340 896.000 656.020 ;
        RECT 4.000 648.180 895.700 649.340 ;
        RECT 4.000 645.980 896.000 648.180 ;
        RECT 4.300 644.820 896.000 645.980 ;
        RECT 4.000 634.780 896.000 644.820 ;
        RECT 4.300 633.620 896.000 634.780 ;
        RECT 4.000 628.060 896.000 633.620 ;
        RECT 4.000 626.900 895.700 628.060 ;
        RECT 4.000 623.580 896.000 626.900 ;
        RECT 4.300 622.420 896.000 623.580 ;
        RECT 4.000 612.380 896.000 622.420 ;
        RECT 4.300 611.220 896.000 612.380 ;
        RECT 4.000 606.780 896.000 611.220 ;
        RECT 4.000 605.620 895.700 606.780 ;
        RECT 4.000 601.180 896.000 605.620 ;
        RECT 4.300 600.020 896.000 601.180 ;
        RECT 4.000 589.980 896.000 600.020 ;
        RECT 4.300 588.820 896.000 589.980 ;
        RECT 4.000 585.500 896.000 588.820 ;
        RECT 4.000 584.340 895.700 585.500 ;
        RECT 4.000 578.780 896.000 584.340 ;
        RECT 4.300 577.620 896.000 578.780 ;
        RECT 4.000 567.580 896.000 577.620 ;
        RECT 4.300 566.420 896.000 567.580 ;
        RECT 4.000 564.220 896.000 566.420 ;
        RECT 4.000 563.060 895.700 564.220 ;
        RECT 4.000 556.380 896.000 563.060 ;
        RECT 4.300 555.220 896.000 556.380 ;
        RECT 4.000 545.180 896.000 555.220 ;
        RECT 4.300 544.020 896.000 545.180 ;
        RECT 4.000 542.940 896.000 544.020 ;
        RECT 4.000 541.780 895.700 542.940 ;
        RECT 4.000 533.980 896.000 541.780 ;
        RECT 4.300 532.820 896.000 533.980 ;
        RECT 4.000 522.780 896.000 532.820 ;
        RECT 4.300 521.660 896.000 522.780 ;
        RECT 4.300 521.620 895.700 521.660 ;
        RECT 4.000 520.500 895.700 521.620 ;
        RECT 4.000 511.580 896.000 520.500 ;
        RECT 4.300 510.420 896.000 511.580 ;
        RECT 4.000 500.380 896.000 510.420 ;
        RECT 4.300 499.220 895.700 500.380 ;
        RECT 4.000 489.180 896.000 499.220 ;
        RECT 4.300 488.020 896.000 489.180 ;
        RECT 4.000 479.100 896.000 488.020 ;
        RECT 4.000 477.980 895.700 479.100 ;
        RECT 4.300 477.940 895.700 477.980 ;
        RECT 4.300 476.820 896.000 477.940 ;
        RECT 4.000 466.780 896.000 476.820 ;
        RECT 4.300 465.620 896.000 466.780 ;
        RECT 4.000 457.820 896.000 465.620 ;
        RECT 4.000 456.660 895.700 457.820 ;
        RECT 4.000 455.580 896.000 456.660 ;
        RECT 4.300 454.420 896.000 455.580 ;
        RECT 4.000 444.380 896.000 454.420 ;
        RECT 4.300 443.220 896.000 444.380 ;
        RECT 4.000 436.540 896.000 443.220 ;
        RECT 4.000 435.380 895.700 436.540 ;
        RECT 4.000 433.180 896.000 435.380 ;
        RECT 4.300 432.020 896.000 433.180 ;
        RECT 4.000 421.980 896.000 432.020 ;
        RECT 4.300 420.820 896.000 421.980 ;
        RECT 4.000 415.260 896.000 420.820 ;
        RECT 4.000 414.100 895.700 415.260 ;
        RECT 4.000 410.780 896.000 414.100 ;
        RECT 4.300 409.620 896.000 410.780 ;
        RECT 4.000 399.580 896.000 409.620 ;
        RECT 4.300 398.420 896.000 399.580 ;
        RECT 4.000 393.980 896.000 398.420 ;
        RECT 4.000 392.820 895.700 393.980 ;
        RECT 4.000 388.380 896.000 392.820 ;
        RECT 4.300 387.220 896.000 388.380 ;
        RECT 4.000 377.180 896.000 387.220 ;
        RECT 4.300 376.020 896.000 377.180 ;
        RECT 4.000 372.700 896.000 376.020 ;
        RECT 4.000 371.540 895.700 372.700 ;
        RECT 4.000 365.980 896.000 371.540 ;
        RECT 4.300 364.820 896.000 365.980 ;
        RECT 4.000 354.780 896.000 364.820 ;
        RECT 4.300 353.620 896.000 354.780 ;
        RECT 4.000 351.420 896.000 353.620 ;
        RECT 4.000 350.260 895.700 351.420 ;
        RECT 4.000 343.580 896.000 350.260 ;
        RECT 4.300 342.420 896.000 343.580 ;
        RECT 4.000 332.380 896.000 342.420 ;
        RECT 4.300 331.220 896.000 332.380 ;
        RECT 4.000 330.140 896.000 331.220 ;
        RECT 4.000 328.980 895.700 330.140 ;
        RECT 4.000 321.180 896.000 328.980 ;
        RECT 4.300 320.020 896.000 321.180 ;
        RECT 4.000 309.980 896.000 320.020 ;
        RECT 4.300 308.860 896.000 309.980 ;
        RECT 4.300 308.820 895.700 308.860 ;
        RECT 4.000 307.700 895.700 308.820 ;
        RECT 4.000 298.780 896.000 307.700 ;
        RECT 4.300 297.620 896.000 298.780 ;
        RECT 4.000 287.580 896.000 297.620 ;
        RECT 4.300 286.420 895.700 287.580 ;
        RECT 4.000 276.380 896.000 286.420 ;
        RECT 4.300 275.220 896.000 276.380 ;
        RECT 4.000 266.300 896.000 275.220 ;
        RECT 4.000 265.180 895.700 266.300 ;
        RECT 4.300 265.140 895.700 265.180 ;
        RECT 4.300 264.020 896.000 265.140 ;
        RECT 4.000 253.980 896.000 264.020 ;
        RECT 4.300 252.820 896.000 253.980 ;
        RECT 4.000 245.020 896.000 252.820 ;
        RECT 4.000 243.860 895.700 245.020 ;
        RECT 4.000 242.780 896.000 243.860 ;
        RECT 4.300 241.620 896.000 242.780 ;
        RECT 4.000 231.580 896.000 241.620 ;
        RECT 4.300 230.420 896.000 231.580 ;
        RECT 4.000 223.740 896.000 230.420 ;
        RECT 4.000 222.580 895.700 223.740 ;
        RECT 4.000 220.380 896.000 222.580 ;
        RECT 4.300 219.220 896.000 220.380 ;
        RECT 4.000 209.180 896.000 219.220 ;
        RECT 4.300 208.020 896.000 209.180 ;
        RECT 4.000 202.460 896.000 208.020 ;
        RECT 4.000 201.300 895.700 202.460 ;
        RECT 4.000 197.980 896.000 201.300 ;
        RECT 4.300 196.820 896.000 197.980 ;
        RECT 4.000 186.780 896.000 196.820 ;
        RECT 4.300 185.620 896.000 186.780 ;
        RECT 4.000 181.180 896.000 185.620 ;
        RECT 4.000 180.020 895.700 181.180 ;
        RECT 4.000 175.580 896.000 180.020 ;
        RECT 4.300 174.420 896.000 175.580 ;
        RECT 4.000 164.380 896.000 174.420 ;
        RECT 4.300 163.220 896.000 164.380 ;
        RECT 4.000 159.900 896.000 163.220 ;
        RECT 4.000 158.740 895.700 159.900 ;
        RECT 4.000 153.180 896.000 158.740 ;
        RECT 4.300 152.020 896.000 153.180 ;
        RECT 4.000 141.980 896.000 152.020 ;
        RECT 4.300 140.820 896.000 141.980 ;
        RECT 4.000 138.620 896.000 140.820 ;
        RECT 4.000 137.460 895.700 138.620 ;
        RECT 4.000 130.780 896.000 137.460 ;
        RECT 4.300 129.620 896.000 130.780 ;
        RECT 4.000 119.580 896.000 129.620 ;
        RECT 4.300 118.420 896.000 119.580 ;
        RECT 4.000 117.340 896.000 118.420 ;
        RECT 4.000 116.180 895.700 117.340 ;
        RECT 4.000 108.380 896.000 116.180 ;
        RECT 4.300 107.220 896.000 108.380 ;
        RECT 4.000 97.180 896.000 107.220 ;
        RECT 4.300 96.060 896.000 97.180 ;
        RECT 4.300 96.020 895.700 96.060 ;
        RECT 4.000 94.900 895.700 96.020 ;
        RECT 4.000 85.980 896.000 94.900 ;
        RECT 4.300 84.820 896.000 85.980 ;
        RECT 4.000 74.780 896.000 84.820 ;
        RECT 4.300 73.620 895.700 74.780 ;
        RECT 4.000 63.580 896.000 73.620 ;
        RECT 4.300 62.420 896.000 63.580 ;
        RECT 4.000 53.500 896.000 62.420 ;
        RECT 4.000 52.380 895.700 53.500 ;
        RECT 4.300 52.340 895.700 52.380 ;
        RECT 4.300 51.220 896.000 52.340 ;
        RECT 4.000 41.180 896.000 51.220 ;
        RECT 4.300 40.020 896.000 41.180 ;
        RECT 4.000 32.220 896.000 40.020 ;
        RECT 4.000 31.060 895.700 32.220 ;
        RECT 4.000 29.980 896.000 31.060 ;
        RECT 4.300 28.820 896.000 29.980 ;
        RECT 4.000 15.540 896.000 28.820 ;
      LAYER Metal4 ;
        RECT 11.340 18.010 21.940 981.030 ;
        RECT 24.140 18.010 98.740 981.030 ;
        RECT 100.940 18.010 175.540 981.030 ;
        RECT 177.740 18.010 252.340 981.030 ;
        RECT 254.540 18.010 329.140 981.030 ;
        RECT 331.340 18.010 405.940 981.030 ;
        RECT 408.140 18.010 482.740 981.030 ;
        RECT 484.940 18.010 559.540 981.030 ;
        RECT 561.740 18.010 636.340 981.030 ;
        RECT 638.540 18.010 713.140 981.030 ;
        RECT 715.340 18.010 789.940 981.030 ;
        RECT 792.140 18.010 866.740 981.030 ;
        RECT 868.940 18.010 888.020 981.030 ;
      LAYER Metal5 ;
        RECT 11.260 130.730 860.100 978.070 ;
  END
END pinmux_top
END LIBRARY

