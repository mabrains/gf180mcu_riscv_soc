VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO uart_i2c_usb_spi_top
  CLASS BLOCK ;
  FOREIGN uart_i2c_usb_spi_top ;
  ORIGIN 0.000 0.000 ;
  SIZE 850.000 BY 1000.000 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 19.940 15.380 26.140 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 119.940 15.380 126.140 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 219.940 15.380 226.140 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 319.940 15.380 326.140 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 419.940 15.380 426.140 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 519.940 15.380 526.140 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 619.940 15.380 626.140 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 719.940 15.380 726.140 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 819.940 15.380 826.140 984.220 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 69.940 15.380 76.140 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 169.940 15.380 176.140 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 269.940 15.380 276.140 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 369.940 15.380 376.140 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 469.940 15.380 476.140 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 569.940 15.380 576.140 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 669.940 15.380 676.140 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 769.940 15.380 776.140 984.220 ;
    END
  END VSS
  PIN app_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 6.720 4.000 7.280 ;
    END
  END app_clk
  PIN i2c_rstn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 593.600 0.000 594.160 4.000 ;
    END
  END i2c_rstn
  PIN i2cm_intr_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 525.280 996.000 525.840 1000.000 ;
    END
  END i2cm_intr_o
  PIN reg_ack
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 992.320 4.000 992.880 ;
    END
  END reg_ack
  PIN reg_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 142.240 4.000 142.800 ;
    END
  END reg_addr[0]
  PIN reg_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 129.920 4.000 130.480 ;
    END
  END reg_addr[1]
  PIN reg_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 117.600 4.000 118.160 ;
    END
  END reg_addr[2]
  PIN reg_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 105.280 4.000 105.840 ;
    END
  END reg_addr[3]
  PIN reg_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 92.960 4.000 93.520 ;
    END
  END reg_addr[4]
  PIN reg_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 80.640 4.000 81.200 ;
    END
  END reg_addr[5]
  PIN reg_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 68.320 4.000 68.880 ;
    END
  END reg_addr[6]
  PIN reg_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 56.000 4.000 56.560 ;
    END
  END reg_addr[7]
  PIN reg_addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 43.680 4.000 44.240 ;
    END
  END reg_addr[8]
  PIN reg_be[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 191.520 4.000 192.080 ;
    END
  END reg_be[0]
  PIN reg_be[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 179.200 4.000 179.760 ;
    END
  END reg_be[1]
  PIN reg_be[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 166.880 4.000 167.440 ;
    END
  END reg_be[2]
  PIN reg_be[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 154.560 4.000 155.120 ;
    END
  END reg_be[3]
  PIN reg_cs
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 19.040 4.000 19.600 ;
    END
  END reg_cs
  PIN reg_rdata[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 980.000 4.000 980.560 ;
    END
  END reg_rdata[0]
  PIN reg_rdata[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 856.800 4.000 857.360 ;
    END
  END reg_rdata[10]
  PIN reg_rdata[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 844.480 4.000 845.040 ;
    END
  END reg_rdata[11]
  PIN reg_rdata[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 832.160 4.000 832.720 ;
    END
  END reg_rdata[12]
  PIN reg_rdata[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 819.840 4.000 820.400 ;
    END
  END reg_rdata[13]
  PIN reg_rdata[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 807.520 4.000 808.080 ;
    END
  END reg_rdata[14]
  PIN reg_rdata[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 795.200 4.000 795.760 ;
    END
  END reg_rdata[15]
  PIN reg_rdata[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 782.880 4.000 783.440 ;
    END
  END reg_rdata[16]
  PIN reg_rdata[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 770.560 4.000 771.120 ;
    END
  END reg_rdata[17]
  PIN reg_rdata[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 758.240 4.000 758.800 ;
    END
  END reg_rdata[18]
  PIN reg_rdata[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 745.920 4.000 746.480 ;
    END
  END reg_rdata[19]
  PIN reg_rdata[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 967.680 4.000 968.240 ;
    END
  END reg_rdata[1]
  PIN reg_rdata[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 733.600 4.000 734.160 ;
    END
  END reg_rdata[20]
  PIN reg_rdata[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 721.280 4.000 721.840 ;
    END
  END reg_rdata[21]
  PIN reg_rdata[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 708.960 4.000 709.520 ;
    END
  END reg_rdata[22]
  PIN reg_rdata[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 696.640 4.000 697.200 ;
    END
  END reg_rdata[23]
  PIN reg_rdata[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 684.320 4.000 684.880 ;
    END
  END reg_rdata[24]
  PIN reg_rdata[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 672.000 4.000 672.560 ;
    END
  END reg_rdata[25]
  PIN reg_rdata[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 659.680 4.000 660.240 ;
    END
  END reg_rdata[26]
  PIN reg_rdata[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 647.360 4.000 647.920 ;
    END
  END reg_rdata[27]
  PIN reg_rdata[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 635.040 4.000 635.600 ;
    END
  END reg_rdata[28]
  PIN reg_rdata[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 622.720 4.000 623.280 ;
    END
  END reg_rdata[29]
  PIN reg_rdata[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 955.360 4.000 955.920 ;
    END
  END reg_rdata[2]
  PIN reg_rdata[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 610.400 4.000 610.960 ;
    END
  END reg_rdata[30]
  PIN reg_rdata[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 598.080 4.000 598.640 ;
    END
  END reg_rdata[31]
  PIN reg_rdata[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 943.040 4.000 943.600 ;
    END
  END reg_rdata[3]
  PIN reg_rdata[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 930.720 4.000 931.280 ;
    END
  END reg_rdata[4]
  PIN reg_rdata[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 918.400 4.000 918.960 ;
    END
  END reg_rdata[5]
  PIN reg_rdata[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 906.080 4.000 906.640 ;
    END
  END reg_rdata[6]
  PIN reg_rdata[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 893.760 4.000 894.320 ;
    END
  END reg_rdata[7]
  PIN reg_rdata[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 881.440 4.000 882.000 ;
    END
  END reg_rdata[8]
  PIN reg_rdata[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 869.120 4.000 869.680 ;
    END
  END reg_rdata[9]
  PIN reg_wdata[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 585.760 4.000 586.320 ;
    END
  END reg_wdata[0]
  PIN reg_wdata[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 462.560 4.000 463.120 ;
    END
  END reg_wdata[10]
  PIN reg_wdata[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 450.240 4.000 450.800 ;
    END
  END reg_wdata[11]
  PIN reg_wdata[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 437.920 4.000 438.480 ;
    END
  END reg_wdata[12]
  PIN reg_wdata[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 425.600 4.000 426.160 ;
    END
  END reg_wdata[13]
  PIN reg_wdata[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 413.280 4.000 413.840 ;
    END
  END reg_wdata[14]
  PIN reg_wdata[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 400.960 4.000 401.520 ;
    END
  END reg_wdata[15]
  PIN reg_wdata[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 388.640 4.000 389.200 ;
    END
  END reg_wdata[16]
  PIN reg_wdata[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 376.320 4.000 376.880 ;
    END
  END reg_wdata[17]
  PIN reg_wdata[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 364.000 4.000 364.560 ;
    END
  END reg_wdata[18]
  PIN reg_wdata[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 351.680 4.000 352.240 ;
    END
  END reg_wdata[19]
  PIN reg_wdata[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 573.440 4.000 574.000 ;
    END
  END reg_wdata[1]
  PIN reg_wdata[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 339.360 4.000 339.920 ;
    END
  END reg_wdata[20]
  PIN reg_wdata[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 327.040 4.000 327.600 ;
    END
  END reg_wdata[21]
  PIN reg_wdata[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 314.720 4.000 315.280 ;
    END
  END reg_wdata[22]
  PIN reg_wdata[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 302.400 4.000 302.960 ;
    END
  END reg_wdata[23]
  PIN reg_wdata[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 290.080 4.000 290.640 ;
    END
  END reg_wdata[24]
  PIN reg_wdata[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 277.760 4.000 278.320 ;
    END
  END reg_wdata[25]
  PIN reg_wdata[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 265.440 4.000 266.000 ;
    END
  END reg_wdata[26]
  PIN reg_wdata[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 253.120 4.000 253.680 ;
    END
  END reg_wdata[27]
  PIN reg_wdata[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 240.800 4.000 241.360 ;
    END
  END reg_wdata[28]
  PIN reg_wdata[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 228.480 4.000 229.040 ;
    END
  END reg_wdata[29]
  PIN reg_wdata[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 561.120 4.000 561.680 ;
    END
  END reg_wdata[2]
  PIN reg_wdata[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 216.160 4.000 216.720 ;
    END
  END reg_wdata[30]
  PIN reg_wdata[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 203.840 4.000 204.400 ;
    END
  END reg_wdata[31]
  PIN reg_wdata[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 548.800 4.000 549.360 ;
    END
  END reg_wdata[3]
  PIN reg_wdata[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 536.480 4.000 537.040 ;
    END
  END reg_wdata[4]
  PIN reg_wdata[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 524.160 4.000 524.720 ;
    END
  END reg_wdata[5]
  PIN reg_wdata[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 511.840 4.000 512.400 ;
    END
  END reg_wdata[6]
  PIN reg_wdata[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 499.520 4.000 500.080 ;
    END
  END reg_wdata[7]
  PIN reg_wdata[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 487.200 4.000 487.760 ;
    END
  END reg_wdata[8]
  PIN reg_wdata[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 474.880 4.000 475.440 ;
    END
  END reg_wdata[9]
  PIN reg_wr
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 31.360 4.000 31.920 ;
    END
  END reg_wr
  PIN scl_pad_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 21.280 996.000 21.840 1000.000 ;
    END
  END scl_pad_i
  PIN scl_pad_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 54.880 996.000 55.440 1000.000 ;
    END
  END scl_pad_o
  PIN scl_pad_oen_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 88.480 996.000 89.040 1000.000 ;
    END
  END scl_pad_oen_o
  PIN sda_pad_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 122.080 996.000 122.640 1000.000 ;
    END
  END sda_pad_i
  PIN sda_pad_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 155.680 996.000 156.240 1000.000 ;
    END
  END sda_pad_o
  PIN sda_padoen_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 189.280 996.000 189.840 1000.000 ;
    END
  END sda_padoen_o
  PIN spi_rstn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 592.480 996.000 593.040 1000.000 ;
    END
  END spi_rstn
  PIN sspim_sck
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 626.080 996.000 626.640 1000.000 ;
    END
  END sspim_sck
  PIN sspim_si
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 659.680 996.000 660.240 1000.000 ;
    END
  END sspim_si
  PIN sspim_so
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 693.280 996.000 693.840 1000.000 ;
    END
  END sspim_so
  PIN sspim_ssn[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 827.680 996.000 828.240 1000.000 ;
    END
  END sspim_ssn[0]
  PIN sspim_ssn[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 794.080 996.000 794.640 1000.000 ;
    END
  END sspim_ssn[1]
  PIN sspim_ssn[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 760.480 996.000 761.040 1000.000 ;
    END
  END sspim_ssn[2]
  PIN sspim_ssn[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 726.880 996.000 727.440 1000.000 ;
    END
  END sspim_ssn[3]
  PIN uart_rstn[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 424.480 0.000 425.040 4.000 ;
    END
  END uart_rstn[0]
  PIN uart_rstn[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 255.360 0.000 255.920 4.000 ;
    END
  END uart_rstn[1]
  PIN uart_rxd[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 222.880 996.000 223.440 1000.000 ;
    END
  END uart_rxd[0]
  PIN uart_rxd[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 290.080 996.000 290.640 1000.000 ;
    END
  END uart_rxd[1]
  PIN uart_txd[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 256.480 996.000 257.040 1000.000 ;
    END
  END uart_txd[0]
  PIN uart_txd[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 323.680 996.000 324.240 1000.000 ;
    END
  END uart_txd[1]
  PIN usb_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 86.240 0.000 86.800 4.000 ;
    END
  END usb_clk
  PIN usb_in_dn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 390.880 996.000 391.440 1000.000 ;
    END
  END usb_in_dn
  PIN usb_in_dp
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 357.280 996.000 357.840 1000.000 ;
    END
  END usb_in_dp
  PIN usb_intr_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 558.880 996.000 559.440 1000.000 ;
    END
  END usb_intr_o
  PIN usb_out_dn
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal2 ;
        RECT 458.080 996.000 458.640 1000.000 ;
    END
  END usb_out_dn
  PIN usb_out_dp
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 424.480 996.000 425.040 1000.000 ;
    END
  END usb_out_dp
  PIN usb_out_tx_oen
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 491.680 996.000 492.240 1000.000 ;
    END
  END usb_out_tx_oen
  PIN usb_rstn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 762.720 0.000 763.280 4.000 ;
    END
  END usb_rstn
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 842.800 984.890 ;
      LAYER Metal2 ;
        RECT 7.420 995.700 20.980 996.660 ;
        RECT 22.140 995.700 54.580 996.660 ;
        RECT 55.740 995.700 88.180 996.660 ;
        RECT 89.340 995.700 121.780 996.660 ;
        RECT 122.940 995.700 155.380 996.660 ;
        RECT 156.540 995.700 188.980 996.660 ;
        RECT 190.140 995.700 222.580 996.660 ;
        RECT 223.740 995.700 256.180 996.660 ;
        RECT 257.340 995.700 289.780 996.660 ;
        RECT 290.940 995.700 323.380 996.660 ;
        RECT 324.540 995.700 356.980 996.660 ;
        RECT 358.140 995.700 390.580 996.660 ;
        RECT 391.740 995.700 424.180 996.660 ;
        RECT 425.340 995.700 457.780 996.660 ;
        RECT 458.940 995.700 491.380 996.660 ;
        RECT 492.540 995.700 524.980 996.660 ;
        RECT 526.140 995.700 558.580 996.660 ;
        RECT 559.740 995.700 592.180 996.660 ;
        RECT 593.340 995.700 625.780 996.660 ;
        RECT 626.940 995.700 659.380 996.660 ;
        RECT 660.540 995.700 692.980 996.660 ;
        RECT 694.140 995.700 726.580 996.660 ;
        RECT 727.740 995.700 760.180 996.660 ;
        RECT 761.340 995.700 793.780 996.660 ;
        RECT 794.940 995.700 827.380 996.660 ;
        RECT 828.540 995.700 842.660 996.660 ;
        RECT 7.420 4.300 842.660 995.700 ;
        RECT 7.420 4.000 85.940 4.300 ;
        RECT 87.100 4.000 255.060 4.300 ;
        RECT 256.220 4.000 424.180 4.300 ;
        RECT 425.340 4.000 593.300 4.300 ;
        RECT 594.460 4.000 762.420 4.300 ;
        RECT 763.580 4.000 842.660 4.300 ;
      LAYER Metal3 ;
        RECT 4.300 992.020 842.710 992.740 ;
        RECT 3.500 980.860 842.710 992.020 ;
        RECT 4.300 979.700 842.710 980.860 ;
        RECT 3.500 968.540 842.710 979.700 ;
        RECT 4.300 967.380 842.710 968.540 ;
        RECT 3.500 956.220 842.710 967.380 ;
        RECT 4.300 955.060 842.710 956.220 ;
        RECT 3.500 943.900 842.710 955.060 ;
        RECT 4.300 942.740 842.710 943.900 ;
        RECT 3.500 931.580 842.710 942.740 ;
        RECT 4.300 930.420 842.710 931.580 ;
        RECT 3.500 919.260 842.710 930.420 ;
        RECT 4.300 918.100 842.710 919.260 ;
        RECT 3.500 906.940 842.710 918.100 ;
        RECT 4.300 905.780 842.710 906.940 ;
        RECT 3.500 894.620 842.710 905.780 ;
        RECT 4.300 893.460 842.710 894.620 ;
        RECT 3.500 882.300 842.710 893.460 ;
        RECT 4.300 881.140 842.710 882.300 ;
        RECT 3.500 869.980 842.710 881.140 ;
        RECT 4.300 868.820 842.710 869.980 ;
        RECT 3.500 857.660 842.710 868.820 ;
        RECT 4.300 856.500 842.710 857.660 ;
        RECT 3.500 845.340 842.710 856.500 ;
        RECT 4.300 844.180 842.710 845.340 ;
        RECT 3.500 833.020 842.710 844.180 ;
        RECT 4.300 831.860 842.710 833.020 ;
        RECT 3.500 820.700 842.710 831.860 ;
        RECT 4.300 819.540 842.710 820.700 ;
        RECT 3.500 808.380 842.710 819.540 ;
        RECT 4.300 807.220 842.710 808.380 ;
        RECT 3.500 796.060 842.710 807.220 ;
        RECT 4.300 794.900 842.710 796.060 ;
        RECT 3.500 783.740 842.710 794.900 ;
        RECT 4.300 782.580 842.710 783.740 ;
        RECT 3.500 771.420 842.710 782.580 ;
        RECT 4.300 770.260 842.710 771.420 ;
        RECT 3.500 759.100 842.710 770.260 ;
        RECT 4.300 757.940 842.710 759.100 ;
        RECT 3.500 746.780 842.710 757.940 ;
        RECT 4.300 745.620 842.710 746.780 ;
        RECT 3.500 734.460 842.710 745.620 ;
        RECT 4.300 733.300 842.710 734.460 ;
        RECT 3.500 722.140 842.710 733.300 ;
        RECT 4.300 720.980 842.710 722.140 ;
        RECT 3.500 709.820 842.710 720.980 ;
        RECT 4.300 708.660 842.710 709.820 ;
        RECT 3.500 697.500 842.710 708.660 ;
        RECT 4.300 696.340 842.710 697.500 ;
        RECT 3.500 685.180 842.710 696.340 ;
        RECT 4.300 684.020 842.710 685.180 ;
        RECT 3.500 672.860 842.710 684.020 ;
        RECT 4.300 671.700 842.710 672.860 ;
        RECT 3.500 660.540 842.710 671.700 ;
        RECT 4.300 659.380 842.710 660.540 ;
        RECT 3.500 648.220 842.710 659.380 ;
        RECT 4.300 647.060 842.710 648.220 ;
        RECT 3.500 635.900 842.710 647.060 ;
        RECT 4.300 634.740 842.710 635.900 ;
        RECT 3.500 623.580 842.710 634.740 ;
        RECT 4.300 622.420 842.710 623.580 ;
        RECT 3.500 611.260 842.710 622.420 ;
        RECT 4.300 610.100 842.710 611.260 ;
        RECT 3.500 598.940 842.710 610.100 ;
        RECT 4.300 597.780 842.710 598.940 ;
        RECT 3.500 586.620 842.710 597.780 ;
        RECT 4.300 585.460 842.710 586.620 ;
        RECT 3.500 574.300 842.710 585.460 ;
        RECT 4.300 573.140 842.710 574.300 ;
        RECT 3.500 561.980 842.710 573.140 ;
        RECT 4.300 560.820 842.710 561.980 ;
        RECT 3.500 549.660 842.710 560.820 ;
        RECT 4.300 548.500 842.710 549.660 ;
        RECT 3.500 537.340 842.710 548.500 ;
        RECT 4.300 536.180 842.710 537.340 ;
        RECT 3.500 525.020 842.710 536.180 ;
        RECT 4.300 523.860 842.710 525.020 ;
        RECT 3.500 512.700 842.710 523.860 ;
        RECT 4.300 511.540 842.710 512.700 ;
        RECT 3.500 500.380 842.710 511.540 ;
        RECT 4.300 499.220 842.710 500.380 ;
        RECT 3.500 488.060 842.710 499.220 ;
        RECT 4.300 486.900 842.710 488.060 ;
        RECT 3.500 475.740 842.710 486.900 ;
        RECT 4.300 474.580 842.710 475.740 ;
        RECT 3.500 463.420 842.710 474.580 ;
        RECT 4.300 462.260 842.710 463.420 ;
        RECT 3.500 451.100 842.710 462.260 ;
        RECT 4.300 449.940 842.710 451.100 ;
        RECT 3.500 438.780 842.710 449.940 ;
        RECT 4.300 437.620 842.710 438.780 ;
        RECT 3.500 426.460 842.710 437.620 ;
        RECT 4.300 425.300 842.710 426.460 ;
        RECT 3.500 414.140 842.710 425.300 ;
        RECT 4.300 412.980 842.710 414.140 ;
        RECT 3.500 401.820 842.710 412.980 ;
        RECT 4.300 400.660 842.710 401.820 ;
        RECT 3.500 389.500 842.710 400.660 ;
        RECT 4.300 388.340 842.710 389.500 ;
        RECT 3.500 377.180 842.710 388.340 ;
        RECT 4.300 376.020 842.710 377.180 ;
        RECT 3.500 364.860 842.710 376.020 ;
        RECT 4.300 363.700 842.710 364.860 ;
        RECT 3.500 352.540 842.710 363.700 ;
        RECT 4.300 351.380 842.710 352.540 ;
        RECT 3.500 340.220 842.710 351.380 ;
        RECT 4.300 339.060 842.710 340.220 ;
        RECT 3.500 327.900 842.710 339.060 ;
        RECT 4.300 326.740 842.710 327.900 ;
        RECT 3.500 315.580 842.710 326.740 ;
        RECT 4.300 314.420 842.710 315.580 ;
        RECT 3.500 303.260 842.710 314.420 ;
        RECT 4.300 302.100 842.710 303.260 ;
        RECT 3.500 290.940 842.710 302.100 ;
        RECT 4.300 289.780 842.710 290.940 ;
        RECT 3.500 278.620 842.710 289.780 ;
        RECT 4.300 277.460 842.710 278.620 ;
        RECT 3.500 266.300 842.710 277.460 ;
        RECT 4.300 265.140 842.710 266.300 ;
        RECT 3.500 253.980 842.710 265.140 ;
        RECT 4.300 252.820 842.710 253.980 ;
        RECT 3.500 241.660 842.710 252.820 ;
        RECT 4.300 240.500 842.710 241.660 ;
        RECT 3.500 229.340 842.710 240.500 ;
        RECT 4.300 228.180 842.710 229.340 ;
        RECT 3.500 217.020 842.710 228.180 ;
        RECT 4.300 215.860 842.710 217.020 ;
        RECT 3.500 204.700 842.710 215.860 ;
        RECT 4.300 203.540 842.710 204.700 ;
        RECT 3.500 192.380 842.710 203.540 ;
        RECT 4.300 191.220 842.710 192.380 ;
        RECT 3.500 180.060 842.710 191.220 ;
        RECT 4.300 178.900 842.710 180.060 ;
        RECT 3.500 167.740 842.710 178.900 ;
        RECT 4.300 166.580 842.710 167.740 ;
        RECT 3.500 155.420 842.710 166.580 ;
        RECT 4.300 154.260 842.710 155.420 ;
        RECT 3.500 143.100 842.710 154.260 ;
        RECT 4.300 141.940 842.710 143.100 ;
        RECT 3.500 130.780 842.710 141.940 ;
        RECT 4.300 129.620 842.710 130.780 ;
        RECT 3.500 118.460 842.710 129.620 ;
        RECT 4.300 117.300 842.710 118.460 ;
        RECT 3.500 106.140 842.710 117.300 ;
        RECT 4.300 104.980 842.710 106.140 ;
        RECT 3.500 93.820 842.710 104.980 ;
        RECT 4.300 92.660 842.710 93.820 ;
        RECT 3.500 81.500 842.710 92.660 ;
        RECT 4.300 80.340 842.710 81.500 ;
        RECT 3.500 69.180 842.710 80.340 ;
        RECT 4.300 68.020 842.710 69.180 ;
        RECT 3.500 56.860 842.710 68.020 ;
        RECT 4.300 55.700 842.710 56.860 ;
        RECT 3.500 44.540 842.710 55.700 ;
        RECT 4.300 43.380 842.710 44.540 ;
        RECT 3.500 32.220 842.710 43.380 ;
        RECT 4.300 31.060 842.710 32.220 ;
        RECT 3.500 19.900 842.710 31.060 ;
        RECT 4.300 18.740 842.710 19.900 ;
        RECT 3.500 7.580 842.710 18.740 ;
        RECT 4.300 6.860 842.710 7.580 ;
      LAYER Metal4 ;
        RECT 10.220 21.930 19.640 981.030 ;
        RECT 26.440 21.930 69.640 981.030 ;
        RECT 76.440 21.930 119.640 981.030 ;
        RECT 126.440 21.930 169.640 981.030 ;
        RECT 176.440 21.930 219.640 981.030 ;
        RECT 226.440 21.930 269.640 981.030 ;
        RECT 276.440 21.930 319.640 981.030 ;
        RECT 326.440 21.930 369.640 981.030 ;
        RECT 376.440 21.930 419.640 981.030 ;
        RECT 426.440 21.930 469.640 981.030 ;
        RECT 476.440 21.930 519.640 981.030 ;
        RECT 526.440 21.930 569.640 981.030 ;
        RECT 576.440 21.930 619.640 981.030 ;
        RECT 626.440 21.930 669.640 981.030 ;
        RECT 676.440 21.930 719.640 981.030 ;
        RECT 726.440 21.930 769.640 981.030 ;
        RECT 776.440 21.930 819.640 981.030 ;
        RECT 826.440 21.930 839.860 981.030 ;
      LAYER Metal5 ;
        RECT 10.700 32.630 828.740 941.170 ;
  END
END uart_i2c_usb_spi_top
END LIBRARY

