VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO pinmux_top
  CLASS BLOCK ;
  FOREIGN pinmux_top ;
  ORIGIN 0.000 0.000 ;
  SIZE 900.000 BY 1000.000 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 15.380 331.040 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 483.040 15.380 484.640 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 636.640 15.380 638.240 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 790.240 15.380 791.840 984.220 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 406.240 15.380 407.840 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 559.840 15.380 561.440 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 713.440 15.380 715.040 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 867.040 15.380 868.640 984.220 ;
    END
  END VSS
  PIN cfg_strap_pad_ctrl
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 45.920 4.000 46.480 ;
    END
  END cfg_strap_pad_ctrl
  PIN digital_io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 31.360 900.000 31.920 ;
    END
  END digital_io_in[0]
  PIN digital_io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 669.760 900.000 670.320 ;
    END
  END digital_io_in[10]
  PIN digital_io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 733.600 900.000 734.160 ;
    END
  END digital_io_in[11]
  PIN digital_io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 797.440 900.000 798.000 ;
    END
  END digital_io_in[12]
  PIN digital_io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 861.280 900.000 861.840 ;
    END
  END digital_io_in[13]
  PIN digital_io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 925.120 900.000 925.680 ;
    END
  END digital_io_in[14]
  PIN digital_io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 863.520 996.000 864.080 1000.000 ;
    END
  END digital_io_in[15]
  PIN digital_io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 846.720 996.000 847.280 1000.000 ;
    END
  END digital_io_in[16]
  PIN digital_io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 829.920 996.000 830.480 1000.000 ;
    END
  END digital_io_in[17]
  PIN digital_io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 813.120 996.000 813.680 1000.000 ;
    END
  END digital_io_in[18]
  PIN digital_io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 796.320 996.000 796.880 1000.000 ;
    END
  END digital_io_in[19]
  PIN digital_io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 95.200 900.000 95.760 ;
    END
  END digital_io_in[1]
  PIN digital_io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 779.520 996.000 780.080 1000.000 ;
    END
  END digital_io_in[20]
  PIN digital_io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 762.720 996.000 763.280 1000.000 ;
    END
  END digital_io_in[21]
  PIN digital_io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 745.920 996.000 746.480 1000.000 ;
    END
  END digital_io_in[22]
  PIN digital_io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 729.120 996.000 729.680 1000.000 ;
    END
  END digital_io_in[23]
  PIN digital_io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 253.120 996.000 253.680 1000.000 ;
    END
  END digital_io_in[24]
  PIN digital_io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 236.320 996.000 236.880 1000.000 ;
    END
  END digital_io_in[25]
  PIN digital_io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 219.520 996.000 220.080 1000.000 ;
    END
  END digital_io_in[26]
  PIN digital_io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 202.720 996.000 203.280 1000.000 ;
    END
  END digital_io_in[27]
  PIN digital_io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 185.920 996.000 186.480 1000.000 ;
    END
  END digital_io_in[28]
  PIN digital_io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 169.120 996.000 169.680 1000.000 ;
    END
  END digital_io_in[29]
  PIN digital_io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 159.040 900.000 159.600 ;
    END
  END digital_io_in[2]
  PIN digital_io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 152.320 996.000 152.880 1000.000 ;
    END
  END digital_io_in[30]
  PIN digital_io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 135.520 996.000 136.080 1000.000 ;
    END
  END digital_io_in[31]
  PIN digital_io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 118.720 996.000 119.280 1000.000 ;
    END
  END digital_io_in[32]
  PIN digital_io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 101.920 996.000 102.480 1000.000 ;
    END
  END digital_io_in[33]
  PIN digital_io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 85.120 996.000 85.680 1000.000 ;
    END
  END digital_io_in[34]
  PIN digital_io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 68.320 996.000 68.880 1000.000 ;
    END
  END digital_io_in[35]
  PIN digital_io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 51.520 996.000 52.080 1000.000 ;
    END
  END digital_io_in[36]
  PIN digital_io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 34.720 996.000 35.280 1000.000 ;
    END
  END digital_io_in[37]
  PIN digital_io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 222.880 900.000 223.440 ;
    END
  END digital_io_in[3]
  PIN digital_io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 286.720 900.000 287.280 ;
    END
  END digital_io_in[4]
  PIN digital_io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 350.560 900.000 351.120 ;
    END
  END digital_io_in[5]
  PIN digital_io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 414.400 900.000 414.960 ;
    END
  END digital_io_in[6]
  PIN digital_io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 478.240 900.000 478.800 ;
    END
  END digital_io_in[7]
  PIN digital_io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 542.080 900.000 542.640 ;
    END
  END digital_io_in[8]
  PIN digital_io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 605.920 900.000 606.480 ;
    END
  END digital_io_in[9]
  PIN digital_io_oen[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 73.920 900.000 74.480 ;
    END
  END digital_io_oen[0]
  PIN digital_io_oen[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 712.320 900.000 712.880 ;
    END
  END digital_io_oen[10]
  PIN digital_io_oen[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 776.160 900.000 776.720 ;
    END
  END digital_io_oen[11]
  PIN digital_io_oen[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 840.000 900.000 840.560 ;
    END
  END digital_io_oen[12]
  PIN digital_io_oen[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 903.840 900.000 904.400 ;
    END
  END digital_io_oen[13]
  PIN digital_io_oen[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 967.680 900.000 968.240 ;
    END
  END digital_io_oen[14]
  PIN digital_io_oen[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 874.720 996.000 875.280 1000.000 ;
    END
  END digital_io_oen[15]
  PIN digital_io_oen[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 857.920 996.000 858.480 1000.000 ;
    END
  END digital_io_oen[16]
  PIN digital_io_oen[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 841.120 996.000 841.680 1000.000 ;
    END
  END digital_io_oen[17]
  PIN digital_io_oen[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal2 ;
        RECT 824.320 996.000 824.880 1000.000 ;
    END
  END digital_io_oen[18]
  PIN digital_io_oen[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 807.520 996.000 808.080 1000.000 ;
    END
  END digital_io_oen[19]
  PIN digital_io_oen[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 137.760 900.000 138.320 ;
    END
  END digital_io_oen[1]
  PIN digital_io_oen[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 790.720 996.000 791.280 1000.000 ;
    END
  END digital_io_oen[20]
  PIN digital_io_oen[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 773.920 996.000 774.480 1000.000 ;
    END
  END digital_io_oen[21]
  PIN digital_io_oen[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 757.120 996.000 757.680 1000.000 ;
    END
  END digital_io_oen[22]
  PIN digital_io_oen[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 740.320 996.000 740.880 1000.000 ;
    END
  END digital_io_oen[23]
  PIN digital_io_oen[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 241.920 996.000 242.480 1000.000 ;
    END
  END digital_io_oen[24]
  PIN digital_io_oen[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 225.120 996.000 225.680 1000.000 ;
    END
  END digital_io_oen[25]
  PIN digital_io_oen[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 208.320 996.000 208.880 1000.000 ;
    END
  END digital_io_oen[26]
  PIN digital_io_oen[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 191.520 996.000 192.080 1000.000 ;
    END
  END digital_io_oen[27]
  PIN digital_io_oen[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 174.720 996.000 175.280 1000.000 ;
    END
  END digital_io_oen[28]
  PIN digital_io_oen[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 157.920 996.000 158.480 1000.000 ;
    END
  END digital_io_oen[29]
  PIN digital_io_oen[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 201.600 900.000 202.160 ;
    END
  END digital_io_oen[2]
  PIN digital_io_oen[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 141.120 996.000 141.680 1000.000 ;
    END
  END digital_io_oen[30]
  PIN digital_io_oen[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 124.320 996.000 124.880 1000.000 ;
    END
  END digital_io_oen[31]
  PIN digital_io_oen[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 107.520 996.000 108.080 1000.000 ;
    END
  END digital_io_oen[32]
  PIN digital_io_oen[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 90.720 996.000 91.280 1000.000 ;
    END
  END digital_io_oen[33]
  PIN digital_io_oen[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 73.920 996.000 74.480 1000.000 ;
    END
  END digital_io_oen[34]
  PIN digital_io_oen[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 57.120 996.000 57.680 1000.000 ;
    END
  END digital_io_oen[35]
  PIN digital_io_oen[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 40.320 996.000 40.880 1000.000 ;
    END
  END digital_io_oen[36]
  PIN digital_io_oen[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 23.520 996.000 24.080 1000.000 ;
    END
  END digital_io_oen[37]
  PIN digital_io_oen[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 265.440 900.000 266.000 ;
    END
  END digital_io_oen[3]
  PIN digital_io_oen[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 329.280 900.000 329.840 ;
    END
  END digital_io_oen[4]
  PIN digital_io_oen[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 393.120 900.000 393.680 ;
    END
  END digital_io_oen[5]
  PIN digital_io_oen[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 456.960 900.000 457.520 ;
    END
  END digital_io_oen[6]
  PIN digital_io_oen[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 520.800 900.000 521.360 ;
    END
  END digital_io_oen[7]
  PIN digital_io_oen[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 584.640 900.000 585.200 ;
    END
  END digital_io_oen[8]
  PIN digital_io_oen[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 648.480 900.000 649.040 ;
    END
  END digital_io_oen[9]
  PIN digital_io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 52.640 900.000 53.200 ;
    END
  END digital_io_out[0]
  PIN digital_io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 691.040 900.000 691.600 ;
    END
  END digital_io_out[10]
  PIN digital_io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 754.880 900.000 755.440 ;
    END
  END digital_io_out[11]
  PIN digital_io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 818.720 900.000 819.280 ;
    END
  END digital_io_out[12]
  PIN digital_io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 882.560 900.000 883.120 ;
    END
  END digital_io_out[13]
  PIN digital_io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 946.400 900.000 946.960 ;
    END
  END digital_io_out[14]
  PIN digital_io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 869.120 996.000 869.680 1000.000 ;
    END
  END digital_io_out[15]
  PIN digital_io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal2 ;
        RECT 852.320 996.000 852.880 1000.000 ;
    END
  END digital_io_out[16]
  PIN digital_io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 835.520 996.000 836.080 1000.000 ;
    END
  END digital_io_out[17]
  PIN digital_io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 818.720 996.000 819.280 1000.000 ;
    END
  END digital_io_out[18]
  PIN digital_io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 801.920 996.000 802.480 1000.000 ;
    END
  END digital_io_out[19]
  PIN digital_io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 116.480 900.000 117.040 ;
    END
  END digital_io_out[1]
  PIN digital_io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 785.120 996.000 785.680 1000.000 ;
    END
  END digital_io_out[20]
  PIN digital_io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 768.320 996.000 768.880 1000.000 ;
    END
  END digital_io_out[21]
  PIN digital_io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 751.520 996.000 752.080 1000.000 ;
    END
  END digital_io_out[22]
  PIN digital_io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 734.720 996.000 735.280 1000.000 ;
    END
  END digital_io_out[23]
  PIN digital_io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 247.520 996.000 248.080 1000.000 ;
    END
  END digital_io_out[24]
  PIN digital_io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 230.720 996.000 231.280 1000.000 ;
    END
  END digital_io_out[25]
  PIN digital_io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 213.920 996.000 214.480 1000.000 ;
    END
  END digital_io_out[26]
  PIN digital_io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 197.120 996.000 197.680 1000.000 ;
    END
  END digital_io_out[27]
  PIN digital_io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 180.320 996.000 180.880 1000.000 ;
    END
  END digital_io_out[28]
  PIN digital_io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 163.520 996.000 164.080 1000.000 ;
    END
  END digital_io_out[29]
  PIN digital_io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 180.320 900.000 180.880 ;
    END
  END digital_io_out[2]
  PIN digital_io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 146.720 996.000 147.280 1000.000 ;
    END
  END digital_io_out[30]
  PIN digital_io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 129.920 996.000 130.480 1000.000 ;
    END
  END digital_io_out[31]
  PIN digital_io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 113.120 996.000 113.680 1000.000 ;
    END
  END digital_io_out[32]
  PIN digital_io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 96.320 996.000 96.880 1000.000 ;
    END
  END digital_io_out[33]
  PIN digital_io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 79.520 996.000 80.080 1000.000 ;
    END
  END digital_io_out[34]
  PIN digital_io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 62.720 996.000 63.280 1000.000 ;
    END
  END digital_io_out[35]
  PIN digital_io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 45.920 996.000 46.480 1000.000 ;
    END
  END digital_io_out[36]
  PIN digital_io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 29.120 996.000 29.680 1000.000 ;
    END
  END digital_io_out[37]
  PIN digital_io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 244.160 900.000 244.720 ;
    END
  END digital_io_out[3]
  PIN digital_io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 308.000 900.000 308.560 ;
    END
  END digital_io_out[4]
  PIN digital_io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 371.840 900.000 372.400 ;
    END
  END digital_io_out[5]
  PIN digital_io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 435.680 900.000 436.240 ;
    END
  END digital_io_out[6]
  PIN digital_io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 499.520 900.000 500.080 ;
    END
  END digital_io_out[7]
  PIN digital_io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 563.360 900.000 563.920 ;
    END
  END digital_io_out[8]
  PIN digital_io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 627.200 900.000 627.760 ;
    END
  END digital_io_out[9]
  PIN e_reset_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 34.720 4.000 35.280 ;
    END
  END e_reset_n
  PIN i2cm_clk_i
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 449.120 0.000 449.680 4.000 ;
    END
  END i2cm_clk_i
  PIN i2cm_clk_o
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 425.600 0.000 426.160 4.000 ;
    END
  END i2cm_clk_o
  PIN i2cm_clk_oen
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 472.640 0.000 473.200 4.000 ;
    END
  END i2cm_clk_oen
  PIN i2cm_data_i
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 543.200 0.000 543.760 4.000 ;
    END
  END i2cm_data_i
  PIN i2cm_data_o
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 519.680 0.000 520.240 4.000 ;
    END
  END i2cm_data_o
  PIN i2cm_data_oen
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 496.160 0.000 496.720 4.000 ;
    END
  END i2cm_data_oen
  PIN i2cm_intr
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 754.880 0.000 755.440 4.000 ;
    END
  END i2cm_intr
  PIN i2cm_rst_n
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 96.320 0.000 96.880 4.000 ;
    END
  END i2cm_rst_n
  PIN mclk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 57.120 4.000 57.680 ;
    END
  END mclk
  PIN p_reset_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 23.520 4.000 24.080 ;
    END
  END p_reset_n
  PIN pulse1m_mclk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 731.360 0.000 731.920 4.000 ;
    END
  END pulse1m_mclk
  PIN reg_ack
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 975.520 4.000 976.080 ;
    END
  END reg_ack
  PIN reg_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 202.720 4.000 203.280 ;
    END
  END reg_addr[0]
  PIN reg_addr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 90.720 4.000 91.280 ;
    END
  END reg_addr[10]
  PIN reg_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 191.520 4.000 192.080 ;
    END
  END reg_addr[1]
  PIN reg_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.408000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 180.320 4.000 180.880 ;
    END
  END reg_addr[2]
  PIN reg_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 169.120 4.000 169.680 ;
    END
  END reg_addr[3]
  PIN reg_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 157.920 4.000 158.480 ;
    END
  END reg_addr[4]
  PIN reg_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 146.720 4.000 147.280 ;
    END
  END reg_addr[5]
  PIN reg_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 135.520 4.000 136.080 ;
    END
  END reg_addr[6]
  PIN reg_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 124.320 4.000 124.880 ;
    END
  END reg_addr[7]
  PIN reg_addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 113.120 4.000 113.680 ;
    END
  END reg_addr[8]
  PIN reg_addr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 101.920 4.000 102.480 ;
    END
  END reg_addr[9]
  PIN reg_be[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 247.520 4.000 248.080 ;
    END
  END reg_be[0]
  PIN reg_be[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 236.320 4.000 236.880 ;
    END
  END reg_be[1]
  PIN reg_be[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 225.120 4.000 225.680 ;
    END
  END reg_be[2]
  PIN reg_be[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 213.920 4.000 214.480 ;
    END
  END reg_be[3]
  PIN reg_cs
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 68.320 4.000 68.880 ;
    END
  END reg_cs
  PIN reg_peri_ack
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 723.520 996.000 724.080 1000.000 ;
    END
  END reg_peri_ack
  PIN reg_peri_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 337.120 996.000 337.680 1000.000 ;
    END
  END reg_peri_addr[0]
  PIN reg_peri_addr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 281.120 996.000 281.680 1000.000 ;
    END
  END reg_peri_addr[10]
  PIN reg_peri_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 331.520 996.000 332.080 1000.000 ;
    END
  END reg_peri_addr[1]
  PIN reg_peri_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 325.920 996.000 326.480 1000.000 ;
    END
  END reg_peri_addr[2]
  PIN reg_peri_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 320.320 996.000 320.880 1000.000 ;
    END
  END reg_peri_addr[3]
  PIN reg_peri_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 314.720 996.000 315.280 1000.000 ;
    END
  END reg_peri_addr[4]
  PIN reg_peri_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 309.120 996.000 309.680 1000.000 ;
    END
  END reg_peri_addr[5]
  PIN reg_peri_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 303.520 996.000 304.080 1000.000 ;
    END
  END reg_peri_addr[6]
  PIN reg_peri_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 297.920 996.000 298.480 1000.000 ;
    END
  END reg_peri_addr[7]
  PIN reg_peri_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 292.320 996.000 292.880 1000.000 ;
    END
  END reg_peri_addr[8]
  PIN reg_peri_addr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 286.720 996.000 287.280 1000.000 ;
    END
  END reg_peri_addr[9]
  PIN reg_peri_be[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 359.520 996.000 360.080 1000.000 ;
    END
  END reg_peri_be[0]
  PIN reg_peri_be[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 353.920 996.000 354.480 1000.000 ;
    END
  END reg_peri_be[1]
  PIN reg_peri_be[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 348.320 996.000 348.880 1000.000 ;
    END
  END reg_peri_be[2]
  PIN reg_peri_be[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 342.720 996.000 343.280 1000.000 ;
    END
  END reg_peri_be[3]
  PIN reg_peri_cs
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 269.920 996.000 270.480 1000.000 ;
    END
  END reg_peri_cs
  PIN reg_peri_rdata[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 717.920 996.000 718.480 1000.000 ;
    END
  END reg_peri_rdata[0]
  PIN reg_peri_rdata[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 661.920 996.000 662.480 1000.000 ;
    END
  END reg_peri_rdata[10]
  PIN reg_peri_rdata[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 656.320 996.000 656.880 1000.000 ;
    END
  END reg_peri_rdata[11]
  PIN reg_peri_rdata[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 650.720 996.000 651.280 1000.000 ;
    END
  END reg_peri_rdata[12]
  PIN reg_peri_rdata[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 645.120 996.000 645.680 1000.000 ;
    END
  END reg_peri_rdata[13]
  PIN reg_peri_rdata[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 639.520 996.000 640.080 1000.000 ;
    END
  END reg_peri_rdata[14]
  PIN reg_peri_rdata[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 633.920 996.000 634.480 1000.000 ;
    END
  END reg_peri_rdata[15]
  PIN reg_peri_rdata[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 628.320 996.000 628.880 1000.000 ;
    END
  END reg_peri_rdata[16]
  PIN reg_peri_rdata[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 622.720 996.000 623.280 1000.000 ;
    END
  END reg_peri_rdata[17]
  PIN reg_peri_rdata[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 617.120 996.000 617.680 1000.000 ;
    END
  END reg_peri_rdata[18]
  PIN reg_peri_rdata[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 611.520 996.000 612.080 1000.000 ;
    END
  END reg_peri_rdata[19]
  PIN reg_peri_rdata[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 712.320 996.000 712.880 1000.000 ;
    END
  END reg_peri_rdata[1]
  PIN reg_peri_rdata[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 605.920 996.000 606.480 1000.000 ;
    END
  END reg_peri_rdata[20]
  PIN reg_peri_rdata[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 600.320 996.000 600.880 1000.000 ;
    END
  END reg_peri_rdata[21]
  PIN reg_peri_rdata[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 594.720 996.000 595.280 1000.000 ;
    END
  END reg_peri_rdata[22]
  PIN reg_peri_rdata[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 589.120 996.000 589.680 1000.000 ;
    END
  END reg_peri_rdata[23]
  PIN reg_peri_rdata[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 583.520 996.000 584.080 1000.000 ;
    END
  END reg_peri_rdata[24]
  PIN reg_peri_rdata[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 577.920 996.000 578.480 1000.000 ;
    END
  END reg_peri_rdata[25]
  PIN reg_peri_rdata[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 572.320 996.000 572.880 1000.000 ;
    END
  END reg_peri_rdata[26]
  PIN reg_peri_rdata[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 566.720 996.000 567.280 1000.000 ;
    END
  END reg_peri_rdata[27]
  PIN reg_peri_rdata[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 561.120 996.000 561.680 1000.000 ;
    END
  END reg_peri_rdata[28]
  PIN reg_peri_rdata[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 555.520 996.000 556.080 1000.000 ;
    END
  END reg_peri_rdata[29]
  PIN reg_peri_rdata[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 706.720 996.000 707.280 1000.000 ;
    END
  END reg_peri_rdata[2]
  PIN reg_peri_rdata[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 549.920 996.000 550.480 1000.000 ;
    END
  END reg_peri_rdata[30]
  PIN reg_peri_rdata[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 544.320 996.000 544.880 1000.000 ;
    END
  END reg_peri_rdata[31]
  PIN reg_peri_rdata[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 701.120 996.000 701.680 1000.000 ;
    END
  END reg_peri_rdata[3]
  PIN reg_peri_rdata[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 695.520 996.000 696.080 1000.000 ;
    END
  END reg_peri_rdata[4]
  PIN reg_peri_rdata[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 689.920 996.000 690.480 1000.000 ;
    END
  END reg_peri_rdata[5]
  PIN reg_peri_rdata[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 684.320 996.000 684.880 1000.000 ;
    END
  END reg_peri_rdata[6]
  PIN reg_peri_rdata[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 678.720 996.000 679.280 1000.000 ;
    END
  END reg_peri_rdata[7]
  PIN reg_peri_rdata[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 673.120 996.000 673.680 1000.000 ;
    END
  END reg_peri_rdata[8]
  PIN reg_peri_rdata[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 667.520 996.000 668.080 1000.000 ;
    END
  END reg_peri_rdata[9]
  PIN reg_peri_wdata[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 538.720 996.000 539.280 1000.000 ;
    END
  END reg_peri_wdata[0]
  PIN reg_peri_wdata[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 482.720 996.000 483.280 1000.000 ;
    END
  END reg_peri_wdata[10]
  PIN reg_peri_wdata[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 477.120 996.000 477.680 1000.000 ;
    END
  END reg_peri_wdata[11]
  PIN reg_peri_wdata[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 471.520 996.000 472.080 1000.000 ;
    END
  END reg_peri_wdata[12]
  PIN reg_peri_wdata[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 465.920 996.000 466.480 1000.000 ;
    END
  END reg_peri_wdata[13]
  PIN reg_peri_wdata[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 460.320 996.000 460.880 1000.000 ;
    END
  END reg_peri_wdata[14]
  PIN reg_peri_wdata[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 454.720 996.000 455.280 1000.000 ;
    END
  END reg_peri_wdata[15]
  PIN reg_peri_wdata[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 449.120 996.000 449.680 1000.000 ;
    END
  END reg_peri_wdata[16]
  PIN reg_peri_wdata[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 443.520 996.000 444.080 1000.000 ;
    END
  END reg_peri_wdata[17]
  PIN reg_peri_wdata[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 437.920 996.000 438.480 1000.000 ;
    END
  END reg_peri_wdata[18]
  PIN reg_peri_wdata[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 432.320 996.000 432.880 1000.000 ;
    END
  END reg_peri_wdata[19]
  PIN reg_peri_wdata[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 533.120 996.000 533.680 1000.000 ;
    END
  END reg_peri_wdata[1]
  PIN reg_peri_wdata[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 426.720 996.000 427.280 1000.000 ;
    END
  END reg_peri_wdata[20]
  PIN reg_peri_wdata[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 421.120 996.000 421.680 1000.000 ;
    END
  END reg_peri_wdata[21]
  PIN reg_peri_wdata[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal2 ;
        RECT 415.520 996.000 416.080 1000.000 ;
    END
  END reg_peri_wdata[22]
  PIN reg_peri_wdata[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 409.920 996.000 410.480 1000.000 ;
    END
  END reg_peri_wdata[23]
  PIN reg_peri_wdata[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 404.320 996.000 404.880 1000.000 ;
    END
  END reg_peri_wdata[24]
  PIN reg_peri_wdata[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 398.720 996.000 399.280 1000.000 ;
    END
  END reg_peri_wdata[25]
  PIN reg_peri_wdata[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 393.120 996.000 393.680 1000.000 ;
    END
  END reg_peri_wdata[26]
  PIN reg_peri_wdata[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 387.520 996.000 388.080 1000.000 ;
    END
  END reg_peri_wdata[27]
  PIN reg_peri_wdata[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 381.920 996.000 382.480 1000.000 ;
    END
  END reg_peri_wdata[28]
  PIN reg_peri_wdata[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 376.320 996.000 376.880 1000.000 ;
    END
  END reg_peri_wdata[29]
  PIN reg_peri_wdata[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 527.520 996.000 528.080 1000.000 ;
    END
  END reg_peri_wdata[2]
  PIN reg_peri_wdata[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 370.720 996.000 371.280 1000.000 ;
    END
  END reg_peri_wdata[30]
  PIN reg_peri_wdata[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 365.120 996.000 365.680 1000.000 ;
    END
  END reg_peri_wdata[31]
  PIN reg_peri_wdata[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 521.920 996.000 522.480 1000.000 ;
    END
  END reg_peri_wdata[3]
  PIN reg_peri_wdata[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 516.320 996.000 516.880 1000.000 ;
    END
  END reg_peri_wdata[4]
  PIN reg_peri_wdata[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 510.720 996.000 511.280 1000.000 ;
    END
  END reg_peri_wdata[5]
  PIN reg_peri_wdata[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 505.120 996.000 505.680 1000.000 ;
    END
  END reg_peri_wdata[6]
  PIN reg_peri_wdata[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 499.520 996.000 500.080 1000.000 ;
    END
  END reg_peri_wdata[7]
  PIN reg_peri_wdata[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 493.920 996.000 494.480 1000.000 ;
    END
  END reg_peri_wdata[8]
  PIN reg_peri_wdata[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 488.320 996.000 488.880 1000.000 ;
    END
  END reg_peri_wdata[9]
  PIN reg_peri_wr
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 275.520 996.000 276.080 1000.000 ;
    END
  END reg_peri_wr
  PIN reg_rdata[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 964.320 4.000 964.880 ;
    END
  END reg_rdata[0]
  PIN reg_rdata[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 852.320 4.000 852.880 ;
    END
  END reg_rdata[10]
  PIN reg_rdata[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 841.120 4.000 841.680 ;
    END
  END reg_rdata[11]
  PIN reg_rdata[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 829.920 4.000 830.480 ;
    END
  END reg_rdata[12]
  PIN reg_rdata[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 818.720 4.000 819.280 ;
    END
  END reg_rdata[13]
  PIN reg_rdata[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 807.520 4.000 808.080 ;
    END
  END reg_rdata[14]
  PIN reg_rdata[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 796.320 4.000 796.880 ;
    END
  END reg_rdata[15]
  PIN reg_rdata[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 785.120 4.000 785.680 ;
    END
  END reg_rdata[16]
  PIN reg_rdata[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 773.920 4.000 774.480 ;
    END
  END reg_rdata[17]
  PIN reg_rdata[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 762.720 4.000 763.280 ;
    END
  END reg_rdata[18]
  PIN reg_rdata[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 751.520 4.000 752.080 ;
    END
  END reg_rdata[19]
  PIN reg_rdata[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 953.120 4.000 953.680 ;
    END
  END reg_rdata[1]
  PIN reg_rdata[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 740.320 4.000 740.880 ;
    END
  END reg_rdata[20]
  PIN reg_rdata[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 729.120 4.000 729.680 ;
    END
  END reg_rdata[21]
  PIN reg_rdata[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 717.920 4.000 718.480 ;
    END
  END reg_rdata[22]
  PIN reg_rdata[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 706.720 4.000 707.280 ;
    END
  END reg_rdata[23]
  PIN reg_rdata[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 695.520 4.000 696.080 ;
    END
  END reg_rdata[24]
  PIN reg_rdata[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 684.320 4.000 684.880 ;
    END
  END reg_rdata[25]
  PIN reg_rdata[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 673.120 4.000 673.680 ;
    END
  END reg_rdata[26]
  PIN reg_rdata[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 661.920 4.000 662.480 ;
    END
  END reg_rdata[27]
  PIN reg_rdata[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 650.720 4.000 651.280 ;
    END
  END reg_rdata[28]
  PIN reg_rdata[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 639.520 4.000 640.080 ;
    END
  END reg_rdata[29]
  PIN reg_rdata[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 941.920 4.000 942.480 ;
    END
  END reg_rdata[2]
  PIN reg_rdata[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 628.320 4.000 628.880 ;
    END
  END reg_rdata[30]
  PIN reg_rdata[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 617.120 4.000 617.680 ;
    END
  END reg_rdata[31]
  PIN reg_rdata[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 930.720 4.000 931.280 ;
    END
  END reg_rdata[3]
  PIN reg_rdata[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 919.520 4.000 920.080 ;
    END
  END reg_rdata[4]
  PIN reg_rdata[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 908.320 4.000 908.880 ;
    END
  END reg_rdata[5]
  PIN reg_rdata[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 897.120 4.000 897.680 ;
    END
  END reg_rdata[6]
  PIN reg_rdata[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 885.920 4.000 886.480 ;
    END
  END reg_rdata[7]
  PIN reg_rdata[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 874.720 4.000 875.280 ;
    END
  END reg_rdata[8]
  PIN reg_rdata[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 863.520 4.000 864.080 ;
    END
  END reg_rdata[9]
  PIN reg_wdata[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 605.920 4.000 606.480 ;
    END
  END reg_wdata[0]
  PIN reg_wdata[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 493.920 4.000 494.480 ;
    END
  END reg_wdata[10]
  PIN reg_wdata[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 482.720 4.000 483.280 ;
    END
  END reg_wdata[11]
  PIN reg_wdata[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 471.520 4.000 472.080 ;
    END
  END reg_wdata[12]
  PIN reg_wdata[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 460.320 4.000 460.880 ;
    END
  END reg_wdata[13]
  PIN reg_wdata[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 449.120 4.000 449.680 ;
    END
  END reg_wdata[14]
  PIN reg_wdata[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 437.920 4.000 438.480 ;
    END
  END reg_wdata[15]
  PIN reg_wdata[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 426.720 4.000 427.280 ;
    END
  END reg_wdata[16]
  PIN reg_wdata[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 415.520 4.000 416.080 ;
    END
  END reg_wdata[17]
  PIN reg_wdata[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 404.320 4.000 404.880 ;
    END
  END reg_wdata[18]
  PIN reg_wdata[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 393.120 4.000 393.680 ;
    END
  END reg_wdata[19]
  PIN reg_wdata[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 594.720 4.000 595.280 ;
    END
  END reg_wdata[1]
  PIN reg_wdata[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 381.920 4.000 382.480 ;
    END
  END reg_wdata[20]
  PIN reg_wdata[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 370.720 4.000 371.280 ;
    END
  END reg_wdata[21]
  PIN reg_wdata[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 359.520 4.000 360.080 ;
    END
  END reg_wdata[22]
  PIN reg_wdata[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 348.320 4.000 348.880 ;
    END
  END reg_wdata[23]
  PIN reg_wdata[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 337.120 4.000 337.680 ;
    END
  END reg_wdata[24]
  PIN reg_wdata[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 325.920 4.000 326.480 ;
    END
  END reg_wdata[25]
  PIN reg_wdata[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 314.720 4.000 315.280 ;
    END
  END reg_wdata[26]
  PIN reg_wdata[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 303.520 4.000 304.080 ;
    END
  END reg_wdata[27]
  PIN reg_wdata[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 292.320 4.000 292.880 ;
    END
  END reg_wdata[28]
  PIN reg_wdata[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 281.120 4.000 281.680 ;
    END
  END reg_wdata[29]
  PIN reg_wdata[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 583.520 4.000 584.080 ;
    END
  END reg_wdata[2]
  PIN reg_wdata[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 269.920 4.000 270.480 ;
    END
  END reg_wdata[30]
  PIN reg_wdata[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 258.720 4.000 259.280 ;
    END
  END reg_wdata[31]
  PIN reg_wdata[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 572.320 4.000 572.880 ;
    END
  END reg_wdata[3]
  PIN reg_wdata[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 561.120 4.000 561.680 ;
    END
  END reg_wdata[4]
  PIN reg_wdata[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 549.920 4.000 550.480 ;
    END
  END reg_wdata[5]
  PIN reg_wdata[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 538.720 4.000 539.280 ;
    END
  END reg_wdata[6]
  PIN reg_wdata[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 527.520 4.000 528.080 ;
    END
  END reg_wdata[7]
  PIN reg_wdata[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 516.320 4.000 516.880 ;
    END
  END reg_wdata[8]
  PIN reg_wdata[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 505.120 4.000 505.680 ;
    END
  END reg_wdata[9]
  PIN reg_wr
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 79.520 4.000 80.080 ;
    END
  END reg_wr
  PIN rtc_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 258.720 996.000 259.280 1000.000 ;
    END
  END rtc_clk
  PIN rtc_intr
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 264.320 996.000 264.880 1000.000 ;
    END
  END rtc_intr
  PIN s_reset_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 848.960 0.000 849.520 4.000 ;
    END
  END s_reset_n
  PIN spim_miso
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 684.320 0.000 684.880 4.000 ;
    END
  END spim_miso
  PIN spim_mosi
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 707.840 0.000 708.400 4.000 ;
    END
  END spim_mosi
  PIN spim_sck
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 566.720 0.000 567.280 4.000 ;
    END
  END spim_sck
  PIN spim_ssn[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 660.800 0.000 661.360 4.000 ;
    END
  END spim_ssn[0]
  PIN spim_ssn[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 637.280 0.000 637.840 4.000 ;
    END
  END spim_ssn[1]
  PIN spim_ssn[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 613.760 0.000 614.320 4.000 ;
    END
  END spim_ssn[2]
  PIN spim_ssn[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 590.240 0.000 590.800 4.000 ;
    END
  END spim_ssn[3]
  PIN sspim_rst_n
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 25.760 0.000 26.320 4.000 ;
    END
  END sspim_rst_n
  PIN uart_rst_n[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 72.800 0.000 73.360 4.000 ;
    END
  END uart_rst_n[0]
  PIN uart_rst_n[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 49.280 0.000 49.840 4.000 ;
    END
  END uart_rst_n[1]
  PIN uart_rxd[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 402.080 0.000 402.640 4.000 ;
    END
  END uart_rxd[0]
  PIN uart_rxd[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 355.040 0.000 355.600 4.000 ;
    END
  END uart_rxd[1]
  PIN uart_txd[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 378.560 0.000 379.120 4.000 ;
    END
  END uart_txd[0]
  PIN uart_txd[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 331.520 0.000 332.080 4.000 ;
    END
  END uart_txd[1]
  PIN usb_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 872.480 0.000 873.040 4.000 ;
    END
  END usb_clk
  PIN usb_dn_i
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 308.000 0.000 308.560 4.000 ;
    END
  END usb_dn_i
  PIN usb_dn_o
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 237.440 0.000 238.000 4.000 ;
    END
  END usb_dn_o
  PIN usb_dp_i
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 284.480 0.000 285.040 4.000 ;
    END
  END usb_dp_i
  PIN usb_dp_o
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 213.920 0.000 214.480 4.000 ;
    END
  END usb_dp_o
  PIN usb_intr
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 778.400 0.000 778.960 4.000 ;
    END
  END usb_intr
  PIN usb_oen
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 260.960 0.000 261.520 4.000 ;
    END
  END usb_oen
  PIN usb_rst_n
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 119.840 0.000 120.400 4.000 ;
    END
  END usb_rst_n
  PIN user_clock1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 801.920 0.000 802.480 4.000 ;
    END
  END user_clock1
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 825.440 0.000 826.000 4.000 ;
    END
  END user_clock2
  PIN user_irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 143.360 0.000 143.920 4.000 ;
    END
  END user_irq[0]
  PIN user_irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 166.880 0.000 167.440 4.000 ;
    END
  END user_irq[1]
  PIN user_irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 190.400 0.000 190.960 4.000 ;
    END
  END user_irq[2]
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 893.200 984.890 ;
      LAYER Metal2 ;
        RECT 7.980 995.700 23.220 996.660 ;
        RECT 24.380 995.700 28.820 996.660 ;
        RECT 29.980 995.700 34.420 996.660 ;
        RECT 35.580 995.700 40.020 996.660 ;
        RECT 41.180 995.700 45.620 996.660 ;
        RECT 46.780 995.700 51.220 996.660 ;
        RECT 52.380 995.700 56.820 996.660 ;
        RECT 57.980 995.700 62.420 996.660 ;
        RECT 63.580 995.700 68.020 996.660 ;
        RECT 69.180 995.700 73.620 996.660 ;
        RECT 74.780 995.700 79.220 996.660 ;
        RECT 80.380 995.700 84.820 996.660 ;
        RECT 85.980 995.700 90.420 996.660 ;
        RECT 91.580 995.700 96.020 996.660 ;
        RECT 97.180 995.700 101.620 996.660 ;
        RECT 102.780 995.700 107.220 996.660 ;
        RECT 108.380 995.700 112.820 996.660 ;
        RECT 113.980 995.700 118.420 996.660 ;
        RECT 119.580 995.700 124.020 996.660 ;
        RECT 125.180 995.700 129.620 996.660 ;
        RECT 130.780 995.700 135.220 996.660 ;
        RECT 136.380 995.700 140.820 996.660 ;
        RECT 141.980 995.700 146.420 996.660 ;
        RECT 147.580 995.700 152.020 996.660 ;
        RECT 153.180 995.700 157.620 996.660 ;
        RECT 158.780 995.700 163.220 996.660 ;
        RECT 164.380 995.700 168.820 996.660 ;
        RECT 169.980 995.700 174.420 996.660 ;
        RECT 175.580 995.700 180.020 996.660 ;
        RECT 181.180 995.700 185.620 996.660 ;
        RECT 186.780 995.700 191.220 996.660 ;
        RECT 192.380 995.700 196.820 996.660 ;
        RECT 197.980 995.700 202.420 996.660 ;
        RECT 203.580 995.700 208.020 996.660 ;
        RECT 209.180 995.700 213.620 996.660 ;
        RECT 214.780 995.700 219.220 996.660 ;
        RECT 220.380 995.700 224.820 996.660 ;
        RECT 225.980 995.700 230.420 996.660 ;
        RECT 231.580 995.700 236.020 996.660 ;
        RECT 237.180 995.700 241.620 996.660 ;
        RECT 242.780 995.700 247.220 996.660 ;
        RECT 248.380 995.700 252.820 996.660 ;
        RECT 253.980 995.700 258.420 996.660 ;
        RECT 259.580 995.700 264.020 996.660 ;
        RECT 265.180 995.700 269.620 996.660 ;
        RECT 270.780 995.700 275.220 996.660 ;
        RECT 276.380 995.700 280.820 996.660 ;
        RECT 281.980 995.700 286.420 996.660 ;
        RECT 287.580 995.700 292.020 996.660 ;
        RECT 293.180 995.700 297.620 996.660 ;
        RECT 298.780 995.700 303.220 996.660 ;
        RECT 304.380 995.700 308.820 996.660 ;
        RECT 309.980 995.700 314.420 996.660 ;
        RECT 315.580 995.700 320.020 996.660 ;
        RECT 321.180 995.700 325.620 996.660 ;
        RECT 326.780 995.700 331.220 996.660 ;
        RECT 332.380 995.700 336.820 996.660 ;
        RECT 337.980 995.700 342.420 996.660 ;
        RECT 343.580 995.700 348.020 996.660 ;
        RECT 349.180 995.700 353.620 996.660 ;
        RECT 354.780 995.700 359.220 996.660 ;
        RECT 360.380 995.700 364.820 996.660 ;
        RECT 365.980 995.700 370.420 996.660 ;
        RECT 371.580 995.700 376.020 996.660 ;
        RECT 377.180 995.700 381.620 996.660 ;
        RECT 382.780 995.700 387.220 996.660 ;
        RECT 388.380 995.700 392.820 996.660 ;
        RECT 393.980 995.700 398.420 996.660 ;
        RECT 399.580 995.700 404.020 996.660 ;
        RECT 405.180 995.700 409.620 996.660 ;
        RECT 410.780 995.700 415.220 996.660 ;
        RECT 416.380 995.700 420.820 996.660 ;
        RECT 421.980 995.700 426.420 996.660 ;
        RECT 427.580 995.700 432.020 996.660 ;
        RECT 433.180 995.700 437.620 996.660 ;
        RECT 438.780 995.700 443.220 996.660 ;
        RECT 444.380 995.700 448.820 996.660 ;
        RECT 449.980 995.700 454.420 996.660 ;
        RECT 455.580 995.700 460.020 996.660 ;
        RECT 461.180 995.700 465.620 996.660 ;
        RECT 466.780 995.700 471.220 996.660 ;
        RECT 472.380 995.700 476.820 996.660 ;
        RECT 477.980 995.700 482.420 996.660 ;
        RECT 483.580 995.700 488.020 996.660 ;
        RECT 489.180 995.700 493.620 996.660 ;
        RECT 494.780 995.700 499.220 996.660 ;
        RECT 500.380 995.700 504.820 996.660 ;
        RECT 505.980 995.700 510.420 996.660 ;
        RECT 511.580 995.700 516.020 996.660 ;
        RECT 517.180 995.700 521.620 996.660 ;
        RECT 522.780 995.700 527.220 996.660 ;
        RECT 528.380 995.700 532.820 996.660 ;
        RECT 533.980 995.700 538.420 996.660 ;
        RECT 539.580 995.700 544.020 996.660 ;
        RECT 545.180 995.700 549.620 996.660 ;
        RECT 550.780 995.700 555.220 996.660 ;
        RECT 556.380 995.700 560.820 996.660 ;
        RECT 561.980 995.700 566.420 996.660 ;
        RECT 567.580 995.700 572.020 996.660 ;
        RECT 573.180 995.700 577.620 996.660 ;
        RECT 578.780 995.700 583.220 996.660 ;
        RECT 584.380 995.700 588.820 996.660 ;
        RECT 589.980 995.700 594.420 996.660 ;
        RECT 595.580 995.700 600.020 996.660 ;
        RECT 601.180 995.700 605.620 996.660 ;
        RECT 606.780 995.700 611.220 996.660 ;
        RECT 612.380 995.700 616.820 996.660 ;
        RECT 617.980 995.700 622.420 996.660 ;
        RECT 623.580 995.700 628.020 996.660 ;
        RECT 629.180 995.700 633.620 996.660 ;
        RECT 634.780 995.700 639.220 996.660 ;
        RECT 640.380 995.700 644.820 996.660 ;
        RECT 645.980 995.700 650.420 996.660 ;
        RECT 651.580 995.700 656.020 996.660 ;
        RECT 657.180 995.700 661.620 996.660 ;
        RECT 662.780 995.700 667.220 996.660 ;
        RECT 668.380 995.700 672.820 996.660 ;
        RECT 673.980 995.700 678.420 996.660 ;
        RECT 679.580 995.700 684.020 996.660 ;
        RECT 685.180 995.700 689.620 996.660 ;
        RECT 690.780 995.700 695.220 996.660 ;
        RECT 696.380 995.700 700.820 996.660 ;
        RECT 701.980 995.700 706.420 996.660 ;
        RECT 707.580 995.700 712.020 996.660 ;
        RECT 713.180 995.700 717.620 996.660 ;
        RECT 718.780 995.700 723.220 996.660 ;
        RECT 724.380 995.700 728.820 996.660 ;
        RECT 729.980 995.700 734.420 996.660 ;
        RECT 735.580 995.700 740.020 996.660 ;
        RECT 741.180 995.700 745.620 996.660 ;
        RECT 746.780 995.700 751.220 996.660 ;
        RECT 752.380 995.700 756.820 996.660 ;
        RECT 757.980 995.700 762.420 996.660 ;
        RECT 763.580 995.700 768.020 996.660 ;
        RECT 769.180 995.700 773.620 996.660 ;
        RECT 774.780 995.700 779.220 996.660 ;
        RECT 780.380 995.700 784.820 996.660 ;
        RECT 785.980 995.700 790.420 996.660 ;
        RECT 791.580 995.700 796.020 996.660 ;
        RECT 797.180 995.700 801.620 996.660 ;
        RECT 802.780 995.700 807.220 996.660 ;
        RECT 808.380 995.700 812.820 996.660 ;
        RECT 813.980 995.700 818.420 996.660 ;
        RECT 819.580 995.700 824.020 996.660 ;
        RECT 825.180 995.700 829.620 996.660 ;
        RECT 830.780 995.700 835.220 996.660 ;
        RECT 836.380 995.700 840.820 996.660 ;
        RECT 841.980 995.700 846.420 996.660 ;
        RECT 847.580 995.700 852.020 996.660 ;
        RECT 853.180 995.700 857.620 996.660 ;
        RECT 858.780 995.700 863.220 996.660 ;
        RECT 864.380 995.700 868.820 996.660 ;
        RECT 869.980 995.700 874.420 996.660 ;
        RECT 875.580 995.700 891.940 996.660 ;
        RECT 7.980 4.300 891.940 995.700 ;
        RECT 7.980 3.500 25.460 4.300 ;
        RECT 26.620 3.500 48.980 4.300 ;
        RECT 50.140 3.500 72.500 4.300 ;
        RECT 73.660 3.500 96.020 4.300 ;
        RECT 97.180 3.500 119.540 4.300 ;
        RECT 120.700 3.500 143.060 4.300 ;
        RECT 144.220 3.500 166.580 4.300 ;
        RECT 167.740 3.500 190.100 4.300 ;
        RECT 191.260 3.500 213.620 4.300 ;
        RECT 214.780 3.500 237.140 4.300 ;
        RECT 238.300 3.500 260.660 4.300 ;
        RECT 261.820 3.500 284.180 4.300 ;
        RECT 285.340 3.500 307.700 4.300 ;
        RECT 308.860 3.500 331.220 4.300 ;
        RECT 332.380 3.500 354.740 4.300 ;
        RECT 355.900 3.500 378.260 4.300 ;
        RECT 379.420 3.500 401.780 4.300 ;
        RECT 402.940 3.500 425.300 4.300 ;
        RECT 426.460 3.500 448.820 4.300 ;
        RECT 449.980 3.500 472.340 4.300 ;
        RECT 473.500 3.500 495.860 4.300 ;
        RECT 497.020 3.500 519.380 4.300 ;
        RECT 520.540 3.500 542.900 4.300 ;
        RECT 544.060 3.500 566.420 4.300 ;
        RECT 567.580 3.500 589.940 4.300 ;
        RECT 591.100 3.500 613.460 4.300 ;
        RECT 614.620 3.500 636.980 4.300 ;
        RECT 638.140 3.500 660.500 4.300 ;
        RECT 661.660 3.500 684.020 4.300 ;
        RECT 685.180 3.500 707.540 4.300 ;
        RECT 708.700 3.500 731.060 4.300 ;
        RECT 732.220 3.500 754.580 4.300 ;
        RECT 755.740 3.500 778.100 4.300 ;
        RECT 779.260 3.500 801.620 4.300 ;
        RECT 802.780 3.500 825.140 4.300 ;
        RECT 826.300 3.500 848.660 4.300 ;
        RECT 849.820 3.500 872.180 4.300 ;
        RECT 873.340 3.500 891.940 4.300 ;
      LAYER Metal3 ;
        RECT 3.500 976.380 896.000 984.060 ;
        RECT 4.300 975.220 896.000 976.380 ;
        RECT 3.500 968.540 896.000 975.220 ;
        RECT 3.500 967.380 895.700 968.540 ;
        RECT 3.500 965.180 896.000 967.380 ;
        RECT 4.300 964.020 896.000 965.180 ;
        RECT 3.500 953.980 896.000 964.020 ;
        RECT 4.300 952.820 896.000 953.980 ;
        RECT 3.500 947.260 896.000 952.820 ;
        RECT 3.500 946.100 895.700 947.260 ;
        RECT 3.500 942.780 896.000 946.100 ;
        RECT 4.300 941.620 896.000 942.780 ;
        RECT 3.500 931.580 896.000 941.620 ;
        RECT 4.300 930.420 896.000 931.580 ;
        RECT 3.500 925.980 896.000 930.420 ;
        RECT 3.500 924.820 895.700 925.980 ;
        RECT 3.500 920.380 896.000 924.820 ;
        RECT 4.300 919.220 896.000 920.380 ;
        RECT 3.500 909.180 896.000 919.220 ;
        RECT 4.300 908.020 896.000 909.180 ;
        RECT 3.500 904.700 896.000 908.020 ;
        RECT 3.500 903.540 895.700 904.700 ;
        RECT 3.500 897.980 896.000 903.540 ;
        RECT 4.300 896.820 896.000 897.980 ;
        RECT 3.500 886.780 896.000 896.820 ;
        RECT 4.300 885.620 896.000 886.780 ;
        RECT 3.500 883.420 896.000 885.620 ;
        RECT 3.500 882.260 895.700 883.420 ;
        RECT 3.500 875.580 896.000 882.260 ;
        RECT 4.300 874.420 896.000 875.580 ;
        RECT 3.500 864.380 896.000 874.420 ;
        RECT 4.300 863.220 896.000 864.380 ;
        RECT 3.500 862.140 896.000 863.220 ;
        RECT 3.500 860.980 895.700 862.140 ;
        RECT 3.500 853.180 896.000 860.980 ;
        RECT 4.300 852.020 896.000 853.180 ;
        RECT 3.500 841.980 896.000 852.020 ;
        RECT 4.300 840.860 896.000 841.980 ;
        RECT 4.300 840.820 895.700 840.860 ;
        RECT 3.500 839.700 895.700 840.820 ;
        RECT 3.500 830.780 896.000 839.700 ;
        RECT 4.300 829.620 896.000 830.780 ;
        RECT 3.500 819.580 896.000 829.620 ;
        RECT 4.300 818.420 895.700 819.580 ;
        RECT 3.500 808.380 896.000 818.420 ;
        RECT 4.300 807.220 896.000 808.380 ;
        RECT 3.500 798.300 896.000 807.220 ;
        RECT 3.500 797.180 895.700 798.300 ;
        RECT 4.300 797.140 895.700 797.180 ;
        RECT 4.300 796.020 896.000 797.140 ;
        RECT 3.500 785.980 896.000 796.020 ;
        RECT 4.300 784.820 896.000 785.980 ;
        RECT 3.500 777.020 896.000 784.820 ;
        RECT 3.500 775.860 895.700 777.020 ;
        RECT 3.500 774.780 896.000 775.860 ;
        RECT 4.300 773.620 896.000 774.780 ;
        RECT 3.500 763.580 896.000 773.620 ;
        RECT 4.300 762.420 896.000 763.580 ;
        RECT 3.500 755.740 896.000 762.420 ;
        RECT 3.500 754.580 895.700 755.740 ;
        RECT 3.500 752.380 896.000 754.580 ;
        RECT 4.300 751.220 896.000 752.380 ;
        RECT 3.500 741.180 896.000 751.220 ;
        RECT 4.300 740.020 896.000 741.180 ;
        RECT 3.500 734.460 896.000 740.020 ;
        RECT 3.500 733.300 895.700 734.460 ;
        RECT 3.500 729.980 896.000 733.300 ;
        RECT 4.300 728.820 896.000 729.980 ;
        RECT 3.500 718.780 896.000 728.820 ;
        RECT 4.300 717.620 896.000 718.780 ;
        RECT 3.500 713.180 896.000 717.620 ;
        RECT 3.500 712.020 895.700 713.180 ;
        RECT 3.500 707.580 896.000 712.020 ;
        RECT 4.300 706.420 896.000 707.580 ;
        RECT 3.500 696.380 896.000 706.420 ;
        RECT 4.300 695.220 896.000 696.380 ;
        RECT 3.500 691.900 896.000 695.220 ;
        RECT 3.500 690.740 895.700 691.900 ;
        RECT 3.500 685.180 896.000 690.740 ;
        RECT 4.300 684.020 896.000 685.180 ;
        RECT 3.500 673.980 896.000 684.020 ;
        RECT 4.300 672.820 896.000 673.980 ;
        RECT 3.500 670.620 896.000 672.820 ;
        RECT 3.500 669.460 895.700 670.620 ;
        RECT 3.500 662.780 896.000 669.460 ;
        RECT 4.300 661.620 896.000 662.780 ;
        RECT 3.500 651.580 896.000 661.620 ;
        RECT 4.300 650.420 896.000 651.580 ;
        RECT 3.500 649.340 896.000 650.420 ;
        RECT 3.500 648.180 895.700 649.340 ;
        RECT 3.500 640.380 896.000 648.180 ;
        RECT 4.300 639.220 896.000 640.380 ;
        RECT 3.500 629.180 896.000 639.220 ;
        RECT 4.300 628.060 896.000 629.180 ;
        RECT 4.300 628.020 895.700 628.060 ;
        RECT 3.500 626.900 895.700 628.020 ;
        RECT 3.500 617.980 896.000 626.900 ;
        RECT 4.300 616.820 896.000 617.980 ;
        RECT 3.500 606.780 896.000 616.820 ;
        RECT 4.300 605.620 895.700 606.780 ;
        RECT 3.500 595.580 896.000 605.620 ;
        RECT 4.300 594.420 896.000 595.580 ;
        RECT 3.500 585.500 896.000 594.420 ;
        RECT 3.500 584.380 895.700 585.500 ;
        RECT 4.300 584.340 895.700 584.380 ;
        RECT 4.300 583.220 896.000 584.340 ;
        RECT 3.500 573.180 896.000 583.220 ;
        RECT 4.300 572.020 896.000 573.180 ;
        RECT 3.500 564.220 896.000 572.020 ;
        RECT 3.500 563.060 895.700 564.220 ;
        RECT 3.500 561.980 896.000 563.060 ;
        RECT 4.300 560.820 896.000 561.980 ;
        RECT 3.500 550.780 896.000 560.820 ;
        RECT 4.300 549.620 896.000 550.780 ;
        RECT 3.500 542.940 896.000 549.620 ;
        RECT 3.500 541.780 895.700 542.940 ;
        RECT 3.500 539.580 896.000 541.780 ;
        RECT 4.300 538.420 896.000 539.580 ;
        RECT 3.500 528.380 896.000 538.420 ;
        RECT 4.300 527.220 896.000 528.380 ;
        RECT 3.500 521.660 896.000 527.220 ;
        RECT 3.500 520.500 895.700 521.660 ;
        RECT 3.500 517.180 896.000 520.500 ;
        RECT 4.300 516.020 896.000 517.180 ;
        RECT 3.500 505.980 896.000 516.020 ;
        RECT 4.300 504.820 896.000 505.980 ;
        RECT 3.500 500.380 896.000 504.820 ;
        RECT 3.500 499.220 895.700 500.380 ;
        RECT 3.500 494.780 896.000 499.220 ;
        RECT 4.300 493.620 896.000 494.780 ;
        RECT 3.500 483.580 896.000 493.620 ;
        RECT 4.300 482.420 896.000 483.580 ;
        RECT 3.500 479.100 896.000 482.420 ;
        RECT 3.500 477.940 895.700 479.100 ;
        RECT 3.500 472.380 896.000 477.940 ;
        RECT 4.300 471.220 896.000 472.380 ;
        RECT 3.500 461.180 896.000 471.220 ;
        RECT 4.300 460.020 896.000 461.180 ;
        RECT 3.500 457.820 896.000 460.020 ;
        RECT 3.500 456.660 895.700 457.820 ;
        RECT 3.500 449.980 896.000 456.660 ;
        RECT 4.300 448.820 896.000 449.980 ;
        RECT 3.500 438.780 896.000 448.820 ;
        RECT 4.300 437.620 896.000 438.780 ;
        RECT 3.500 436.540 896.000 437.620 ;
        RECT 3.500 435.380 895.700 436.540 ;
        RECT 3.500 427.580 896.000 435.380 ;
        RECT 4.300 426.420 896.000 427.580 ;
        RECT 3.500 416.380 896.000 426.420 ;
        RECT 4.300 415.260 896.000 416.380 ;
        RECT 4.300 415.220 895.700 415.260 ;
        RECT 3.500 414.100 895.700 415.220 ;
        RECT 3.500 405.180 896.000 414.100 ;
        RECT 4.300 404.020 896.000 405.180 ;
        RECT 3.500 393.980 896.000 404.020 ;
        RECT 4.300 392.820 895.700 393.980 ;
        RECT 3.500 382.780 896.000 392.820 ;
        RECT 4.300 381.620 896.000 382.780 ;
        RECT 3.500 372.700 896.000 381.620 ;
        RECT 3.500 371.580 895.700 372.700 ;
        RECT 4.300 371.540 895.700 371.580 ;
        RECT 4.300 370.420 896.000 371.540 ;
        RECT 3.500 360.380 896.000 370.420 ;
        RECT 4.300 359.220 896.000 360.380 ;
        RECT 3.500 351.420 896.000 359.220 ;
        RECT 3.500 350.260 895.700 351.420 ;
        RECT 3.500 349.180 896.000 350.260 ;
        RECT 4.300 348.020 896.000 349.180 ;
        RECT 3.500 337.980 896.000 348.020 ;
        RECT 4.300 336.820 896.000 337.980 ;
        RECT 3.500 330.140 896.000 336.820 ;
        RECT 3.500 328.980 895.700 330.140 ;
        RECT 3.500 326.780 896.000 328.980 ;
        RECT 4.300 325.620 896.000 326.780 ;
        RECT 3.500 315.580 896.000 325.620 ;
        RECT 4.300 314.420 896.000 315.580 ;
        RECT 3.500 308.860 896.000 314.420 ;
        RECT 3.500 307.700 895.700 308.860 ;
        RECT 3.500 304.380 896.000 307.700 ;
        RECT 4.300 303.220 896.000 304.380 ;
        RECT 3.500 293.180 896.000 303.220 ;
        RECT 4.300 292.020 896.000 293.180 ;
        RECT 3.500 287.580 896.000 292.020 ;
        RECT 3.500 286.420 895.700 287.580 ;
        RECT 3.500 281.980 896.000 286.420 ;
        RECT 4.300 280.820 896.000 281.980 ;
        RECT 3.500 270.780 896.000 280.820 ;
        RECT 4.300 269.620 896.000 270.780 ;
        RECT 3.500 266.300 896.000 269.620 ;
        RECT 3.500 265.140 895.700 266.300 ;
        RECT 3.500 259.580 896.000 265.140 ;
        RECT 4.300 258.420 896.000 259.580 ;
        RECT 3.500 248.380 896.000 258.420 ;
        RECT 4.300 247.220 896.000 248.380 ;
        RECT 3.500 245.020 896.000 247.220 ;
        RECT 3.500 243.860 895.700 245.020 ;
        RECT 3.500 237.180 896.000 243.860 ;
        RECT 4.300 236.020 896.000 237.180 ;
        RECT 3.500 225.980 896.000 236.020 ;
        RECT 4.300 224.820 896.000 225.980 ;
        RECT 3.500 223.740 896.000 224.820 ;
        RECT 3.500 222.580 895.700 223.740 ;
        RECT 3.500 214.780 896.000 222.580 ;
        RECT 4.300 213.620 896.000 214.780 ;
        RECT 3.500 203.580 896.000 213.620 ;
        RECT 4.300 202.460 896.000 203.580 ;
        RECT 4.300 202.420 895.700 202.460 ;
        RECT 3.500 201.300 895.700 202.420 ;
        RECT 3.500 192.380 896.000 201.300 ;
        RECT 4.300 191.220 896.000 192.380 ;
        RECT 3.500 181.180 896.000 191.220 ;
        RECT 4.300 180.020 895.700 181.180 ;
        RECT 3.500 169.980 896.000 180.020 ;
        RECT 4.300 168.820 896.000 169.980 ;
        RECT 3.500 159.900 896.000 168.820 ;
        RECT 3.500 158.780 895.700 159.900 ;
        RECT 4.300 158.740 895.700 158.780 ;
        RECT 4.300 157.620 896.000 158.740 ;
        RECT 3.500 147.580 896.000 157.620 ;
        RECT 4.300 146.420 896.000 147.580 ;
        RECT 3.500 138.620 896.000 146.420 ;
        RECT 3.500 137.460 895.700 138.620 ;
        RECT 3.500 136.380 896.000 137.460 ;
        RECT 4.300 135.220 896.000 136.380 ;
        RECT 3.500 125.180 896.000 135.220 ;
        RECT 4.300 124.020 896.000 125.180 ;
        RECT 3.500 117.340 896.000 124.020 ;
        RECT 3.500 116.180 895.700 117.340 ;
        RECT 3.500 113.980 896.000 116.180 ;
        RECT 4.300 112.820 896.000 113.980 ;
        RECT 3.500 102.780 896.000 112.820 ;
        RECT 4.300 101.620 896.000 102.780 ;
        RECT 3.500 96.060 896.000 101.620 ;
        RECT 3.500 94.900 895.700 96.060 ;
        RECT 3.500 91.580 896.000 94.900 ;
        RECT 4.300 90.420 896.000 91.580 ;
        RECT 3.500 80.380 896.000 90.420 ;
        RECT 4.300 79.220 896.000 80.380 ;
        RECT 3.500 74.780 896.000 79.220 ;
        RECT 3.500 73.620 895.700 74.780 ;
        RECT 3.500 69.180 896.000 73.620 ;
        RECT 4.300 68.020 896.000 69.180 ;
        RECT 3.500 57.980 896.000 68.020 ;
        RECT 4.300 56.820 896.000 57.980 ;
        RECT 3.500 53.500 896.000 56.820 ;
        RECT 3.500 52.340 895.700 53.500 ;
        RECT 3.500 46.780 896.000 52.340 ;
        RECT 4.300 45.620 896.000 46.780 ;
        RECT 3.500 35.580 896.000 45.620 ;
        RECT 4.300 34.420 896.000 35.580 ;
        RECT 3.500 32.220 896.000 34.420 ;
        RECT 3.500 31.060 895.700 32.220 ;
        RECT 3.500 24.380 896.000 31.060 ;
        RECT 4.300 23.220 896.000 24.380 ;
        RECT 3.500 15.540 896.000 23.220 ;
      LAYER Metal4 ;
        RECT 16.940 24.730 21.940 982.150 ;
        RECT 24.140 24.730 98.740 982.150 ;
        RECT 100.940 24.730 175.540 982.150 ;
        RECT 177.740 24.730 252.340 982.150 ;
        RECT 254.540 24.730 329.140 982.150 ;
        RECT 331.340 24.730 405.940 982.150 ;
        RECT 408.140 24.730 482.740 982.150 ;
        RECT 484.940 24.730 559.540 982.150 ;
        RECT 561.740 24.730 636.340 982.150 ;
        RECT 638.540 24.730 713.140 982.150 ;
        RECT 715.340 24.730 789.940 982.150 ;
        RECT 792.140 24.730 866.740 982.150 ;
        RECT 868.940 24.730 888.020 982.150 ;
      LAYER Metal5 ;
        RECT 24.700 216.230 812.500 981.670 ;
  END
END pinmux_top
END LIBRARY

