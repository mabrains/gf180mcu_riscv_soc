magic
tech gf180mcuD
magscale 1 5
timestamp 1700411252
<< obsm1 >>
rect 672 754 24304 39230
<< obsm2 >>
rect 798 765 24066 39219
<< metal3 >>
rect 0 38416 200 38472
rect 0 35952 200 36008
rect 0 33488 200 33544
rect 0 31024 200 31080
rect 0 28560 200 28616
rect 0 26096 200 26152
rect 0 23632 200 23688
rect 0 21168 200 21224
rect 0 18704 200 18760
rect 0 16240 200 16296
rect 0 13776 200 13832
rect 0 11312 200 11368
rect 0 8848 200 8904
rect 0 6384 200 6440
rect 0 3920 200 3976
rect 0 1456 200 1512
<< obsm3 >>
rect 126 38502 24071 39214
rect 230 38386 24071 38502
rect 126 36038 24071 38386
rect 230 35922 24071 36038
rect 126 33574 24071 35922
rect 230 33458 24071 33574
rect 126 31110 24071 33458
rect 230 30994 24071 31110
rect 126 28646 24071 30994
rect 230 28530 24071 28646
rect 126 26182 24071 28530
rect 230 26066 24071 26182
rect 126 23718 24071 26066
rect 230 23602 24071 23718
rect 126 21254 24071 23602
rect 230 21138 24071 21254
rect 126 18790 24071 21138
rect 230 18674 24071 18790
rect 126 16326 24071 18674
rect 230 16210 24071 16326
rect 126 13862 24071 16210
rect 230 13746 24071 13862
rect 126 11398 24071 13746
rect 230 11282 24071 11398
rect 126 8934 24071 11282
rect 230 8818 24071 8934
rect 126 6470 24071 8818
rect 230 6354 24071 6470
rect 126 4006 24071 6354
rect 230 3890 24071 4006
rect 126 1542 24071 3890
rect 230 1426 24071 1542
rect 126 770 24071 1426
<< metal4 >>
rect 2224 754 2384 39230
rect 9904 754 10064 39230
rect 17584 754 17744 39230
<< obsm4 >>
rect 1134 1857 2194 33815
rect 2414 1857 9874 33815
rect 10094 1857 17554 33815
rect 17774 1857 19978 33815
<< labels >>
rlabel metal4 s 2224 754 2384 39230 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 17584 754 17744 39230 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 9904 754 10064 39230 6 VSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 1456 200 1512 6 io_in[0]
port 3 nsew signal input
rlabel metal3 s 0 3920 200 3976 6 io_in[1]
port 4 nsew signal input
rlabel metal3 s 0 6384 200 6440 6 io_in[2]
port 5 nsew signal input
rlabel metal3 s 0 8848 200 8904 6 io_in[3]
port 6 nsew signal input
rlabel metal3 s 0 11312 200 11368 6 io_in[4]
port 7 nsew signal input
rlabel metal3 s 0 13776 200 13832 6 io_in[5]
port 8 nsew signal input
rlabel metal3 s 0 16240 200 16296 6 io_in[6]
port 9 nsew signal input
rlabel metal3 s 0 18704 200 18760 6 io_in[7]
port 10 nsew signal input
rlabel metal3 s 0 21168 200 21224 6 io_out[0]
port 11 nsew signal output
rlabel metal3 s 0 23632 200 23688 6 io_out[1]
port 12 nsew signal output
rlabel metal3 s 0 26096 200 26152 6 io_out[2]
port 13 nsew signal output
rlabel metal3 s 0 28560 200 28616 6 io_out[3]
port 14 nsew signal output
rlabel metal3 s 0 31024 200 31080 6 io_out[4]
port 15 nsew signal output
rlabel metal3 s 0 33488 200 33544 6 io_out[5]
port 16 nsew signal output
rlabel metal3 s 0 35952 200 36008 6 io_out[6]
port 17 nsew signal output
rlabel metal3 s 0 38416 200 38472 6 io_out[7]
port 18 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 25000 40000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 2924842
string GDS_FILE /home/farag/carvel_riscv_soc/gf180mcu_riscv_soc/openlane/temp_sensor/runs/23_11_19_18_21/results/signoff/temp_sensor.magic.gds
string GDS_START 439110
<< end >>

